* NGSPICE file created from team_02_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt team_02_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_0_20_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09671_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\] net895 net939 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08731__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11834__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08622_ net73 net1708 net954 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11618__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08553_ _04214_ _04215_ _04224_ net793 net1502 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08484_ _03321_ _04182_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12665__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1071_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14446__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1169_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10693__B _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09105_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\] net710 _04616_ _04618_
+ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09036_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\] net925 net921 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout796_A _06105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold340 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10357__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 team_02_WB.instance_to_wrap.top.a1.row2\[25\] vssd1 vssd1 vccd1 vccd1 net1809
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09762__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A _03027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16874__1418 vssd1 vssd1 vccd1 vccd1 _16874__1418/HI net1418 sky130_fd_sc_hd__conb_1
Xfanout820 _04520_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08970__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15741__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10109__A0 _05580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 net832 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_8
Xfanout842 _04403_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_4
X_09938_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\] net819 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\]
+ _05454_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a221o_1
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_6
XFILLER_0_42_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout864 _04543_ vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout875 _04539_ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_2
XANTENNA__09514__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout886 _04536_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_8
Xfanout897 _04531_ vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_4
X_09869_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\] net740 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\]
+ _05385_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a221o_1
Xhold1040 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11744__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net341 net1902 net489 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__mux2_1
Xhold1062 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1073 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12880_ _07387_ _07399_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__nand2_1
Xhold1084 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1095 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
X_11831_ net337 net2364 net592 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10587__C _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14550_ net1095 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
X_11762_ net333 net2547 net599 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ net1668 _04268_ _04346_ team_02_WB.instance_to_wrap.top.ru.next_read_i vssd1
+ vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__o31a_1
XFILLER_0_3_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10713_ team_02_WB.instance_to_wrap.top.pc\[22\] _06177_ _06229_ vssd1 vssd1 vccd1
+ vccd1 _06230_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14481_ net1118 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XANTENNA__12575__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16247__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11693_ _07138_ _07174_ _07178_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__a21o_1
X_16220_ clknet_leaf_45_wb_clk_i _02360_ _01028_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_16725__1280 vssd1 vssd1 vccd1 vccd1 _16725__1280/HI net1280 sky130_fd_sc_hd__conb_1
XFILLER_0_3_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12034__A0 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input92_A wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] _03023_ _03039_ vssd1
+ vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__o21ai_2
X_10644_ _04338_ _06160_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__or2_2
XFILLER_0_82_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16151_ clknet_leaf_14_wb_clk_i _02291_ _00959_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13363_ net1659 net1017 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[25\]
+ sky130_fd_sc_hd__and2_1
X_10575_ net530 net404 _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15102_ net1098 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
XANTENNA__10060__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ net250 net1875 net565 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__mux2_1
X_16082_ clknet_leaf_3_wb_clk_i _02222_ _00890_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13294_ net2395 net983 net965 _02996_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15033_ net1201 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
XANTENNA__11919__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ net244 net2141 net573 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10348__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12176_ net344 net2309 net462 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08961__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11560__A2 _07046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11848__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11058_ _06431_ _06433_ net396 vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__mux2_1
XANTENNA__09505__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15935_ clknet_leaf_111_wb_clk_i _02075_ _00743_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_60_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10009_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\] net780 net720 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a22o_1
X_15866_ clknet_leaf_120_wb_clk_i _02006_ _00674_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08529__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14817_ net1211 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15797_ clknet_leaf_41_wb_clk_i _01937_ _00605_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14748_ net1149 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12485__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14679_ net1174 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07579__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16418_ clknet_leaf_67_wb_clk_i _02553_ _01226_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11379__A2 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16349_ clknet_leaf_51_wb_clk_i _02489_ _01157_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08244__A2 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10051__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11829__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09744__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07984_ _03601_ _03662_ _03675_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09723_ _05233_ _05235_ _05237_ _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout377_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09654_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\] net787 net703 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08439__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08605_ net91 net2305 net954 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__mux2_1
X_09585_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\] net748 _05097_ _05098_
+ _05101_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[0\] _04177_ vssd1 vssd1 vccd1
+ vccd1 _04221_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout711_A _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12395__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ net1655 net1006 net981 _04167_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout809_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08398_ _04105_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__nor2_1
Xwire506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_85_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire528 _05146_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10360_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09983__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11739__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ _04297_ net943 _04509_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__and3_4
XFILLER_0_131_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10291_ _05788_ _05806_ net968 vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__mux2_1
X_12030_ net320 net1843 net474 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__mux2_1
Xhold170 net134 vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold181 net144 vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout650 _04332_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_2
Xfanout661 net663 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_4
Xfanout672 _05964_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__buf_2
Xfanout683 net685 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_4
X_13981_ net1080 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
Xfanout694 net697 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13295__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15720_ clknet_leaf_19_wb_clk_i _01860_ _00528_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12932_ team_02_WB.instance_to_wrap.top.pc\[26\] _06150_ vssd1 vssd1 vccd1 vccd1
+ _07452_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15651_ clknet_leaf_2_wb_clk_i _01791_ _00459_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12863_ _07381_ _07382_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13047__A2 _07332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14602_ net1142 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11814_ net268 net2701 net589 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15582_ clknet_leaf_114_wb_clk_i _01722_ _00390_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15637__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12794_ net377 _06534_ _07076_ _07127_ _06037_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_55_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09120__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14533_ net1094 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
X_11745_ net265 net2612 net598 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14464_ net1158 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
XANTENNA__10281__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11676_ _05187_ _05206_ _05979_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16203_ clknet_leaf_16_wb_clk_i _02343_ _01011_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13415_ _03018_ _03024_ _03025_ _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_133_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10627_ team_02_WB.instance_to_wrap.top.pc\[27\] _06143_ vssd1 vssd1 vccd1 vccd1
+ _06144_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15787__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14395_ net1157 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16134_ clknet_leaf_44_wb_clk_i _02274_ _00942_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10033__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13346_ team_02_WB.instance_to_wrap.ramload\[8\] net1015 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[8\] sky130_fd_sc_hd__and2_1
X_10558_ _04755_ net386 vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16065_ clknet_leaf_121_wb_clk_i _02205_ _00873_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13277_ team_02_WB.instance_to_wrap.top.pc\[21\] net1053 _06679_ net934 vssd1 vssd1
+ vccd1 vccd1 _02988_ sky130_fd_sc_hd__a22o_1
X_10489_ _05919_ _06005_ _05920_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09187__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15016_ net1235 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12810__A_N _04422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09726__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ net1757 net298 net617 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12159_ net295 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\] net464 vssd1
+ vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13286__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10789__A _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15918_ clknet_leaf_10_wb_clk_i _02058_ _00726_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15849_ clknet_leaf_103_wb_clk_i _01989_ _00657_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09370_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\] net895 net939 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09111__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ _04028_ _04032_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16873__1417 vssd1 vssd1 vccd1 vccd1 _16873__1417/HI net1417 sky130_fd_sc_hd__conb_1
X_08252_ _03957_ _03960_ _03945_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07673__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10272__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08183_ _03882_ _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09818__A _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11221__A1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09965__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput220 net220 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1034_A _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09717__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1201_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07967_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] _03687_ _03688_ vssd1 vssd1
+ vccd1 vccd1 _03690_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout661_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16092__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout759_A _04374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\] net700 _05219_ _05220_
+ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a2111o_1
X_07898_ _03591_ _03620_ _03596_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09350__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09637_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\] net864 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout926_A _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09568_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\] net724 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\]
+ _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09102__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ team_02_WB.instance_to_wrap.top.a1.data\[4\] net958 vssd1 vssd1 vccd1 vccd1
+ _04208_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09499_ _05009_ _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11530_ _06037_ net382 _06296_ _07021_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__a31oi_1
XANTENNA__10263__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11461_ _05512_ _05514_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13200_ net1022 _02953_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__or2_4
X_10412_ _05465_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__or2_1
XANTENNA__10015__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14180_ net1132 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11392_ net606 _06884_ _06890_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__and3_4
XFILLER_0_116_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13131_ _06887_ net232 _02898_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__o22a_1
X_10343_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\] net725 net677 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__a22o_1
XANTENNA__11696__C _07177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09708__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ _07455_ _07456_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__nand2b_1
X_10274_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\] net832 net820 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\]
+ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16435__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net251 net2138 net476 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16821_ net1365 vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__buf_2
XFILLER_0_79_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_50_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout491 _07196_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_122_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16752_ net1296 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_122_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13964_ net1236 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
XANTENNA__11279__B2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09341__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15703_ clknet_leaf_15_wb_clk_i _01843_ _00511_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12915_ _07359_ _07434_ _07358_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16683_ clknet_leaf_73_wb_clk_i _02800_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13895_ net1251 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
XANTENNA__11304__A1_N net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11932__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15634_ clknet_leaf_8_wb_clk_i _01774_ _00442_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ _05061_ _06186_ vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ clknet_leaf_33_wb_clk_i _01705_ _00373_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12777_ _06548_ _06674_ _07266_ _07300_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_48_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ net1074 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10254__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ net333 net2371 net602 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15496_ clknet_leaf_19_wb_clk_i _01636_ _00304_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14447_ net1113 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
X_11659_ _05832_ _05910_ _06429_ _07142_ _07144_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__a41o_1
XFILLER_0_126_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12400__A0 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10006__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11203__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14378_ net1139 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10791__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold906 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16117_ clknet_leaf_43_wb_clk_i _02257_ _00925_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold917 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap636 net637 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_2
X_13329_ team_02_WB.instance_to_wrap.top.a1.nextHex\[2\] team_02_WB.instance_to_wrap.top.a1.nextHex\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[0\] sky130_fd_sc_hd__or2_1
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold939 team_02_WB.instance_to_wrap.ramaddr\[6\] vssd1 vssd1 vccd1 vccd1 net2397
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16048_ clknet_leaf_39_wb_clk_i _02188_ _00856_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_45 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08870_ net1055 net1031 team_02_WB.instance_to_wrap.wb.prev_BUSY_O vssd1 vssd1 vccd1
+ vccd1 _04432_ sky130_fd_sc_hd__or3b_1
XFILLER_0_97_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07821_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] _03541_ _03542_ vssd1 vssd1
+ vccd1 vccd1 _03544_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09092__B _04608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ _03461_ _03462_ _03453_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_105_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12003__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10312__A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07683_ _03375_ _03404_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15952__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11842__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\] net891 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13342__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\] net778 _04868_ _04869_
+ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a211o_1
XANTENNA__08438__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout242_A _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13431__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08304_ net2312 net1007 net982 _04018_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10245__A2 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09284_ _04794_ _04796_ _04798_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__nor4_2
XTAP_TAPCELL_ROW_60_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08235_ _03950_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nand2_2
XANTENNA__12673__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09399__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1249_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08166_ _03839_ net226 _03838_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09938__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15332__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11289__S net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16458__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08097_ net2698 net1007 net982 _03817_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout876_A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09571__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ net1056 _04499_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_76_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09323__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_117_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_67_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ _06078_ _06100_ net408 vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11752__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net356 net1855 net430 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13680_ _03206_ _03210_ net1241 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a21oi_1
X_10892_ net380 _06404_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__or2_1
X_12631_ net1740 net330 net555 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10236__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ clknet_leaf_87_wb_clk_i _01490_ _00163_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_12562_ net321 net2457 net443 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ net1082 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
X_11513_ net669 _06995_ _06996_ net837 _07005_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__o221a_1
XFILLER_0_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12583__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15281_ clknet_leaf_78_wb_clk_i _01425_ _00094_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12493_ net305 net2025 net557 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__mux2_1
XANTENNA__10892__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14232_ net1196 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
XANTENNA__09929__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11444_ _06848_ _06939_ net394 vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14163_ net1163 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11375_ _06873_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_128_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13114_ net978 _07420_ _02882_ _02885_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__o31ai_1
X_10326_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\] net824 net917 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14094_ net1114 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11927__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _07436_ _02827_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12697__A0 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\] net720 net845 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__A2_N net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1220 net1225 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1231 net1237 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__buf_4
XFILLER_0_24_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16872__1416 vssd1 vssd1 vccd1 vccd1 _16872__1416/HI net1416 sky130_fd_sc_hd__conb_1
X_10188_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\] net813 net910 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\]
+ _05704_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__a221o_1
Xfanout1242 net1250 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1253 net1254 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__buf_4
Xfanout1264 net1265 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__buf_2
X_16804_ net1348 vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_2
X_14996_ net1223 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
XANTENNA__09314__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16735_ net1281 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
X_13947_ net1216 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14539__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16666_ clknet_leaf_74_wb_clk_i _02785_ _01408_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15205__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ net1263 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15617_ clknet_leaf_122_wb_clk_i _01757_ _00425_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12829_ team_02_WB.instance_to_wrap.top.i_ready team_02_WB.instance_to_wrap.top.testpc.en_latched
+ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_29_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16597_ clknet_leaf_97_wb_clk_i _02716_ _01390_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10227__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15548_ clknet_leaf_49_wb_clk_i _01688_ _00356_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15479_ clknet_leaf_115_wb_clk_i _01619_ _00287_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ _03733_ _03737_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold703 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold714 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold736 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold758 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09971_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\] net728 _05470_ _05482_
+ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a2111oi_2
Xhold769 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11837__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ net1493 _04443_ net930 vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07616__A team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08853_ net141 net1037 net1034 net1575 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a22o_1
X_07804_ _03481_ _03513_ _03526_ _03485_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08784_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\] net778 net750 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a22o_1
XANTENNA__13637__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09305__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13101__B2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ _03420_ _03427_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__and2_1
XANTENNA__12668__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11112__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1199_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07666_ _03356_ _03360_ _03357_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_62_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10696__B _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09405_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\] net783 net735 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07597_ net1776 net1005 net981 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a21o_1
X_09336_ _04846_ _04848_ _04850_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__or4_1
XANTENNA__10218__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09267_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\] net775 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__a22o_1
XANTENNA__16280__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08831__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ _03918_ _03927_ _03917_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__and3b_1
XANTENNA__13168__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09198_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout993_A _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08149_ _03863_ _03866_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_56_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16819__1363 vssd1 vssd1 vccd1 vccd1 _16819__1363/HI net1363 sky130_fd_sc_hd__conb_1
XFILLER_0_114_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09792__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ net421 _06666_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11747__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\] net828 net824 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11091_ _05972_ _06023_ _06597_ _05975_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _05557_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__nand2_2
XANTENNA__12789__D _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10154__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold30 team_02_WB.instance_to_wrap.top.a1.data\[7\] vssd1 vssd1 vccd1 vccd1 net1488
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_02_WB.instance_to_wrap.top.a1.data\[0\] vssd1 vssd1 vccd1 vccd1 net1499
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 net130 vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ net1202 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold63 _02621_ vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold74 team_02_WB.instance_to_wrap.ramstore\[27\] vssd1 vssd1 vccd1 vccd1 net1532
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_02_WB.START_ADDR_VAL_REG\[1\] vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\] _03284_
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\] vssd1 vssd1 vccd1
+ vccd1 _03287_ sky130_fd_sc_hd__a21o_1
Xhold96 team_02_WB.instance_to_wrap.ramstore\[20\] vssd1 vssd1 vccd1 vccd1 net1554
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14781_ net1087 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
XANTENNA__12578__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ net298 net2161 net479 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10887__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ clknet_leaf_28_wb_clk_i _02654_ _01327_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13732_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\] _03240_ vssd1 vssd1 vccd1
+ vccd1 _03242_ sky130_fd_sc_hd__and2_1
X_10944_ net838 _06426_ _06454_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16451_ clknet_leaf_64_wb_clk_i net1626 _01259_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dfrtp_1
XANTENNA__15378__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13663_ net1468 _04086_ net852 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__mux2_1
X_10875_ net369 _06099_ _06389_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__o21ai_1
X_15402_ clknet_leaf_129_wb_clk_i _01542_ _00210_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12614_ net2297 net262 net553 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__mux2_1
XANTENNA__10209__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16382_ clknet_leaf_92_wb_clk_i _02517_ _01190_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09075__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ _03141_ _03144_ _03146_ _03147_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_22_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_85_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15333_ clknet_leaf_46_wb_clk_i _01476_ _00146_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12545_ net250 net2408 net442 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XANTENNA__08822__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_14_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10090__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15264_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[23\]
+ _00077_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_12476_ net247 net2641 net558 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14215_ net1107 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
XANTENNA_5 _06657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _06922_ _06923_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_39_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15195_ net1261 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09783__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ net1207 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
X_11358_ net952 _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16003__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\] net712 _05822_ _05823_
+ _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_120_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14077_ net1082 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
X_11289_ net2409 net292 net642 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09535__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13028_ _07545_ _07546_ net230 vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1050 team_02_WB.instance_to_wrap.top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1
+ net1050 sky130_fd_sc_hd__clkbuf_2
Xfanout1061 team_02_WB.instance_to_wrap.top.a1.instruction\[5\] vssd1 vssd1 vccd1
+ vccd1 net1061 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1072 net1079 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__buf_4
Xfanout1083 net1088 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1094 net1097 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12488__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ net1238 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13173__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16718_ net1446 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16649_ clknet_leaf_99_wb_clk_i _02768_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_98_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13901__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09066__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09121_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\] net914 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08813__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ _04566_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08003_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] _03723_ _03724_ _03722_ vssd1
+ vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__o211a_1
Xhold500 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold533 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold544 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08730__A team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold555 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold577 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09954_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\] net724 net708 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold599 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1114_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ net1506 _04434_ net930 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09885_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__a22o_1
Xhold1200 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout574_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1211 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08836_ net1540 net1039 net1035 team_02_WB.instance_to_wrap.ramstore\[28\] vssd1
+ vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
Xhold1222 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] vssd1
+ vssd1 vccd1 vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1233 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1244 net184 vssd1 vssd1 vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1277 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\] net786 net736 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\]
+ _04395_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__a221o_1
XANTENNA__12398__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A _04379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1288 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 team_02_WB.instance_to_wrap.ramload\[15\] vssd1 vssd1 vccd1 vccd1 net2757
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16646__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ _03402_ _03429_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08698_ net1001 net849 vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__nand2_1
XANTENNA__08501__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ _03370_ _03371_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10660_ _06128_ _06176_ _04490_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09057__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15670__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09319_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\] net779 net763 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\]
+ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08804__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16871__1415 vssd1 vssd1 vccd1 vccd1 _16871__1415/HI net1415 sky130_fd_sc_hd__conb_1
XFILLER_0_36_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10591_ net379 _06107_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__nor2_1
XANTENNA__10072__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ net318 net2376 net565 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ net296 net1877 net574 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14000_ net1091 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
XANTENNA__09765__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ net414 _06716_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__nand2_1
X_12192_ net294 net2130 net577 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13258__A _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ _06229_ _06650_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13313__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15951_ clknet_leaf_36_wb_clk_i _02091_ _00759_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11074_ _06583_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__inv_2
X_14902_ net1136 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
X_10025_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\] net811 _04559_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\]
+ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__a221o_1
X_15882_ clknet_leaf_128_wb_clk_i _02022_ _00690_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14833_ net1106 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14764_ net1080 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
XANTENNA__12101__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ net241 net2343 net481 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09296__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13715_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\] _03231_ net1240 vssd1
+ vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__a21oi_1
X_16503_ clknet_leaf_28_wb_clk_i _02637_ _01310_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ _06439_ _06440_ net393 vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__mux2_1
X_14695_ net1117 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16434_ clknet_leaf_103_wb_clk_i net1603 _01242_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dfrtp_1
X_13646_ _03109_ _03113_ net1249 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a21o_1
XANTENNA__09048__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10858_ _05966_ _05967_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__nand2_2
XFILLER_0_2_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16365_ clknet_leaf_23_wb_clk_i _02505_ _01173_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13577_ _03106_ net962 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__nand2b_1
X_10789_ _05356_ net406 vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15316_ clknet_leaf_85_wb_clk_i _01459_ _00129_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_12528_ net317 net2555 net446 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16296_ clknet_leaf_19_wb_clk_i _02436_ _01104_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15247_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[6\]
+ _00060_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12459_ net296 net2466 net451 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09756__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15178_ net1243 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XANTENNA__09220__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14129_ net1118 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
XANTENNA__10291__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout309 net311 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09508__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13304__B2 _03001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15543__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_98_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09670_ net521 vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08621_ net74 net1723 net956 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12011__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ _04211_ _04212_ net653 net794 net1513 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a32o_1
XANTENNA__11618__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09287__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16818__1362 vssd1 vssd1 vccd1 vccd1 _16818__1362/HI net1362 sky130_fd_sc_hd__conb_1
XFILLER_0_33_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08483_ net1009 _04168_ net1046 _04181_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__o31a_1
XFILLER_0_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11850__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09039__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13350__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09104_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\] net694 _04619_ _04620_
+ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09035_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\] net800 net861 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12681__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1231_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10990__A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16199__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold330 net120 vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold341 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout691_A _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold352 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09211__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold363 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A _04362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold385 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 net812 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__buf_4
Xfanout821 _04514_ vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_8
Xfanout832 _04508_ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__buf_4
X_09937_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\] net908 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__a22o_1
XANTENNA__10109__A1 _05625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout843 net846 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout956_A _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 _04559_ vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_6
Xfanout865 _04543_ vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout876 _04539_ vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_8
Xfanout887 _04536_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_4
X_09868_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\] net774 net772 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__a22o_1
Xfanout898 _04526_ vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_8
Xhold1030 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1041 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1052 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ net109 net1041 net991 net1680 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__a22o_1
Xhold1063 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\] net922 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__a22o_1
Xhold1085 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1096 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ net332 net2163 net591 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09278__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ net325 net1885 net599 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11760__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14637__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ net1016 team_02_WB.instance_to_wrap.top.ru.next_dready vssd1 vssd1 vccd1
+ vccd1 _00005_ sky130_fd_sc_hd__or2_1
X_10712_ _06178_ _06228_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__and2_1
XANTENNA__10293__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14480_ net1091 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11692_ _04461_ _06109_ _07177_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__or3b_1
XFILLER_0_76_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13431_ team_02_WB.instance_to_wrap.top.lcd.currentState\[5\] net962 net1065 vssd1
+ vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__o21a_1
X_10643_ net1001 _06156_ _06158_ _06159_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__or4b_1
XANTENNA__13231__B1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10045__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16150_ clknet_leaf_47_wb_clk_i _02290_ _00958_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08789__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09986__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13362_ team_02_WB.instance_to_wrap.ramload\[24\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[24\] sky130_fd_sc_hd__and2_1
XFILLER_0_1_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input85_A wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10574_ _05061_ net404 vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09450__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ net1104 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12313_ net252 net1791 net568 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16081_ clknet_leaf_50_wb_clk_i _02221_ _00889_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12591__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13293_ _06883_ _02959_ team_02_WB.instance_to_wrap.top.pc\[13\] net1052 vssd1 vssd1
+ vccd1 vccd1 _02996_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__09738__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15032_ net1203 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
X_12244_ net242 net1698 net575 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__mux2_1
XANTENNA__09202__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_107_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12175_ net348 net2293 net464 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11126_ _06632_ _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__and2_1
XANTENNA__13298__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ net407 _06429_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__or2_1
X_15934_ clknet_leaf_114_wb_clk_i _02074_ _00742_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09910__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\] net764 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__a22o_1
X_15865_ clknet_leaf_112_wb_clk_i _02005_ _00673_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14816_ net1160 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09269__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15796_ clknet_leaf_10_wb_clk_i _01936_ _00604_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11959_ net296 net2108 net586 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14747_ net1156 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
XANTENNA__13470__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10284__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14678_ net1093 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16417_ clknet_leaf_67_wb_clk_i _02552_ _01225_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13629_ _03023_ _03106_ _03169_ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13222__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10036__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11379__A3 _06388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16348_ clknet_leaf_49_wb_clk_i _02488_ _01156_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16341__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09441__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16279_ clknet_leaf_13_wb_clk_i _02419_ _01087_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09729__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10339__A1 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11536__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13101__A1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16491__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12006__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07983_ _03677_ _03704_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__xor2_2
XANTENNA__13289__B1 _06830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11845__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\] net824 net885 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\]
+ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a221o_1
X_16870__1414 vssd1 vssd1 vccd1 vccd1 _16870__1414/HI net1414 sky130_fd_sc_hd__conb_1
XFILLER_0_39_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13345__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\] net719 net711 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08604_ net92 net1624 net956 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XANTENNA__11146__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09584_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\] net676 _05099_ _05100_
+ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08535_ team_02_WB.instance_to_wrap.top.a1.data\[0\] net959 vssd1 vssd1 vccd1 vccd1
+ _04220_ sky130_fd_sc_hd__or2_1
XANTENNA__12676__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13461__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10985__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11580__S net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10275__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15439__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08466_ _04164_ _04166_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09680__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08483__A3 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13213__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout704_A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ _04092_ _04099_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire507 _05667_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_2
Xwire518 _05400_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_2
XANTENNA__10027__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09968__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15589__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10924__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09018_ _04504_ _04519_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10290_ _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold160 team_02_WB.instance_to_wrap.ramstore\[3\] vssd1 vssd1 vccd1 vccd1 net1618
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _02600_ vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _02576_ vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold193 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\] vssd1
+ vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11755__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout651 _04332_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_4
X_13980_ net1145 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
Xfanout673 _04469_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_4
Xfanout684 net685 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_6
Xfanout695 net697 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_4
X_12931_ team_02_WB.instance_to_wrap.top.pc\[27\] _06147_ vssd1 vssd1 vccd1 vccd1
+ _07451_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16214__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15650_ clknet_leaf_123_wb_clk_i _01790_ _00458_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12862_ net514 _05444_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11813_ net261 net2153 net590 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__mux2_1
X_14601_ net1109 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
X_15581_ clknet_leaf_51_wb_clk_i _01721_ _00389_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12793_ net377 _06432_ _07041_ _07316_ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__o211a_1
XANTENNA__12586__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14532_ net1132 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
X_11744_ net258 net2318 net598 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09671__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ net1182 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11675_ _04865_ _05985_ _06531_ _07160_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__or4_2
XFILLER_0_126_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16202_ clknet_leaf_130_wb_clk_i _02342_ _01010_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13414_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09959__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ _06128_ _06142_ _04490_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_24_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14394_ net1167 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
XANTENNA_output191_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09423__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16133_ clknet_leaf_30_wb_clk_i _02273_ _00941_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13345_ team_02_WB.instance_to_wrap.ramload\[7\] net1014 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[7\] sky130_fd_sc_hd__and2_1
XANTENNA__15198__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10557_ _06072_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16064_ clknet_leaf_108_wb_clk_i _02204_ _00872_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13276_ net2289 net984 net964 _02987_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10488_ _05649_ _06004_ _05624_ _05646_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11518__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15015_ net1233 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
X_12227_ net1933 net311 net618 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__mux2_1
X_16817__1361 vssd1 vssd1 vccd1 vccd1 _16817__1361/HI net1361 sky130_fd_sc_hd__conb_1
XFILLER_0_110_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14830__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ net284 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\] net464 vssd1
+ vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11109_ _04470_ _06596_ _06617_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__o21bai_4
XANTENNA_max_cap502_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12089_ net2566 net274 net581 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10789__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15917_ clknet_leaf_24_wb_clk_i _02057_ _00725_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15848_ clknet_leaf_15_wb_clk_i _01988_ _00656_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12496__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15779_ clknet_leaf_2_wb_clk_i _01919_ _00587_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10257__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08320_ _04032_ _04033_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09662__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08251_ _03945_ _03957_ _03960_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__and3_1
XANTENNA__10009__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11206__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ _03888_ _03893_ _03862_ _03878_ _03887_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_83_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput210 net210 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_0_112_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput221 net221 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_101_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08925__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout487_A _07198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13356__A team_02_WB.instance_to_wrap.ramload\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07966_ _03687_ _03688_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10699__B _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\] net715 net845 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\]
+ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07897_ _03588_ _03598_ _03595_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__nor3b_1
XANTENNA_fanout654_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09636_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\] net832 net824 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\]
+ _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__a221o_1
XANTENNA__11307__C net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09567_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\] net744 net704 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout821_A _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout919_A _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08518_ _04207_ net1638 net850 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\] net740 _05011_ _05013_
+ _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_110_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09653__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10799__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08449_ _04153_ _03321_ net1005 net1750 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ net2410 net321 net643 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XANTENNA__09405__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10411_ net517 _05419_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11391_ net976 _06206_ _06885_ _06889_ _06837_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__a311o_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13130_ _07375_ _07376_ _07415_ net977 vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a31o_1
X_10342_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\] net752 net717 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13061_ team_02_WB.instance_to_wrap.top.pc\[25\] _07349_ _02837_ _02841_ vssd1 vssd1
+ vccd1 vccd1 _01506_ sky130_fd_sc_hd__o22a_1
X_10273_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\] _04530_ net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12012_ net239 net2127 net474 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
XANTENNA__08916__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16820_ net1364 vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout470 _07208_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_8
Xfanout481 _07204_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16751_ net1295 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
Xfanout492 _07196_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_122_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13963_ net1251 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15702_ clknet_leaf_62_wb_clk_i _01842_ _00510_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12914_ _04802_ _06150_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__o21bai_1
X_16682_ clknet_leaf_73_wb_clk_i _02799_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13894_ net1239 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
XANTENNA__09892__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15633_ clknet_leaf_50_wb_clk_i _01773_ _00441_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12845_ _05016_ _06184_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10239__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12776_ _06825_ _06854_ _06876_ _06925_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_48_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ clknet_leaf_15_wb_clk_i _01704_ _00372_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09644__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ net1164 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
X_11727_ net325 net2164 net602 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15495_ clknet_leaf_24_wb_clk_i _01635_ _00303_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08852__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11658_ _05830_ _05908_ _05907_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__a21oi_1
X_14446_ net1163 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XANTENNA__11739__A0 _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ net552 _04491_ _04494_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14377_ net1100 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
X_11589_ _05910_ net664 _06113_ _05783_ _07077_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold907 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold918 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16116_ clknet_leaf_11_wb_clk_i _02256_ _00924_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13328_ net1491 _03010_ _03012_ _03292_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[1\]
+ sky130_fd_sc_hd__a22o_1
Xhold929 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16047_ clknet_leaf_34_wb_clk_i _02187_ _00855_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13259_ _02964_ _02976_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12164__A0 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ _03541_ _03542_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15284__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07751_ _03471_ _03472_ _03467_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_105_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10312__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13904__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ _03393_ _03394_ _03369_ _03373_ _03374_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09421_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\] net822 net818 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\]
+ _04931_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09352_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\] net738 net722 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a22o_1
XANTENNA__09096__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09635__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08303_ _04000_ _04007_ _04016_ _03992_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__a31o_2
XFILLER_0_75_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09283_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\] net779 net723 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\]
+ _04799_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08234_ _03897_ _03922_ _03923_ _03913_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08165_ _03880_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout402_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08096_ _03815_ _03816_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09564__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout771_A _04371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08998_ _04295_ net944 _04507_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__and3_4
XANTENNA__07582__B1 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ _03632_ _03634_ _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15777__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _06471_ _06472_ net414 vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09874__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\] net740 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\]
+ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10891_ net410 _06404_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12630_ net2051 net334 net555 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__mux2_1
XANTENNA__11334__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input102_A wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16816__1360 vssd1 vssd1 vccd1 vccd1 _16816__1360/HI net1360 sky130_fd_sc_hd__conb_1
XFILLER_0_116_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09626__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ net317 net2487 net442 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08834__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11512_ net796 _07001_ _07002_ net656 _07004_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__o221a_1
X_14300_ net1151 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15280_ clknet_leaf_78_wb_clk_i _01424_ _00093_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ net298 net2403 net558 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14231_ net1121 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11443_ _06896_ _06938_ net366 vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11197__A1 _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14162_ net1121 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11374_ net423 _06406_ _06872_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__o21a_1
XANTENNA__10944__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ net229 _02884_ _06811_ net233 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10325_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\] net873 _05841_ vssd1
+ vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_128_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14093_ net1132 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _07356_ _07357_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__nand2b_1
X_10256_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\] net744 net740 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1210 net1212 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__buf_4
Xfanout1221 net1223 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1232 net1237 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_4
XANTENNA__12104__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10187_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\] net886 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1243 net1246 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__buf_4
Xfanout1254 net1264 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16803_ net1347 vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_2
Xfanout1265 net38 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14995_ net1221 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
XANTENNA__11943__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16734_ net1458 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
X_13946_ net1216 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09865__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16665_ clknet_leaf_74_wb_clk_i _02784_ _01407_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13877_ net1255 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ clknet_leaf_108_wb_clk_i _01756_ _00424_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09078__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ team_02_WB.instance_to_wrap.top.i_ready team_02_WB.instance_to_wrap.top.testpc.en_latched
+ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16596_ clknet_leaf_97_wb_clk_i _02715_ _01389_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09617__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08825__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15547_ clknet_leaf_127_wb_clk_i _01687_ _00355_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12759_ _04610_ _04653_ _04735_ _04949_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15478_ clknet_leaf_46_wb_clk_i _01618_ _00286_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16082__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14429_ net1081 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold704 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09250__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold715 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold737 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold748 team_02_WB.instance_to_wrap.top.a1.row2\[43\] vssd1 vssd1 vccd1 vccd1 net2206
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\] net676 _05483_ _05486_
+ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a211o_1
Xhold759 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08921_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] net1008 _04232_ _04442_ vssd1
+ vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08852_ net142 net1037 net1033 net1592 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a22o_1
XANTENNA__12014__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10163__A2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ _03481_ _03494_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__nor2_1
X_08783_ _04296_ net848 _04363_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__and3_4
XANTENNA__11853__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07734_ _03419_ _03444_ _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__o21a_2
XANTENNA__11112__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09856__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07665_ _03356_ _03357_ _03361_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__and3b_1
XFILLER_0_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout352_A _07087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09404_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\] net778 _04917_ _04918_
+ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1094_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09069__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07596_ net1009 _03317_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__nand2_4
XFILLER_0_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09335_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\] net810 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\]
+ _04851_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08816__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12684__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1261_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ _04777_ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_79_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08217_ _03900_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__or2_1
XANTENNA__13168__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09197_ net615 vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12376__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11179__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08148_ _03863_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09241__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout986_A _02956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08079_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] _03796_ _03797_ _03798_ vssd1
+ vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__12713__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] net792 net652 _05626_
+ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_120_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11090_ _05127_ _06598_ _05124_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10041_ _05534_ _05556_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__or2_1
XANTENNA__11351__A1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[9\] vssd1 vssd1 vccd1 vccd1
+ net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 team_02_WB.instance_to_wrap.top.a1.data\[4\] vssd1 vssd1 vccd1 vccd1 net1489
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_02_WB.instance_to_wrap.ramaddr\[18\] vssd1 vssd1 vccd1 vccd1 net1500
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold53 _02625_ vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 net182 vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold75 _02589_ vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11763__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13800_ net1552 _03284_ _03286_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__a21oi_1
Xhold86 net113 vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold97 _02582_ vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ net310 net2691 net481 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14780_ net1152 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09847__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13731_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\] _03240_ vssd1 vssd1 vccd1
+ vccd1 _03241_ sky130_fd_sc_hd__or2_1
X_10943_ net668 _06446_ _06455_ _06456_ _06428_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_93_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08992__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11064__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16450_ clknet_leaf_45_wb_clk_i net1632 _01258_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13662_ net1471 _04100_ net852 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10874_ net390 _06074_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15401_ clknet_leaf_120_wb_clk_i _01541_ _00209_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12613_ net2128 net264 net553 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08807__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12594__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11406__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13593_ team_02_WB.instance_to_wrap.top.a1.row2\[1\] _03126_ _03023_ vssd1 vssd1
+ vccd1 vccd1 _03147_ sky130_fd_sc_hd__a21o_1
X_16381_ clknet_leaf_92_wb_clk_i _02516_ _01189_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15332_ clknet_leaf_64_wb_clk_i _01475_ _00145_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12544_ net253 net2345 net445 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15263_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[22\]
+ _00076_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_12475_ net241 net1840 net560 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11426_ net414 _06483_ net423 vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__a21oi_1
X_14214_ net1090 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
X_15194_ net1262 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
XANTENNA__09232__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_6 _06657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_54_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_39_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ net1211 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
XANTENNA__11938__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ net837 _06844_ _06856_ _06842_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15942__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10308_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\] net748 _05824_ vssd1
+ vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__a21o_1
X_14076_ net1149 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
X_11288_ net606 _06783_ _06790_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__and3_4
XANTENNA__10475__A_N net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ _07444_ _07445_ _07446_ _07537_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\] net928 net920 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\]
+ _05755_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_98_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10145__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1040 _04245_ vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__buf_2
Xfanout1051 net1052 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
Xfanout1062 team_02_WB.instance_to_wrap.top.a1.instruction\[4\] vssd1 vssd1 vccd1
+ vccd1 net1062 sky130_fd_sc_hd__buf_2
XFILLER_0_83_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1073 net1079 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
Xfanout1084 net1088 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_4
Xfanout1095 net1097 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09299__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14978_ net1255 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16717_ net1276 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_77_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13929_ net1221 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
XANTENNA__15322__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16648_ clknet_leaf_95_wb_clk_i _02767_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_98_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16579_ clknet_leaf_95_wb_clk_i _02698_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dfxtp_1
X_09120_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\] net833 net829 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\]
+ _04636_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15472__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09471__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09051_ net547 _04565_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08002_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] _03723_ _03724_ vssd1 vssd1
+ vccd1 vccd1 _03725_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09223__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold501 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10908__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold512 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11848__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 team_02_WB.instance_to_wrap.top.a1.row2\[16\] vssd1 vssd1 vccd1 vccd1 net1981
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13629__A _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold534 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold556 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold578 team_02_WB.instance_to_wrap.ramstore\[23\] vssd1 vssd1 vccd1 vccd1 net2036
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09953_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\] net772 net744 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__a22o_1
Xhold589 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11149__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ net1045 _04187_ _04199_ net1008 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__a32o_1
XANTENNA__10136__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\] net813 net906 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1107_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1201 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1223 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ net1615 net1037 net1033 team_02_WB.instance_to_wrap.ramstore\[29\] vssd1
+ vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12679__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1234 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout567_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1245 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] vssd1
+ vssd1 vccd1 vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\] net740 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__a22o_1
Xhold1278 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07717_ _03438_ _03439_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__or2_1
X_08697_ net1001 net849 vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout734_A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08501__A2 _04185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ _03342_ _03360_ _03339_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07579_ net2571 net187 _00017_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout901_A _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12708__A _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\] net731 net707 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__a22o_1
XANTENNA__10941__A2_N net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__A team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10590_ net409 _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09249_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\] _04529_ _04530_
+ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\] _04765_ vssd1 vssd1 vccd1
+ vccd1 _04766_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12349__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15965__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13546__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12260_ net309 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\] net576 vssd1
+ vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09214__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11758__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ _06605_ _06715_ net400 vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12191_ net286 net2593 net579 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__mux2_1
X_11142_ _06178_ _06228_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13313__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11073_ _06104_ _06122_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__nor2_2
X_15950_ clknet_leaf_8_wb_clk_i _02090_ _00758_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10127__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14901_ net1187 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
X_10024_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\] net916 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12589__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15881_ clknet_leaf_103_wb_clk_i _02021_ _00689_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15345__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14832_ net1077 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13077__B2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_101_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14763_ net1200 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11975_ net647 _07203_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16502_ clknet_leaf_37_wb_clk_i _02636_ _01309_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13714_ net1240 _03230_ _03231_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__nor3_1
XFILLER_0_135_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10926_ _06334_ _06337_ net366 vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__mux2_1
X_14694_ net1074 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16433_ clknet_leaf_64_wb_clk_i net1597 _01241_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10857_ net2686 net244 net641 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__mux2_1
X_13645_ net1730 net963 _03192_ net1067 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ clknet_leaf_21_wb_clk_i _02504_ _01172_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ net517 net402 vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__and2_1
X_13576_ team_02_WB.instance_to_wrap.top.a1.row1\[120\] _03116_ _03121_ team_02_WB.instance_to_wrap.top.a1.row1\[112\]
+ _03130_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10063__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10063__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15315_ clknet_leaf_103_wb_clk_i _01458_ _00128_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12527_ net313 net2219 net446 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
X_16295_ clknet_leaf_24_wb_clk_i _02435_ _01103_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15246_ clknet_leaf_61_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[5\]
+ _00059_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09205__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ net308 net1962 net453 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11409_ net837 _06895_ _06902_ _06117_ _06906_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__o221a_1
XFILLER_0_111_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12389_ net285 net2107 net460 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__mux2_1
X_15177_ net1244 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XANTENNA__10366__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16120__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ net1109 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13304__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14059_ net1203 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
XANTENNA__10118__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12499__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08620_ net75 net1784 net955 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10601__A _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08278__A team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08551_ _04208_ _04209_ net653 net793 net1559 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11618__A2 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12815__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08482_ _00017_ _04170_ _04176_ _04180_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09103_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\] net698 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14743__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout315_A _06914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09034_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\] net913 _04530_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\]
+ _04549_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13359__A team_02_WB.instance_to_wrap.ramload\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold320 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _02616_ vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1224_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11554__B2 _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout684_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout800 _04542_ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_4
Xhold386 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 net812 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold397 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08970__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout822 _04514_ vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__buf_4
X_09936_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\] net815 net900 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\]
+ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__a221o_1
Xfanout833 net836 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout844 net846 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__buf_4
Xfanout855 net857 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__buf_6
Xfanout866 net869 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout877 _04539_ vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
X_09867_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\] net766 net754 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\]
+ _05383_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout851_A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1020 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 _04536_ vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_8
Xhold1031 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 _04526_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_4
Xhold1042 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ net1622 net1041 net990 team_02_WB.instance_to_wrap.ramaddr\[13\] vssd1 vssd1
+ vccd1 vccd1 _02607_ sky130_fd_sc_hd__a22o_1
XANTENNA__12202__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09798_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__a22o_1
Xhold1064 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1075 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1097 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08749_ _04296_ net847 _04370_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11760_ net324 net2360 net599 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09683__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _06181_ _06227_ _06182_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11691_ _05738_ _05916_ _07141_ _07176_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__or4_2
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11342__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10642_ _04268_ _06155_ _06157_ _04311_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13430_ _03038_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09435__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13231__B2 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13361_ net2764 net1017 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[23\]
+ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ _05187_ net387 _06089_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14653__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15100_ net1078 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16143__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12312_ net239 net1916 net565 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16080_ clknet_leaf_39_wb_clk_i _02220_ _00888_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13292_ net2004 net983 net965 _02995_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input78_A wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12243_ _04291_ net647 _07188_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__or3_1
X_15031_ net1150 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10348__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12174_ net362 net1968 net465 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16293__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ net410 _06347_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__nand2_1
XANTENNA__08961__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13298__B2 _02998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15933_ clknet_leaf_49_wb_clk_i _02073_ _00741_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11056_ _05950_ _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10007_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\] net696 _05521_ _05523_
+ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11517__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12112__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15864_ clknet_leaf_54_wb_clk_i _02004_ _00672_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14815_ net1182 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
XANTENNA__08529__C _04215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15795_ clknet_leaf_55_wb_clk_i _01935_ _00603_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11951__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14746_ net1181 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
X_11958_ net311 net2650 net588 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__mux2_1
XANTENNA__09674__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10909_ _06419_ _06423_ net607 _06416_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__o211a_4
XFILLER_0_89_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14677_ net1217 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11889_ net300 net2439 net488 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16416_ clknet_leaf_66_wb_clk_i _02551_ _01224_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13628_ team_02_WB.instance_to_wrap.top.a1.row1\[60\] _03117_ _03160_ team_02_WB.instance_to_wrap.top.a1.row1\[108\]
+ _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__a221o_1
XANTENNA__09426__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16347_ clknet_leaf_127_wb_clk_i _02487_ _01155_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13559_ net1050 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] vssd1 vssd1 vccd1
+ vccd1 _03114_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16278_ clknet_leaf_52_wb_clk_i _02418_ _01086_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15229_ clknet_leaf_70_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[20\]
+ _00042_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_114_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11536__A1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07982_ _03677_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__or2_1
XANTENNA__13289__B2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\] net800 net861 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09652_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\] net783 net759 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a22o_1
XANTENNA__12022__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08603_ net93 net1587 net957 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
X_09583_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\] net700 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14738__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08534_ _04219_ net1588 net850 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__mux2_1
XANTENNA__09665__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08465_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] _04158_ _04160_ vssd1 vssd1
+ vccd1 vccd1 _04166_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout432_A _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1174_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16166__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09417__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04070_ vssd1 vssd1 vccd1
+ vccd1 _04105_ sky130_fd_sc_hd__xor2_4
XFILLER_0_18_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire508 net509 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire519 net520 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13285__A1_N _06782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12692__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08471__A team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout899_A _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ _04510_ _04516_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold150 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold161 _02565_ vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold172 team_02_WB.instance_to_wrap.top.a1.row1\[2\] vssd1 vssd1 vccd1 vccd1 net1630
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 team_02_WB.instance_to_wrap.top.a1.hexop\[2\] vssd1 vssd1 vccd1 vccd1 net1641
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold194 team_02_WB.START_ADDR_VAL_REG\[5\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13817__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout641 net642 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_8
Xfanout652 _04331_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_6
X_09919_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\] net736 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__a22o_1
Xfanout663 _06112_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_2
Xfanout674 _04412_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_8
Xfanout685 _04402_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_4
Xfanout696 net697 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_8
X_12930_ team_02_WB.instance_to_wrap.top.pc\[28\] _06143_ vssd1 vssd1 vccd1 vccd1
+ _07450_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_124_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12861_ net514 _05444_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__or2_1
X_14600_ net1178 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11812_ net264 net2628 net590 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__mux2_1
X_15580_ clknet_leaf_45_wb_clk_i _01720_ _00388_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16509__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12792_ _06054_ _06296_ net382 vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11463__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14531_ net1147 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
XANTENNA__09120__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11743_ net249 net1848 net597 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14462_ net1192 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XANTENNA__09408__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11674_ _06373_ _07158_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__or3_1
XANTENNA__10018__A1 _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16201_ clknet_leaf_105_wb_clk_i _02341_ _01009_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13413_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_92_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10625_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] net995 vssd1 vssd1 vccd1
+ vccd1 _06142_ sky130_fd_sc_hd__nand2_1
XANTENNA__15533__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16659__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14393_ net1137 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16132_ clknet_leaf_0_wb_clk_i _02272_ _00940_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09477__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13344_ net1771 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[6\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08092__C1 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10556_ _04802_ net404 vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__nor2_1
XANTENNA_output184_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ clknet_leaf_109_wb_clk_i _02203_ _00871_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13275_ _06648_ _02959_ team_02_WB.instance_to_wrap.top.pc\[22\] net1053 vssd1 vssd1
+ vccd1 vccd1 _02987_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12107__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10487_ _05913_ _06003_ _05914_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11518__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15014_ net1235 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
XANTENNA__15683__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09187__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12226_ net1880 net301 net617 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11946__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12157_ net272 net2006 net462 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11108_ net671 _06603_ _06609_ _06104_ _06616_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12088_ net1751 net288 net582 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
XANTENNA__16039__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15916_ clknet_leaf_25_wb_clk_i _02056_ _00724_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11039_ _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__inv_2
XANTENNA__10151__A team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15847_ clknet_leaf_29_wb_clk_i _01987_ _00655_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15778_ clknet_leaf_125_wb_clk_i _01918_ _00586_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08556__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09111__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14729_ net1099 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08250_ _03956_ _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08181_ _03886_ _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12017__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput200 net200 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput211 net211 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput222 net222 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11856__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10193__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07965_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] _03670_ _03672_ vssd1 vssd1
+ vccd1 vccd1 _03688_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout382_A _06084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09704_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\] net745 net842 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07896_ _03596_ _03597_ _03588_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a21o_1
XANTENNA__09886__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09350__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\] net820 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a22o_1
XANTENNA__12687__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09566_ _05082_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__inv_2
XANTENNA__09638__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09102__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08517_ net1046 _04205_ _04206_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout814_A _04521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09497_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\] net788 net714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08448_ _04149_ _04150_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_81_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08379_ _04084_ _04085_ _04081_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07962__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ _05468_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_22_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11390_ _06200_ net654 _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] _06888_
+ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09810__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\] net773 net749 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13060_ _04280_ _02839_ _02840_ net229 net1027 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__a221o_1
XANTENNA__09169__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10272_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\] net827 net892 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12011_ net244 net2087 net476 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XANTENNA__11766__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10184__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 _07220_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_6
XFILLER_0_79_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout471 _07208_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16750_ net1294 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_45_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout482 net485 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_6
Xfanout493 _07196_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_4
X_13962_ net1251 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15701_ clknet_leaf_43_wb_clk_i _01841_ _00509_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16331__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09341__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ _04842_ _06172_ _07432_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_79_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16681_ clknet_leaf_73_wb_clk_i _02798_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12597__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ net1253 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
X_15632_ clknet_leaf_40_wb_clk_i _01772_ _00440_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12844_ _04971_ _06180_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15563_ clknet_leaf_116_wb_clk_i _01703_ _00371_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12775_ _06360_ _06452_ _07297_ _07298_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16481__CLK clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14514_ net1119 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11726_ net321 net2548 net602 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ clknet_leaf_49_wb_clk_i _01634_ _00302_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14445_ net1141 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
X_11657_ _05832_ _05910_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ net1175 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
X_11588_ _05909_ net658 vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__nand2_1
XANTENNA__09801__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16115_ clknet_leaf_57_wb_clk_i _02255_ _00923_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold908 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13327_ _00009_ team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] vssd1 vssd1 vccd1
+ vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[2\] sky130_fd_sc_hd__or2_1
X_10539_ _05489_ net402 vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold919 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16046_ clknet_leaf_9_wb_clk_i _02186_ _00854_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13258_ _06458_ _02963_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12209_ net346 net2053 net577 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13189_ _04280_ _07395_ _02945_ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a31o_1
XANTENNA__15429__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07750_ _03471_ _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09868__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09332__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09670__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire615_A _04713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ _03393_ _03394_ _03369_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_126_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15579__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16879_ net1423 vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__buf_2
XFILLER_0_36_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09420_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\] net814 net883 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\]
+ _04936_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a221o_1
XANTENNA__12300__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09351_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\] net787 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08302_ _04000_ _04007_ _04016_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__and3_1
X_09282_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\] net751 net738 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08233_ _03913_ _03927_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout228_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09399__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ _03840_ net226 _03847_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08095_ _03782_ _03786_ _03811_ _03785_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_77_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1137_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08359__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout597_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10166__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09571__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _04297_ net943 _04503_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_3_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07948_ _03631_ _03634_ _03637_ _03622_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10602__A2_N _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout931_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07879_ _03571_ _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09618_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\] net692 net843 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__a22o_1
X_10890_ _06404_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09549_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\] net813 net809 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\]
+ _05065_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ net314 net2090 net442 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ net667 _06053_ net377 _07003_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__o31a_1
X_12491_ net310 net2501 net560 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__mux2_1
XANTENNA__08771__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ net1096 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_126_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11442_ _06301_ _06304_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14161_ net1106 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
X_11373_ net374 _06665_ _06871_ net379 vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09177__D _04692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10324_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\] net913 net889 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a22o_1
XANTENNA_input60_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ _07516_ _02883_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__xnor2_1
X_14092_ net1081 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ team_02_WB.instance_to_wrap.top.pc\[28\] _07349_ _02822_ _02826_ vssd1 vssd1
+ vccd1 vccd1 _01509_ sky130_fd_sc_hd__o22a_1
X_10255_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\] net716 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\]
+ _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10157__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1200 net1202 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_4
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1222 net1223 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_4
X_10186_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\] net805 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\]
+ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_33_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1233 net1235 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1244 net1246 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__buf_2
X_16802_ net1346 vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_2
Xfanout1255 net1256 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_4
X_14994_ net1221 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09314__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16733_ net1457 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
XFILLER_0_96_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13945_ net1216 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11525__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12120__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16664_ clknet_leaf_101_wb_clk_i _02783_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13876_ net1261 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15615_ clknet_leaf_110_wb_clk_i _01755_ _00423_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12827_ team_02_WB.instance_to_wrap.top.a1.state\[0\] _07343_ _07345_ _07347_ vssd1
+ vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16595_ clknet_leaf_98_wb_clk_i _02714_ _01388_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15546_ clknet_leaf_119_wb_clk_i _01686_ _00354_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12758_ _05648_ _05915_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16227__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11709_ net250 net2106 net601 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
X_15477_ clknet_leaf_43_wb_clk_i _01617_ _00285_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12689_ net309 net1714 net433 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ net1147 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14359_ net1172 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
Xhold705 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold716 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold727 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold738 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 net181 vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12803__B net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16029_ clknet_leaf_48_wb_clk_i _02169_ _00837_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08920_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] net959 _04212_ _04173_ vssd1
+ vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_1678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09002__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10148__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09553__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ net1669 net1037 net1033 net1663 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a22o_1
XANTENNA__11419__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08761__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _03512_ _03524_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08782_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\] net754 net710 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\]
+ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__a221o_1
XANTENNA__09305__A2 _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ _03413_ _03416_ _03445_ _03455_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08728__B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12030__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07664_ _03384_ _03385_ _03351_ _03383_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_81_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10320__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09403_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\] net727 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\]
+ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07595_ net1009 _03317_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1087_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\] net922 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08816__B2 team_02_WB.instance_to_wrap.ramaddr\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09265_ net538 _04775_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1254_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ _03884_ _03899_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09196_ _04702_ _04707_ _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_75_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11179__A2 _06679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08147_ _03829_ net226 _03835_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_56_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08078_ _03797_ _03798_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__and2_1
XANTENNA__09792__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout979_A _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10139__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ _05534_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold10 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[11\] vssd1 vssd1 vccd1 vccd1
+ net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_02_WB.instance_to_wrap.ramstore\[15\] vssd1 vssd1 vccd1 vccd1 net1479
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 net180 vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 _02612_ vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_02_WB.instance_to_wrap.top.a1.data\[1\] vssd1 vssd1 vccd1 vccd1 net1512
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_02_WB.instance_to_wrap.ramstore\[21\] vssd1 vssd1 vccd1 vccd1 net1523
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_02_WB.instance_to_wrap.top.a1.row1\[105\] vssd1 vssd1 vccd1 vccd1 net1534
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 _02610_ vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11991_ net300 net2332 net479 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
Xhold98 team_02_WB.START_ADDR_VAL_REG\[25\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ _03240_ net949 _03239_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__and3b_1
X_10942_ _04693_ net662 _06453_ net796 vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_129_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13661_ net1478 _04111_ net851 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10873_ _06382_ _06387_ net413 vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15400_ clknet_leaf_14_wb_clk_i _01540_ _00208_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12612_ net1846 net258 net553 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16380_ clknet_leaf_78_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[4\] _01188_
+ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_130_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13592_ team_02_WB.instance_to_wrap.top.a1.row1\[57\] _03117_ _03119_ team_02_WB.instance_to_wrap.top.a1.row1\[1\]
+ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15331_ clknet_leaf_64_wb_clk_i _01474_ _00144_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12543_ net239 net2712 net442 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15262_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[21\]
+ _00075_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10090__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12474_ _04292_ _04452_ _07201_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__or3_4
XFILLER_0_123_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14213_ net1086 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11425_ net375 _06716_ _06921_ net383 vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__a22o_1
X_15193_ net1262 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
XANTENNA_7 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14144_ net1207 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11356_ net667 _06845_ _06852_ _06855_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__o211a_1
XANTENNA__09783__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13316__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10307_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\] net720 net704 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__a22o_1
XANTENNA__12115__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14075_ net1159 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
X_11287_ net974 _06784_ _06789_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13026_ _07444_ _07445_ _07446_ _07537_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__nand4_1
XANTENNA__09535__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11878__A0 _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_89_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\] net884 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1030 _04430_ vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__buf_2
XFILLER_0_98_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11954__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_23_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10169_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\] net877 _05675_ _05685_
+ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a211o_1
Xfanout1052 net1054 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
Xfanout1074 net1079 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_4
Xfanout1085 net1088 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__buf_2
Xfanout1096 net1097 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_4
X_14977_ net1255 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13928_ net1194 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16716_ net1275 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XANTENNA__10302__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16647_ clknet_leaf_99_wb_clk_i _02766_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13859_ net1226 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16578_ clknet_leaf_96_wb_clk_i _00004_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15529_ clknet_leaf_105_wb_clk_i _01669_ _00337_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09050_ net547 _04565_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10081__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08001_ _03305_ net255 _03689_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15767__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10369__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold513 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11030__A1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold524 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold535 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 team_02_WB.instance_to_wrap.ramaddr\[14\] vssd1 vssd1 vccd1 vccd1 net2004
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13307__B1 _07026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold557 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold568 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12025__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09952_ _05468_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__inv_2
Xhold579 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09526__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08903_ team_02_WB.instance_to_wrap.top.edg2.flip2 _04179_ _04182_ team_02_WB.instance_to_wrap.top.edg2.flip1
+ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__and4bb_1
X_09883_ _05384_ _05390_ _05399_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nor3_2
XFILLER_0_42_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout295_A _06791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] vssd1 vssd1 vccd1 vccd1
+ net2660 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ net162 net1040 net1036 net1481 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a22o_1
Xhold1213 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 team_02_WB.instance_to_wrap.ramstore\[28\] vssd1 vssd1 vccd1 vccd1 net2682
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1002_A _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1235 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07643__A team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1246 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 team_02_WB.instance_to_wrap.wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net2715
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13364__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ net847 _04363_ _04364_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout462_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1268 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] vssd1
+ vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1279 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
X_07716_ _03403_ net425 _03408_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__a21boi_1
X_08696_ _04323_ _04324_ _04307_ _04322_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07647_ _03343_ _03360_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__nor2_2
XANTENNA__12695__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout727_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15297__CLK clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07578_ team_02_WB.instance_to_wrap.top.pad.count\[1\] team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__nor2_1
XFILLER_0_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09317_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\] net675 _04824_ _04827_
+ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\] net895 net939 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a22o_1
XANTENNA__10072__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09179_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\] net726 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11210_ _06662_ _06714_ net371 vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__mux2_1
XANTENNA__09765__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12190_ net274 net2530 net577 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11141_ net953 _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__nand2_1
XANTENNA__10244__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09517__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ _04864_ net660 _06122_ _06357_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput100 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14900_ net1075 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
XANTENNA__11774__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\] net928 net884 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\]
+ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__a221o_1
X_15880_ clknet_leaf_16_wb_clk_i _02020_ _00688_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14831_ net1113 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12285__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14762_ net1167 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
X_11974_ _07188_ _07201_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__nor2_1
XANTENNA__09150__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16501_ clknet_leaf_28_wb_clk_i _02635_ _01308_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13713_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\]
+ _03227_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10925_ _06309_ _06331_ net366 vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__mux2_1
X_14693_ net1136 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14386__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16432_ clknet_leaf_64_wb_clk_i net1643 _01240_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dfrtp_1
X_13644_ _03023_ _03185_ _03189_ _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__or4_1
X_10856_ net947 _06365_ _06371_ net607 vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__o211a_4
XFILLER_0_71_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16363_ clknet_leaf_117_wb_clk_i _02503_ _01171_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13575_ team_02_WB.instance_to_wrap.top.a1.row2\[40\] _03123_ _03125_ team_02_WB.instance_to_wrap.top.a1.row2\[32\]
+ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a22o_1
X_10787_ _06299_ _06302_ net365 vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__mux2_1
XANTENNA__10419__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15314_ clknet_leaf_64_wb_clk_i _01457_ _00127_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11260__A1 _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ net304 net2102 net446 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__mux2_1
X_16294_ clknet_leaf_43_wb_clk_i _02434_ _01102_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11949__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15245_ clknet_leaf_61_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[4\]
+ _00058_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12457_ net300 net2088 net451 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09756__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _06037_ _06903_ _06905_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__a21oi_1
X_15176_ net1243 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
X_12388_ net273 net2502 net458 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14127_ net1165 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11339_ net946 _06830_ _06839_ net606 vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__o211a_2
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09508__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ net1163 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
X_13009_ team_02_WB.instance_to_wrap.top.pc\[23\] _06177_ _07528_ vssd1 vssd1 vccd1
+ vccd1 _07529_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire528_A _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08550_ _04205_ _04206_ net653 net793 net1560 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a32o_1
XFILLER_0_134_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09141__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08481_ team_02_WB.instance_to_wrap.top.a1.state\[0\] _04168_ vssd1 vssd1 vccd1 vccd1
+ _04180_ sky130_fd_sc_hd__nand2_2
XANTENNA__14296__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08495__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12809__A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\] net770 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10054__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09033_ net944 _04528_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__nor2_4
XFILLER_0_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11859__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout308_A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09747__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold332 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold343 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold354 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold376 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1217_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net804 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_4
Xfanout812 _04522_ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_8
X_09935_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\] net928 net924 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__a22o_1
Xfanout823 _04514_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_6
XFILLER_0_102_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout834 net836 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__buf_4
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout677_A _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net846 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_6
XANTENNA__13700__B1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout856 net857 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_2
Xfanout867 net869 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_4
X_09866_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\] net778 net720 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__a22o_1
Xfanout878 net881 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_8
Xhold1010 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout889 _04536_ vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_4
Xhold1032 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ net1660 net1041 net990 team_02_WB.instance_to_wrap.ramaddr\[14\] vssd1 vssd1
+ vccd1 vccd1 _02608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1043 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout844_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1054 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ net519 vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__inv_2
Xhold1065 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1087 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ _04302_ net848 _04365_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1098 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08679_ team_02_WB.instance_to_wrap.top.a1.instruction\[4\] _04266_ vssd1 vssd1 vccd1
+ vccd1 _04308_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15932__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10710_ team_02_WB.instance_to_wrap.top.pc\[20\] _06184_ _06226_ vssd1 vssd1 vccd1
+ vccd1 _06227_ sky130_fd_sc_hd__a21o_1
XANTENNA__10293__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ _07140_ _07143_ _07161_ _07175_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10641_ _04272_ _04277_ _04276_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10045__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ team_02_WB.instance_to_wrap.ramload\[22\] net1014 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[22\] sky130_fd_sc_hd__and2_1
XFILLER_0_10_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10572_ net525 net387 vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__nand2_1
XANTENNA__09986__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12311_ net244 net2251 net566 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__mux2_1
XANTENNA__11769__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13291_ _06857_ _02959_ team_02_WB.instance_to_wrap.top.pc\[14\] net1052 vssd1 vssd1
+ vccd1 vccd1 _02995_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08651__B net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15030_ net1206 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09199__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09738__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ net1768 net344 net616 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08946__B1 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12173_ net352 net2639 net464 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11124_ net411 _06631_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13298__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15932_ clknet_leaf_49_wb_clk_i _02072_ _00740_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11055_ _04865_ _05949_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__nor2_1
XANTENNA__15462__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09371__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\] net845 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\]
+ _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__a221o_1
XANTENNA__09910__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15863_ clknet_leaf_14_wb_clk_i _02003_ _00671_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14814_ net1192 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15794_ clknet_leaf_3_wb_clk_i _01934_ _00602_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14745_ net1142 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11957_ net301 net2473 net586 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13470__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10908_ net999 _06422_ _06420_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__o21bai_1
XANTENNA__10284__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14676_ net1075 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ net295 net2276 net489 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16415_ clknet_leaf_66_wb_clk_i _02550_ _01223_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13627_ team_02_WB.instance_to_wrap.top.a1.row1\[12\] _03109_ _03114_ _03177_ vssd1
+ vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__a31o_1
X_10839_ net546 net423 vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__or2_4
XFILLER_0_55_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11233__A1 _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16346_ clknet_leaf_117_wb_clk_i _02486_ _01154_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10036__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ net1049 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] vssd1 vssd1 vccd1
+ vccd1 _03113_ sky130_fd_sc_hd__nor2_2
XFILLER_0_82_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12509_ net244 net2269 net446 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__mux2_1
X_16277_ clknet_leaf_50_wb_clk_i _02417_ _01085_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13489_ team_02_WB.START_ADDR_VAL_REG\[29\] _04260_ vssd1 vssd1 vccd1 vccd1 net213
+ sky130_fd_sc_hd__and2_1
XFILLER_0_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16701__1439 vssd1 vssd1 vccd1 vccd1 net1439 _16701__1439/LO sky130_fd_sc_hd__conb_1
XFILLER_0_67_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09729__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15228_ clknet_leaf_70_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[19\]
+ _00041_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15159_ net1245 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15805__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07981_ _03698_ _03703_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12811__B _04422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\] net920 net808 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\]
+ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a221o_1
XANTENNA__12303__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10612__A team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ net527 _05165_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__nand2_1
X_08602_ net95 net1636 net956 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
X_09582_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\] net768 net732 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08533_ net1046 _04217_ _04218_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08468__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13461__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08736__B team_02_WB.instance_to_wrap.top.a1.instruction\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _06530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10985__C _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11472__A1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10275__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08464_ net1687 net1006 net981 _04165_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08395_ _04095_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11224__A1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire509 _05578_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10027__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09968__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11224__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09016_ net944 _04505_ _04509_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__and3_4
XFILLER_0_66_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold140 team_02_WB.instance_to_wrap.ramaddr\[20\] vssd1 vssd1 vccd1 vccd1 net1598
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 net122 vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold162 team_02_WB.instance_to_wrap.top.a1.row2\[8\] vssd1 vssd1 vccd1 vccd1 net1620
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 net154 vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15485__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold184 net166 vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_02_WB.instance_to_wrap.ramload\[16\] vssd1 vssd1 vccd1 vccd1 net1653
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout642 net644 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_6
X_09918_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\] net772 net720 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout653 _04224_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12213__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 _06111_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_4
Xfanout675 _04412_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13205__A2_N net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout686 _04399_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__buf_6
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout697 _04394_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11337__B _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09849_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\] net825 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12860_ net518 _07378_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11811_ net258 net2534 net590 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _06612_ _06641_ _07314_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__and3_1
X_14530_ net1207 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11742_ net252 net2268 net600 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14461_ net1084 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
X_11673_ _04783_ _06467_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16200_ clknet_leaf_16_wb_clk_i _02340_ _01008_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13412_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _03024_
+ sky130_fd_sc_hd__or3b_1
X_10624_ team_02_WB.instance_to_wrap.top.pc\[28\] _06139_ vssd1 vssd1 vccd1 vccd1
+ _06141_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09959__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input90_A wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14392_ net1196 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16131_ clknet_leaf_125_wb_clk_i _02271_ _00939_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13343_ team_02_WB.instance_to_wrap.ramload\[5\] net1014 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[5\] sky130_fd_sc_hd__and2_1
XFILLER_0_106_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10555_ _04842_ net386 vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16062_ clknet_leaf_112_wb_clk_i _02202_ _00870_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13274_ team_02_WB.instance_to_wrap.ramaddr\[23\] net983 net964 _02986_ vssd1 vssd1
+ vccd1 vccd1 _01442_ sky130_fd_sc_hd__a22o_1
X_10486_ net420 net501 _05738_ _06002_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15013_ net1234 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
XANTENNA__11518__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12225_ net1823 net292 net616 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09592__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ net290 net1767 net464 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
XANTENNA__08601__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ net668 _06612_ _06615_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12123__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ net2420 net278 net583 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
XANTENNA__09344__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11038_ net408 _06403_ _06545_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__a21oi_2
X_15915_ clknet_leaf_115_wb_clk_i _02055_ _00723_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11962__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15846_ clknet_leaf_49_wb_clk_i _01986_ _00654_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ clknet_leaf_117_wb_clk_i _01917_ _00585_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12989_ _07480_ _07508_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11454__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10257__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14728_ net1178 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14659_ net1145 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10009__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11206__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ _03888_ _03893_ _03862_ _03878_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__o211a_2
XFILLER_0_7_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08083__B1 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16329_ clknet_leaf_120_wb_clk_i _02469_ _01137_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput201 net201 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput212 net212 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XANTENNA__12706__A1 team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput223 net223 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09583__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11390__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07964_ _03670_ _03672_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1
+ vccd1 vccd1 _03687_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12033__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09335__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\] net741 net709 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__a22o_1
X_07895_ _03614_ _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14749__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\] net928 net815 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\]
+ _05150_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11693__A1 _07138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09565_ _05061_ _05080_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_84_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10248__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[5\] net980 vssd1 vssd1 vccd1
+ vccd1 _04206_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09496_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\] net776 net760 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\]
+ _05012_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08447_ _04141_ _04146_ _04151_ _04136_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16283__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout807_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08378_ _04081_ _04086_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10340_ net388 vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13828__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10271_ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__inv_2
X_12010_ net243 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\] net477 vssd1
+ vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
XANTENNA__09574__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16795__1339 vssd1 vssd1 vccd1 vccd1 _16795__1339/HI net1339 sky130_fd_sc_hd__conb_1
XFILLER_0_100_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 net453 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09326__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout461 _07220_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout472 _07208_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13961_ net1251 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 net485 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout494 _06252_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11782__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ _07360_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15700_ clknet_leaf_12_wb_clk_i _01840_ _00508_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_16680_ clknet_leaf_73_wb_clk_i _02797_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13892_ net1239 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16700__1438 vssd1 vssd1 vccd1 vccd1 net1438 _16700__1438/LO sky130_fd_sc_hd__conb_1
X_15631_ clknet_leaf_40_wb_clk_i _01771_ _00439_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12843_ _04928_ _06177_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16626__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15562_ clknet_leaf_126_wb_clk_i _01702_ _00370_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10239__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ _06482_ _06517_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_48_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14513_ net1106 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11725_ net317 net2311 net601 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__mux2_1
X_15493_ clknet_leaf_32_wb_clk_i _01633_ _00301_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08852__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13189__A1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14444_ net1071 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
X_11656_ net368 _06287_ _05877_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ _05962_ _06036_ _06121_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__or3_4
X_14375_ net1102 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_135_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12118__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ net378 _06470_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16114_ clknet_leaf_6_wb_clk_i _02254_ _00922_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13326_ _03292_ _03011_ _03010_ team_02_WB.instance_to_wrap.top.a1.hexop\[3\] vssd1
+ vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] sky130_fd_sc_hd__a2bb2o_1
Xhold909 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_111_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10538_ net510 net402 vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16006__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11957__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16045_ clknet_leaf_23_wb_clk_i _02185_ _00853_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ net1579 net985 net966 _02975_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__a22o_1
X_10469_ _05231_ _05251_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12208_ net350 net2045 net580 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13188_ _07084_ net232 net228 _02946_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10175__B2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ net354 net1929 net467 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13113__B2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07680_ _03399_ _03400_ _03402_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__a21o_1
X_16878_ net1422 vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__buf_2
XFILLER_0_126_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15829_ clknet_leaf_41_wb_clk_i _01969_ _00637_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09350_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\] net754 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__a22o_1
XANTENNA__09096__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08301_ _04009_ _04014_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_118_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09281_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\] net763 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\]
+ _04797_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_60_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08232_ _03943_ _03944_ _03946_ _03935_ _03919_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_34_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13222__A1_N net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08163_ _03806_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12028__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ _03801_ _03808_ _03812_ _03814_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_43_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11867__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09556__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13367__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout492_A _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08996_ _04313_ net944 _04507_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__and3_4
XANTENNA__09308__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__A _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07947_ _03641_ _03661_ _03662_ _03663_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__a41o_2
XTAP_TAPCELL_ROW_3_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12698__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15523__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout757_A _04375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07878_ _03574_ _03599_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__xnor2_4
XANTENNA__10800__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09617_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\] net708 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16694__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout924_A _04513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09548_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\] net926 net922 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a22o_1
XANTENNA__09087__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ _04993_ _04995_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_134_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11631__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ _05921_ net658 _05923_ net664 vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12490_ net302 net2326 net558 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16029__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11441_ _05468_ _06009_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14160_ net1099 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
X_11372_ _06870_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11777__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ _07468_ _07469_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nor2_1
X_10323_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\] net893 net885 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\]
+ _05839_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14091_ net1201 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_128_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16179__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09547__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ net229 _02824_ _02825_ _04280_ net1027 vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__a221o_1
XANTENNA_input53_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10254_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\] net688 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__clkbuf_4
Xfanout1212 net1213 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1223 net1224 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_4
X_10185_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\] net821 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__buf_4
X_16801_ net1345 vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_2
Xfanout1245 net1246 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__buf_4
Xfanout1256 net1264 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__clkbuf_4
X_14993_ net1223 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
Xfanout280 net283 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11106__B1 _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout291 _06712_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_2
X_16732_ net1456 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__12401__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13944_ net1236 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
X_13875_ net1261 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
X_16663_ clknet_leaf_101_wb_clk_i _02782_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15614_ clknet_leaf_114_wb_clk_i _01754_ _00422_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12826_ _07346_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__inv_2
XANTENNA__11409__B2 _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09078__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16594_ clknet_leaf_98_wb_clk_i _02713_ _01387_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12757_ _05737_ _05831_ _05909_ _07128_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__or4b_1
X_15545_ clknet_leaf_18_wb_clk_i _01685_ _00353_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08825__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10093__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11708_ net251 net1842 net604 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15476_ clknet_leaf_10_wb_clk_i _01616_ _00284_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12688_ net301 net2729 net431 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08038__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14427_ net1181 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
XANTENNA__13031__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ net947 _07122_ _07125_ net607 vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09786__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14358_ net1094 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09250__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold706 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ team_02_WB.instance_to_wrap.top.pc\[5\] net1051 _07046_ _02960_ vssd1 vssd1
+ vccd1 vccd1 _03004_ sky130_fd_sc_hd__a22o_2
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold728 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold739 team_02_WB.instance_to_wrap.ramload\[10\] vssd1 vssd1 vccd1 vccd1 net2197
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ net1106 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16028_ clknet_leaf_45_wb_clk_i _02168_ _00836_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09002__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15546__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ net1639 net1039 net1035 team_02_WB.instance_to_wrap.ramstore\[14\] vssd1
+ vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XANTENNA__08210__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07801_ _03519_ _03520_ _03492_ _03517_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__and4b_1
X_08781_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\] net758 net730 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07732_ _03423_ _03454_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__nor2_1
XANTENNA__11648__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09710__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10856__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _03384_ _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_66_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09402_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\] net747 net844 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09069__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07594_ net1007 _03317_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__nor2_2
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09333_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\] net814 net911 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\]
+ _04849_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13270__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10766__S net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A _06424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16794__1338 vssd1 vssd1 vccd1 vccd1 _16794__1338/HI net1338 sky130_fd_sc_hd__conb_1
XFILLER_0_30_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09264_ net538 _04776_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08215_ _03902_ _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13022__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09195_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\] net766 _04709_ _04710_
+ _04711_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_69_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08146_ _03833_ _03863_ _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__o21ba_1
XANTENNA__16321__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09241__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08077_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _03762_ _03787_ vssd1 vssd1
+ vccd1 vccd1 _03798_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09529__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13325__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout874_A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__B1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16471__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold11 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[2\] vssd1 vssd1 vccd1 vccd1
+ net1469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold22 _02577_ vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold33 team_02_WB.instance_to_wrap.top.a1.hexop\[4\] vssd1 vssd1 vccd1 vccd1 net1491
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ net1062 net1060 _04267_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__a21o_1
Xhold44 team_02_WB.instance_to_wrap.top.a1.row1\[106\] vssd1 vssd1 vccd1 vccd1 net1502
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13089__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 team_02_WB.instance_to_wrap.top.a1.row1\[107\] vssd1 vssd1 vccd1 vccd1 net1513
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 _02583_ vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_02_WB.START_ADDR_VAL_REG\[8\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12221__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold88 net121 vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net292 net1920 net478 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__mux2_1
Xhold99 net161 vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09701__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11345__B _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ _04694_ net660 _04695_ net665 vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_85_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13660_ _04125_ net851 _03197_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__a21oi_1
X_10872_ _06386_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ net1724 net250 net554 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13261__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13591_ team_02_WB.instance_to_wrap.top.a1.row1\[9\] _03110_ _03111_ team_02_WB.instance_to_wrap.top.a1.row1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__a22o_1
XANTENNA__08807__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15330_ clknet_leaf_63_wb_clk_i _01473_ _00143_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10075__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12542_ net246 net2706 net444 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15261_ clknet_leaf_59_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[20\]
+ _00074_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12473_ net345 net2255 net450 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14212_ net1132 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
XANTENNA__09768__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11424_ _06819_ _06920_ net397 vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15192_ net1249 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
XANTENNA__08670__A team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09232__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_8 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14143_ net1183 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11355_ _05295_ _06111_ net656 _06854_ _06846_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_39_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13316__B2 _03007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\] net780 net768 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__a22o_1
X_14074_ net1186 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
X_11286_ _06190_ net655 _06788_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13025_ _06368_ net233 vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ _05747_ _05749_ _05751_ _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1020 net1022 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1031 _04429_ vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_4
Xfanout1042 net1043 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09940__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10168_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\] net941 net893 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a22o_1
Xfanout1053 net1054 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_98_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1075 net1079 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_4
Xfanout1086 net1088 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__buf_4
XANTENNA__12131__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1097 net1199 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10440__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09299__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10099_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\] net680 _05605_ _05608_
+ _05615_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a2111o_1
X_14976_ net1245 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_63_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16715_ net1274 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_88_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13927_ net1204 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14847__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11970__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16646_ clknet_leaf_100_wb_clk_i _02765_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13858_ net1226 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12809_ net791 _07332_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__nand2_1
X_16577_ clknet_leaf_95_wb_clk_i _00003_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13789_ _03278_ _03279_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15528_ clknet_leaf_16_wb_clk_i _01668_ _00336_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16344__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09471__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15459_ clknet_leaf_125_wb_clk_i _01599_ _00267_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08000_ _03689_ net255 vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__nand2_1
XANTENNA__09759__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09223__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold503 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16494__CLK clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold514 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12306__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold525 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13307__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _05465_ _05466_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__nor2_2
Xhold558 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08902_ net2 net1029 net987 net1731 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09882_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\] net726 _05391_ _05392_
+ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12830__A _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08833_ net163 net1039 net1035 net1561 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__a22o_1
XANTENNA__09931__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1203 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1214 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1236 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\] vssd1
+ vssd1 vccd1 vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\] net718 _04390_ _04392_
+ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a211o_1
XANTENNA__12041__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1258 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
X_07715_ _03408_ net425 _03403_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__and3b_1
X_08695_ net1058 _03298_ _04271_ _04318_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout455_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1197_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07646_ _03363_ _03368_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07577_ net2738 net188 _00017_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\] net718 _04829_ _04830_
+ _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10057__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09462__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ _04757_ _04759_ _04761_ _04763_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09178_ _04693_ _04694_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__nand2b_2
XANTENNA__09214__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout991_A _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12724__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ _03829_ _03836_ _03837_ _03848_ _03807_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_31_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12216__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__A _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11140_ _04470_ _06627_ _06647_ net670 _06646_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__o221a_2
XANTENNA__15861__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__B _05760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _04865_ _06110_ net662 _04863_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__a22o_1
Xinput101 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_1
X_10022_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\] net912 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a22o_1
XANTENNA__13053__A1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16217__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830_ net1163 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11973_ net344 net2188 net585 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__mux2_1
XANTENNA__08489__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ net1100 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11790__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16500_ clknet_leaf_6_wb_clk_i _02634_ _01307_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10296__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10924_ _06432_ _06437_ net414 vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__mux2_1
X_13712_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] _03227_ net1670 vssd1
+ vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14692_ net1126 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16367__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16431_ clknet_leaf_103_wb_clk_i net1693 _01239_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13234__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ net975 _06366_ _06369_ _06370_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__a211o_1
X_13643_ team_02_WB.instance_to_wrap.top.a1.row1\[111\] _03160_ _03161_ _03190_ vssd1
+ vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10048__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09989__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16362_ clknet_leaf_129_wb_clk_i _02502_ _01170_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ team_02_WB.instance_to_wrap.top.a1.row2\[8\] _03122_ _03126_ team_02_WB.instance_to_wrap.top.a1.row2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a22o_1
X_10786_ _06300_ _06301_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15313_ clknet_leaf_64_wb_clk_i _01456_ _00126_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12525_ net297 net2329 net447 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__mux2_1
XANTENNA__15391__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16293_ clknet_leaf_32_wb_clk_i _02433_ _01101_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15244_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[3\]
+ _00057_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_12456_ net293 net2236 net451 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__mux2_1
XANTENNA__08604__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09205__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11407_ _05381_ _06110_ _06901_ _06104_ _06904_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15175_ net1250 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12387_ net291 net1903 net460 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__mux2_1
XANTENNA__12126__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ net1096 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
X_11338_ net974 _06212_ _06831_ _06838_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11965__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ net1109 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
X_11269_ _06714_ _06771_ net371 vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13008_ _07457_ _07527_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16793__1337 vssd1 vssd1 vccd1 vccd1 _16793__1337/HI net1337 sky130_fd_sc_hd__conb_1
XFILLER_0_24_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14959_ net1115 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13473__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10287__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08480_ net1063 _04170_ _04173_ net959 vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__o211a_1
XANTENNA__12809__B _07332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16629_ clknet_leaf_100_wb_clk_i _02748_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13225__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09444__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09101_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\] net766 net843 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\]
+ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13420__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09032_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\] net831 net905 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08514__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12036__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold311 team_02_WB.instance_to_wrap.top.a1.row1\[12\] vssd1 vssd1 vccd1 vccd1 net1769
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold322 team_02_WB.instance_to_wrap.top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1 net1780
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold333 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold344 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold366 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11875__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net804 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
XFILLER_0_110_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09934_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\] net807 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\]
+ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__a221o_1
Xhold399 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout813 _04521_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_6
XFILLER_0_102_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1112_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout824 _04514_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_8
Xfanout846 _04400_ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_4
XANTENNA__09904__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout857 _04550_ vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__buf_8
X_09865_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\] net730 net714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__a22o_1
Xhold1000 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout572_A _07217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 net869 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_6
Xfanout879 net881 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_4
Xhold1011 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08816_ net1647 net1042 net992 team_02_WB.instance_to_wrap.ramaddr\[15\] vssd1 vssd1
+ vccd1 vccd1 _02609_ sky130_fd_sc_hd__a22o_1
Xhold1033 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1044 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ _05306_ _05308_ _05310_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nor4_1
XFILLER_0_119_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1055 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net847 _04363_ _04368_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__and3_4
Xhold1088 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout837_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08678_ _04305_ _04285_ _04290_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__or3b_1
XANTENNA__09683__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07629_ _03349_ _03350_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__nand2_1
XANTENNA__13216__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ _04277_ net1057 net1059 vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09435__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10571_ net424 net412 vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12310_ net242 net1989 net568 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15111__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13290_ team_02_WB.instance_to_wrap.ramaddr\[15\] net985 net966 _02994_ vssd1 vssd1
+ vccd1 vccd1 _01434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12241_ net1717 net349 net618 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10202__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12172_ net357 net1766 net462 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11785__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net398 _06630_ _06628_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15607__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07564__A team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11054_ net2174 net267 net641 vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__mux2_1
X_15931_ clknet_leaf_125_wb_clk_i _02071_ _00739_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10702__B _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10005_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\] net744 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15862_ clknet_leaf_62_wb_clk_i _02002_ _00670_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14813_ net1081 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15793_ clknet_leaf_51_wb_clk_i _01933_ _00601_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15757__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10269__A0 _05740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14744_ net1196 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11956_ net294 net1969 net587 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__mux2_1
XANTENNA__09674__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10907_ _06271_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14675_ net1166 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
X_11887_ net284 net2716 net487 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16414_ clknet_leaf_67_wb_clk_i _02549_ _01222_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10838_ _06348_ _06352_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nand2_1
X_13626_ net1047 net1050 team_02_WB.instance_to_wrap.top.a1.row2\[12\] _03103_ vssd1
+ vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09426__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16345_ clknet_leaf_17_wb_clk_i _02485_ _01153_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10769_ _05877_ net385 vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nor2_1
X_13557_ _03289_ net1048 vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12508_ net242 net2498 net448 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__mux2_1
X_13488_ team_02_WB.START_ADDR_VAL_REG\[28\] net1070 net1003 vssd1 vssd1 vccd1 vccd1
+ net212 sky130_fd_sc_hd__a21o_1
X_16276_ clknet_leaf_11_wb_clk_i _02416_ _01084_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15227_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[18\]
+ _00040_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_12439_ net349 net2158 net456 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15158_ net1246 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14109_ net1081 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
X_07980_ _03670_ _03700_ _03702_ _03698_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__a22o_1
X_15089_ net1078 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15287__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire540_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13694__B1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09650_ net527 _05165_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08601_ net96 net1595 net956 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09581_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\] net736 net712 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__a22o_1
X_08532_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[1\] net980 vssd1 vssd1 vccd1
+ vccd1 _04218_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09665__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08463_ _04154_ _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08394_ _04090_ _04093_ _04099_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_114_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09417__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout320_A _06936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout418_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10983__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09015_ net1056 _04297_ _04313_ net951 vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__and4b_1
XFILLER_0_116_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16062__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12185__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold130 team_02_WB.instance_to_wrap.top.a1.row1\[1\] vssd1 vssd1 vccd1 vccd1 net1588
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold141 _02614_ vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _02618_ vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__A0 _07013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold163 team_02_WB.instance_to_wrap.top.a1.row1\[104\] vssd1 vssd1 vccd1 vccd1 net1621
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _02585_ vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _02567_ vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold196 team_02_WB.instance_to_wrap.top.a1.row1\[0\] vssd1 vssd1 vccd1 vccd1 net1654
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09917_ _05422_ _05426_ _05430_ _05433_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout643 net644 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_8
XANTENNA__16697__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_2
XANTENNA_fanout954_A _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout665 _06111_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_2
Xfanout676 _04412_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout687 _04399_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_4
X_09848_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\] net805 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\]
+ _05364_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__a221o_1
Xfanout698 net701 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\] net718 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ net248 net2418 net589 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _06698_ _06671_ _06670_ _06669_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__and4b_1
XFILLER_0_95_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09656__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ net239 net2525 net597 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14460_ net1146 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
X_11672_ _04695_ _07157_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09408__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__A _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10623_ _06139_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__inv_2
X_13411_ _03018_ _03020_ _03021_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__or4_4
XFILLER_0_3_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14391_ net1172 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16792__1336 vssd1 vssd1 vccd1 vccd1 _16792__1336/HI net1336 sky130_fd_sc_hd__conb_1
XFILLER_0_91_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13342_ team_02_WB.instance_to_wrap.ramload\[4\] net1014 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[4\] sky130_fd_sc_hd__and2_1
X_16130_ clknet_leaf_122_wb_clk_i _02270_ _00938_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10554_ _06070_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input83_A wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10974__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16061_ clknet_leaf_52_wb_clk_i _02201_ _00869_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13273_ team_02_WB.instance_to_wrap.top.pc\[23\] net1052 _06618_ net935 vssd1 vssd1
+ vccd1 vccd1 _02986_ sky130_fd_sc_hd__a22o_1
X_10485_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15012_ net1233 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
X_12224_ net2734 net286 net618 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__mux2_1
XANTENNA__09774__A _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10726__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ net276 net2034 net463 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12404__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11106_ _05983_ net665 _06117_ _06613_ _06614_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__o221a_1
X_12086_ net2018 net282 net583 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
XANTENNA__11528__B _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15914_ clknet_leaf_130_wb_clk_i _02054_ _00722_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11037_ net423 _06547_ _06357_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15845_ clknet_leaf_32_wb_clk_i _01985_ _00653_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ clknet_leaf_113_wb_clk_i _01916_ _00584_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ team_02_WB.instance_to_wrap.top.pc\[9\] _05537_ _07507_ vssd1 vssd1 vccd1
+ vccd1 _07508_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_103_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14727_ net1101 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08855__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11939_ net344 net1958 net482 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09949__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14658_ net1205 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16085__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13609_ _03112_ _03127_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nor2_1
XANTENNA__11206__A2 _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14589_ net1085 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16328_ clknet_leaf_14_wb_clk_i _02468_ _01136_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09280__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16259_ clknet_leaf_13_wb_clk_i _02399_ _01067_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput202 net202 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput213 net213 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XANTENNA__09032__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11914__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15922__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12314__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10623__A _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11390__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07963_ _03651_ _03685_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_71_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10455__A_N _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09702_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\] net757 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\]
+ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13131__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07894_ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09886__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\] net827 net924 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a22o_1
XANTENNA__16667__D _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12890__A1 _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout270_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09564_ _05061_ _05080_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09099__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ team_02_WB.instance_to_wrap.top.a1.data\[5\] net958 vssd1 vssd1 vccd1 vccd1
+ _04205_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09495_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\] net704 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a22o_1
XANTENNA__16428__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14765__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08446_ _04130_ _04139_ _04142_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08377_ _04081_ _04084_ _04085_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout702_A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09271__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09810__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10270_ net792 _04492_ _05786_ net652 vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12224__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10184__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout440 net441 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_6
XFILLER_0_100_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout451 net453 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_4
Xfanout462 net465 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout473 _07208_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13960_ net1238 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
Xfanout484 net485 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_8
Xfanout495 _06252_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09877__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12911_ _07361_ _07430_ _07362_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_31_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13891_ net1253 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15630_ clknet_leaf_25_wb_clk_i _01770_ _00438_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12842_ _04494_ _04886_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__or2_1
XANTENNA__09629__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12633__A1 _07051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15561_ clknet_leaf_104_wb_clk_i _01701_ _00369_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08837__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12773_ net546 _06118_ _06402_ _07296_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__and4_1
XFILLER_0_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ net1095 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11724_ net313 net2447 net601 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15492_ clknet_leaf_2_wb_clk_i _01632_ _00300_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14443_ net1203 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
X_11655_ _05649_ _05922_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10606_ _04461_ _06114_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_88_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11586_ _05910_ _06000_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__xor2_1
X_14374_ net1073 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09801__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16113_ clknet_leaf_21_wb_clk_i _02253_ _00921_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10537_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_17_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13325_ net1641 _03010_ _03012_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ clknet_leaf_25_wb_clk_i _02184_ _00852_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13256_ team_02_WB.instance_to_wrap.top.pc\[29\] net1054 net935 _02974_ vssd1 vssd1
+ vccd1 vccd1 _02975_ sky130_fd_sc_hd__a22o_1
X_10468_ _05212_ _05977_ _05980_ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__or4_1
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ net362 net2244 net579 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__mux2_1
XANTENNA__12134__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ _07495_ _07498_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__xor2_1
X_10399_ _05691_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__nor2_2
XFILLER_0_104_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12849__A_N _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12138_ net359 net2422 net466 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11973__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12069_ net339 net2279 net473 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09868__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16877_ net1421 vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__buf_2
XFILLER_0_35_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15828_ clknet_leaf_12_wb_clk_i _01968_ _00636_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire503_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15759_ clknet_leaf_36_wb_clk_i _01899_ _00567_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12624__A1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08828__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08300_ _03985_ _04010_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__xnor2_1
X_09280_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\] net731 net715 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08231_ _03947_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08162_ _03840_ _03847_ _03859_ _03841_ _03802_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_1675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09253__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08093_ _03759_ _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12833__A _04631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08522__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08359__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13219__A2_N net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10166__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08995_ net943 _04503_ _04505_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__and3_1
XANTENNA__11883__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ _03666_ _03668_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11115__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16791__1335 vssd1 vssd1 vccd1 vccd1 _16791__1335/HI net1335 sky130_fd_sc_hd__conb_1
XFILLER_0_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ _03574_ _03599_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16250__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09616_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\] net768 _05130_ _05132_
+ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08819__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\] net833 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\]
+ _05063_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__a221o_1
XANTENNA__14495__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout917_A _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ _04970_ _04991_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08429_ _04128_ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_43_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12219__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11440_ net2351 net317 net642 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09244__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11051__B1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _06772_ _06869_ net397 vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13110_ _07371_ _07419_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__nor2_1
X_10322_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\] net925 net881 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14090_ net1168 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13041_ _07355_ _07437_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_128_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10253_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\] net748 _05767_ _05768_
+ _05769_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_128_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10157__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input46_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\] net801 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\]
+ _05700_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__a221o_1
Xfanout1202 net1212 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1213 net1265 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_33_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1224 net1225 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11793__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16800_ net1344 vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_2
Xfanout1235 net1237 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_4
Xfanout1246 net1250 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__clkbuf_4
X_14992_ net1221 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
Xfanout1257 net1260 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_4
XANTENNA__08668__A team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout281 net283 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16731_ net1455 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
Xfanout292 _06791_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
X_13943_ net1236 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16662_ clknet_leaf_101_wb_clk_i _02781_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13874_ net1259 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15613_ clknet_leaf_49_wb_clk_i _01753_ _00421_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12825_ _03319_ _07340_ _07341_ _04172_ _03317_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__o32a_1
X_16593_ clknet_leaf_96_wb_clk_i _02712_ _01386_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15544_ clknet_leaf_53_wb_clk_i _01684_ _00352_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12756_ _05647_ _05691_ _07278_ _07279_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__or4_1
XANTENNA__08607__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ net237 net2569 net601 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
X_15475_ clknet_leaf_56_wb_clk_i _01615_ _00283_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12129__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ net292 net2265 net432 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14426_ net1182 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11638_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] _04347_ net953 _07124_ vssd1
+ vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11968__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14357_ net1187 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ net417 _06694_ _06898_ net375 _07055_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__a221o_2
XFILLER_0_53_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold707 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13308_ net2397 net984 net965 _03003_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16123__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold718 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold729 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ net1113 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16027_ clknet_leaf_127_wb_clk_i _02167_ _00835_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13239_ _02953_ _02958_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__nand2_1
XANTENNA__10148__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09002__A3 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16273__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ _03515_ _03522_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__nand2b_2
XANTENNA__08761__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08780_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\] net770 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\]
+ _04408_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10901__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07731_ _03386_ _03411_ _03418_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10620__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07662_ _03347_ _03379_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_66_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10320__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\] net751 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07593_ team_02_WB.instance_to_wrap.top.a1.state\[1\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ _03317_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_62_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09332_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\] net899 net887 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09474__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09263_ _04779_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12039__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout233_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08214_ _03901_ _03921_ _03927_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09226__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09194_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\] net730 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11878__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08145_ _03829_ _03836_ net226 vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout400_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__A1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08076_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _03787_ _03762_ vssd1 vssd1
+ vccd1 vccd1 _03797_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10139__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__A1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout867_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold12 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[7\] vssd1 vssd1 vccd1 vccd1
+ net1470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_02_WB.instance_to_wrap.ramstore\[30\] vssd1 vssd1 vccd1 vccd1 net1481
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12502__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ net1062 net1060 _04267_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__a21oi_1
Xhold34 team_02_WB.instance_to_wrap.top.a1.nextHex\[3\] vssd1 vssd1 vccd1 vccd1 net1492
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 net127 vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15640__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold56 team_02_WB.instance_to_wrap.top.a1.data\[9\] vssd1 vssd1 vccd1 vccd1 net1514
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_02_WB.instance_to_wrap.ramstore\[10\] vssd1 vssd1 vccd1 vccd1 net1525
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] _03648_ _03649_ _03650_ vssd1
+ vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__o211a_1
XANTENNA__11639__A2 _07122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold78 team_02_WB.instance_to_wrap.top.a1.row1\[114\] vssd1 vssd1 vccd1 vccd1 net1536
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold89 _02617_ vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11118__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10940_ _06355_ _06452_ net657 vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10871_ _06384_ _06385_ net401 vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12610_ net2096 net253 net555 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11642__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input100_A wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ team_02_WB.instance_to_wrap.top.a1.row2\[41\] _03123_ _03125_ team_02_WB.instance_to_wrap.top.a1.row2\[33\]
+ _03143_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a221o_1
XANTENNA__09465__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13261__B2 _02978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12541_ net242 net2536 net445 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15260_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[19\]
+ _00073_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12472_ net348 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\] net453 vssd1
+ vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08951__A _04463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11788__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14211_ net1131 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
X_11423_ _06868_ _06919_ net367 vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15191_ net1248 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08670__B team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10378__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14142_ net1189 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07567__A team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11354_ _06354_ _06853_ _06850_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_39_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10705__B _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16296__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\] net716 _05820_ _05821_
+ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__a211o_1
XANTENNA__13316__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11285_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] net494 _06787_ _04263_ net496
+ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__a221o_1
X_14073_ net1140 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13024_ net1027 _07543_ net1025 team_02_WB.instance_to_wrap.top.pc\[31\] vssd1 vssd1
+ vccd1 vccd1 _01512_ sky130_fd_sc_hd__a2bb2o_1
X_10236_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\] net803 net799 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\]
+ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_89_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1010 _03014_ vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1021 net1022 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__buf_1
XFILLER_0_105_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1032 _04429_ vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__dlymetal6s2s_1
X_10167_ _05677_ _05679_ _05681_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__or4_1
XANTENNA__12412__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__buf_4
Xfanout1054 team_02_WB.instance_to_wrap.top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1054 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1065 _00018_ vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_2
XANTENNA__13221__A1_N net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1076 net1077 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__buf_4
X_10098_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\] net716 _05612_ _05613_
+ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__a2111o_1
Xfanout1087 net1088 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_4
X_14975_ net1247 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
Xfanout1098 net1103 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_4
X_16714_ net1273 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_117_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13926_ net1203 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10302__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16645_ clknet_leaf_99_wb_clk_i _02764_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13857_ net1226 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15024__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ _07330_ _07331_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__and2b_2
X_16576_ clknet_leaf_99_wb_clk_i _00002_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09456__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13788_ net2432 _03276_ net960 vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15527_ clknet_leaf_32_wb_clk_i _01667_ _00335_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_32_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12739_ net796 _06108_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15458_ clknet_leaf_122_wb_clk_i _01598_ _00266_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16790__1334 vssd1 vssd1 vccd1 vccd1 _16790__1334/HI net1334 sky130_fd_sc_hd__conb_1
X_14409_ net1100 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15513__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15389_ clknet_leaf_50_wb_clk_i _01529_ _00197_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10369__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold504 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold515 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10615__B _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13307__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold548 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09950_ _05466_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold559 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08901_ net13 net1031 net989 net2067 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a22o_1
XANTENNA__15663__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09692__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\] net710 _05394_ _05395_
+ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12830__B _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08832_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] _03301_ team_02_WB.instance_to_wrap.wb.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__and3b_4
XANTENNA__12322__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1204 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1215 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1237 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\] net722 net698 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__a22o_1
Xhold1259 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07714_ _03431_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13942__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08694_ net1061 _04309_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__nor2_1
X_07645_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] _03364_ _03365_ _03366_ vssd1
+ vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_95_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1092_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout448_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ team_02_WB.instance_to_wrap.top.pad.count\[1\] team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__and2b_1
XFILLER_0_48_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09447__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09315_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\] net783 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\]
+ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold1298_A team_02_WB.instance_to_wrap.ramstore\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_119_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\] net830 net814 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\]
+ _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13389__A team_02_WB.instance_to_wrap.ramload\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09177_ _04656_ _04661_ _04671_ _04692_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__or4_4
XFILLER_0_50_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08490__B _04177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08128_ _03846_ _03847_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10765__C1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout984_A _02956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08059_ _03736_ _03777_ _03778_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_43_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11070_ net379 _06579_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput102 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
X_10021_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\] net896 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__a22o_1
XANTENNA__15109__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08725__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14760_ net1177 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09686__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ net349 net1890 net588 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09150__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ net2508 _03227_ _03229_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10923_ _06436_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14691_ net1134 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16430_ clknet_leaf_103_wb_clk_i net1619 _01238_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13642_ team_02_WB.instance_to_wrap.top.a1.row1\[15\] _03113_ _03109_ vssd1 vssd1
+ vccd1 vccd1 _03190_ sky130_fd_sc_hd__o21a_1
X_10854_ _06131_ net655 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[30\] net497
+ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16361_ clknet_leaf_104_wb_clk_i _02501_ _01169_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13573_ _03107_ _03127_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__nor2_2
XFILLER_0_137_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10785_ _05440_ net402 vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15312_ clknet_leaf_103_wb_clk_i _01455_ _00125_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12524_ net308 net1813 net447 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16292_ clknet_leaf_3_wb_clk_i _02432_ _01100_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15243_ clknet_leaf_63_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[2\]
+ _00056_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12455_ net286 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\] net452 vssd1
+ vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12407__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15686__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11406_ _05378_ net661 net658 _05379_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15174_ net1241 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12386_ net276 net2058 net458 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08964__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14125_ net1154 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11337_ _06836_ _06837_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14056_ net1175 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
X_11268_ _05103_ net387 _06089_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__o21ai_1
X_13007_ _07458_ _07526_ _07459_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_24_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10219_ net422 net501 vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__nor2_1
XANTENNA__12142__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11199_ _04469_ _06687_ _06704_ net672 _06703_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__a221o_1
XANTENNA__10451__A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11981__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14958_ net1163 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09677__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16311__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13175__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09141__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ net1222 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
X_14889_ net1109 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16628_ clknet_leaf_100_wb_clk_i _02747_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13225__B2 _05602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10039__A1 _05555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16559_ clknet_leaf_93_wb_clk_i _02683_ _01366_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14593__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08101__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09100_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\] net682 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08591__A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09031_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\] net819 net869 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12317__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11539__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13113__A1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold301 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold312 _02696_ vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold323 team_02_WB.instance_to_wrap.top.a1.row1\[10\] vssd1 vssd1 vccd1 vccd1 net1781
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold334 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold367 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09933_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\] net904 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a22o_1
Xfanout803 net804 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_6
XANTENNA__08530__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout814 _04521_ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_4
Xfanout825 net828 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout398_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout836 _04506_ vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout847 _04359_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__buf_2
X_09864_ _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__inv_2
XANTENNA__12052__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout858 net861 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_8
XANTENNA__15409__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1105_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 _04541_ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_4
Xhold1012 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ net1544 net1041 net990 team_02_WB.instance_to_wrap.ramaddr\[16\] vssd1 vssd1
+ vccd1 vccd1 _02610_ sky130_fd_sc_hd__a22o_1
Xhold1023 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\] net738 net714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\]
+ _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a221o_1
Xhold1034 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11891__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout565_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1056 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ _04302_ net847 _04365_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__and3_4
XFILLER_0_9_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1078 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09668__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1089 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08677_ _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout732_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07628_ team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] _03348_ vssd1 vssd1 vccd1
+ vccd1 _03351_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13216__B2 _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07559_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[3\] vssd1 vssd1 vccd1 vccd1
+ _03300_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10570_ net419 net413 vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09840__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\] net844 _04740_ _04742_
+ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_23_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12227__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09199__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ net1798 net361 net619 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__mux2_1
X_12171_ net342 net2425 net465 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__mux2_1
XANTENNA__13847__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11122_ _06576_ _06629_ net370 vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold890 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13152__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11053_ net947 _06556_ _06563_ net607 vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__o211a_2
X_15930_ clknet_leaf_119_wb_clk_i _02070_ _00738_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10004_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\] net788 net732 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09371__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ clknet_leaf_43_wb_clk_i _02001_ _00669_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14812_ net1149 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
X_15792_ clknet_leaf_33_wb_clk_i _01932_ _00600_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09659__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10269__A1 _05785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14743_ net1124 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11955_ net284 net1994 net587 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__mux2_1
XANTENNA__16484__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output115_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ team_02_WB.instance_to_wrap.top.pc\[29\] _06270_ vssd1 vssd1 vccd1 vccd1
+ _06421_ sky130_fd_sc_hd__nor2_1
X_14674_ net1123 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11886_ net274 net2687 net486 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16413_ clknet_leaf_67_wb_clk_i _02548_ _01221_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13625_ net1522 net963 _03176_ net1067 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10837_ _06352_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16344_ clknet_leaf_51_wb_clk_i _02484_ _01152_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13556_ net1049 _03290_ _03109_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__and3_1
XANTENNA__08615__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ _04611_ _06033_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__xor2_1
XFILLER_0_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12507_ net645 _07203_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12137__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16275_ clknet_leaf_85_wb_clk_i _02415_ _01083_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13487_ team_02_WB.START_ADDR_VAL_REG\[27\] net1068 net1002 vssd1 vssd1 vccd1 vccd1
+ net211 sky130_fd_sc_hd__a21o_1
XFILLER_0_54_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10446__A _04464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10699_ team_02_WB.instance_to_wrap.top.pc\[17\] _06190_ vssd1 vssd1 vccd1 vccd1
+ _06216_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15226_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[17\]
+ _00039_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_125_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12438_ net361 net1991 net455 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15157_ net1243 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12369_ net341 net2281 net564 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14108_ net1150 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
X_15088_ net1078 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ net1121 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire533_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09362__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15701__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ _04249_ _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__nand2_2
XANTENNA__12600__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09580_ _05085_ _05089_ _05093_ _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11457__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ team_02_WB.instance_to_wrap.top.a1.data\[1\] net959 vssd1 vssd1 vccd1 vccd1
+ _04217_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08462_ _04158_ _04160_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1
+ vccd1 vccd1 _04164_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16885__1429 vssd1 vssd1 vccd1 vccd1 _16885__1429/HI net1429 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08393_ _04082_ _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12836__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09822__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16207__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12047__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09014_ _04297_ _04313_ _04500_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11886__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold120 team_02_WB.START_ADDR_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08928__A2 _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold131 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1
+ net1589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 net129 vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 net132 vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15231__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11932__A1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16357__CLK clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 net110 vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold175 team_02_WB.instance_to_wrap.ramaddr\[1\] vssd1 vssd1 vccd1 vccd1 net1633
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1
+ net1644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout682_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout600 _07191_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_4
Xhold197 team_02_WB.instance_to_wrap.top.a1.row2\[1\] vssd1 vssd1 vccd1 vccd1 net1655
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09916_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\] net780 _05431_ _05432_
+ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout644 _04454_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_4
XANTENNA__09889__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout655 _06247_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_4
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_2
XANTENNA__09353__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout677 _04412_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09847_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\] net906 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__a22o_1
Xfanout688 _04399_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout699 net701 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_4
XANTENNA_fanout947_A _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14498__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12510__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09778_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] net931 vssd1 vssd1 vccd1
+ vccd1 _04358_ sky130_fd_sc_hd__and2_1
XANTENNA__11448__B1 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11740_ net246 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\] net597 vssd1
+ vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__mux2_1
XANTENNA__10120__B1 _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10671__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ _04569_ _04611_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__and2b_1
XANTENNA__08943__B _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__or4b_1
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10622_ net552 _06128_ _06138_ _06126_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__a31o_2
X_14390_ net1095 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09813__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ net2393 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[3\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10553_ _06054_ _06069_ net413 vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__mux2_2
XFILLER_0_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10266__A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10974__A2 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16060_ clknet_leaf_45_wb_clk_i _02200_ _00868_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13272_ net1682 net985 net966 _02985_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a22o_1
XANTENNA_input76_A wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10484_ _05907_ _06000_ _05908_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15011_ net1233 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11796__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ net2209 net274 net616 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10187__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ net280 net2532 net463 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__mux2_1
XANTENNA__09592__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11105_ _04907_ _06113_ _06116_ _04908_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12085_ net2115 net269 net583 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
XANTENNA__09344__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15913_ clknet_leaf_104_wb_clk_i _02053_ _00721_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11036_ net410 _06546_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__nor2_1
X_16893_ net1437 vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__buf_2
XFILLER_0_95_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15844_ clknet_leaf_1_wb_clk_i _01984_ _00652_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12420__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15775_ clknet_leaf_109_wb_clk_i _01915_ _00583_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _07505_ _07506_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_103_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08304__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ net1072 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10111__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__A1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11938_ net350 net1960 net485 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14657_ net1210 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
X_11869_ net360 net2035 net492 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13608_ _03115_ _03120_ _03116_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__a21o_1
X_14588_ net1149 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
XANTENNA__09804__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16327_ clknet_leaf_24_wb_clk_i _02467_ _01135_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13539_ team_02_WB.instance_to_wrap.top.edg2.button_i _03074_ _03083_ _03087_ vssd1
+ vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14871__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15254__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16258_ clknet_leaf_125_wb_clk_i _02398_ _01066_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15209_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[0\]
+ _00022_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput203 net203 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16189_ clknet_leaf_52_wb_clk_i _02329_ _00997_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput214 net214 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10904__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09583__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07962_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] _03648_ _03670_ _03672_ vssd1
+ vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_71_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09701_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\] net775 net773 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__a22o_1
XANTENNA__09335__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07893_ _03580_ _03606_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\] net805 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\]
+ _05148_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__a221o_1
XANTENNA__12330__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09563_ net971 net631 net543 vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_77_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout263_A _06595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16739__1284 vssd1 vssd1 vccd1 vccd1 _16739__1284/HI net1284 sky130_fd_sc_hd__conb_1
XFILLER_0_37_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13950__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ _04204_ net1781 net850 vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10102__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\] net752 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\]
+ _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10653__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08445_ _04141_ _04146_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout430_A _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1172_A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08376_ net1700 net1005 net981 _04086_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08074__A2 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15747__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12505__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__A _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09574__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08782__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 _07229_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_126_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout441 _07226_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15897__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09326__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_8
Xfanout463 net465 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout474 _07206_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout485 _07200_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12910_ _04928_ _06177_ _07429_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__a21o_1
Xfanout496 _06250_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15117__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12240__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ net1251 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
XANTENNA__10341__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12841_ _04494_ _04886_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__and2_1
XANTENNA__14956__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15560_ clknet_leaf_19_wb_clk_i _01700_ _00368_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12772_ _06579_ _06606_ net379 vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14511_ net1113 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ net307 net1931 net601 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ clknet_leaf_116_wb_clk_i _01631_ _00299_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14442_ net1139 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11654_ _05468_ _07139_ _06011_ _06956_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_71_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10708__B _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10605_ _04461_ _06114_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__nor2_2
XFILLER_0_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14373_ net1094 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14691__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11585_ net417 _06726_ _06921_ net375 _07073_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__a221o_2
XFILLER_0_49_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16112_ clknet_leaf_39_wb_clk_i _02252_ _00920_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13324_ _04169_ _03010_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_94_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _06044_ _06052_ net396 vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16043_ clknet_leaf_117_wb_clk_i _02183_ _00851_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13255_ _02965_ _02973_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12415__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ _04951_ _05983_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12206_ net352 net2699 net579 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_57_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13186_ _07389_ _07393_ _07394_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10398_ net505 _05690_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__and2_1
X_16884__1428 vssd1 vssd1 vccd1 vccd1 _16884__1428/HI net1428 sky130_fd_sc_hd__conb_1
X_12137_ net341 net2709 net468 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09317__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12068_ net331 net1970 net472 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11019_ net2110 net258 net641 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__mux2_1
XANTENNA__12150__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10332__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16876_ net1420 vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__buf_2
XFILLER_0_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15827_ clknet_leaf_55_wb_clk_i _01967_ _00635_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15758_ clknet_leaf_9_wb_clk_i _01898_ _00566_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ net1215 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15689_ clknet_leaf_118_wb_clk_i _01829_ _00497_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08230_ _03935_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_60_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10618__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08161_ _03840_ _03847_ net226 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08092_ _03771_ _03776_ _03781_ _03787_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12833__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12325__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09556__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08104__A team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11362__A1_N net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ net944 _04507_ _04509_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__and3_4
XANTENNA__09308__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _03626_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__xor2_2
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout478_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12060__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ net316 _03597_ _03586_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10323__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\] net720 net704 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\]
+ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09546_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\] net870 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08774__A team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16545__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ _04970_ _04992_ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_138_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10809__A _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08428_ net1743 net1005 net981 _04134_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10528__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08359_ net1849 net1006 net982 _04070_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11370_ _06818_ _06868_ net366 vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09795__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10321_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\] net832 net869 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\]
+ _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12235__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10544__A _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14016__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11339__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12000__A0 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13040_ _07535_ _02823_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09547__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10252_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\] net776 net708 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10183_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\] net918 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1203 net1206 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__buf_4
Xfanout1214 net1215 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__buf_4
X_16759__1303 vssd1 vssd1 vccd1 vccd1 _16759__1303/HI net1303 sky130_fd_sc_hd__conb_1
Xfanout1225 net1237 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1236 net1237 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__buf_4
XANTENNA_input39_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ net1222 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
Xfanout1247 net1249 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__buf_4
Xfanout260 net263 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
Xfanout1258 net1260 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_2
XANTENNA__08668__B team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout271 _06626_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11106__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_2
X_16730_ net1454 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
X_13942_ net1236 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
Xfanout293 _06791_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_1
XFILLER_0_92_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09180__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ clknet_leaf_101_wb_clk_i _02780_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13873_ net1229 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15612_ clknet_leaf_47_wb_clk_i _01752_ _00420_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12824_ team_02_WB.instance_to_wrap.top.a1.state\[1\] _07343_ _07345_ _07341_ vssd1
+ vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__o22a_1
X_16592_ clknet_leaf_98_wb_clk_i _02711_ _01385_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08684__A team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_104_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15543_ clknet_leaf_116_wb_clk_i _01683_ _00351_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12755_ _05736_ _05783_ _05829_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_57_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11314__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11706_ net245 net2511 net603 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XANTENNA__10093__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ clknet_leaf_11_wb_clk_i _01614_ _00282_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ net284 net2614 net432 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ net1136 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
X_11637_ net1001 net994 _07123_ team_02_WB.instance_to_wrap.top.pc\[1\] vssd1 vssd1
+ vccd1 vccd1 _07124_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09786__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__B2 _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14356_ net1091 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11568_ _05738_ _06001_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ team_02_WB.instance_to_wrap.top.pc\[6\] net1052 _07026_ net935 vssd1 vssd1
+ vccd1 vccd1 _03003_ sky130_fd_sc_hd__a22o_2
XFILLER_0_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold708 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10519_ net669 _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__nor2_1
Xhold719 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12145__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14287_ net1111 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10454__A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11499_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _06833_ _06837_ _06992_ vssd1
+ vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__a211o_1
XFILLER_0_106_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16026_ clknet_leaf_120_wb_clk_i _02166_ _00834_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13238_ team_02_WB.instance_to_wrap.top.ru.next_write_i _00006_ vssd1 vssd1 vccd1
+ vccd1 _02959_ sky130_fd_sc_hd__nor2_4
XANTENNA__09538__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16738__1283 vssd1 vssd1 vccd1 vccd1 _16738__1283/HI net1283 sky130_fd_sc_hd__conb_1
XFILLER_0_42_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11984__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16418__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13169_ net1026 _02931_ net1023 team_02_WB.instance_to_wrap.top.pc\[7\] vssd1 vssd1
+ vccd1 vccd1 _01488_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08210__A2 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10901__B _06415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _03443_ _03447_ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wire613_A _05230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09171__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10856__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09710__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ _03344_ _03370_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__xnor2_4
X_16859_ net1403 vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_2
XFILLER_0_36_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09400_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\] net775 net715 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\]
+ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_81_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07592_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] _03316_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\]
+ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 _03317_
+ sky130_fd_sc_hd__or4b_4
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09331_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\] net834 net830 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\]
+ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__a221o_1
XANTENNA__15592__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13270__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__A team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09262_ _04777_ _04778_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08213_ _03929_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09193_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\] net714 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08144_ _03829_ _03835_ net226 vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08075_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _03787_ vssd1 vssd1 vccd1
+ vccd1 _03796_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12055__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1135_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09529__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11894__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout595_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[10\] vssd1 vssd1 vccd1 vccd1
+ net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _02592_ vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _04491_ _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout762_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 team_02_WB.instance_to_wrap.top.a1.data\[3\] vssd1 vssd1 vccd1 vccd1 net1493
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 _02623_ vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08488__B _04185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 net124 vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _03649_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold68 _02572_ vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 team_02_WB.START_ADDR_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09162__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10847__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ _03540_ _03544_ _03545_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__nand3_1
XANTENNA__10847__B2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10870_ _06058_ _06063_ net365 vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09529_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\] net730 net698 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__a22o_1
XANTENNA__11642__B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13261__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10539__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ net645 _07205_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__nand2_1
X_16883__1427 vssd1 vssd1 vccd1 vccd1 _16883__1427/HI net1427 sky130_fd_sc_hd__conb_1
XANTENNA__10075__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ net363 net2377 net452 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08951__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ net1210 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
X_11422_ net517 net384 _06061_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__a21o_1
XANTENNA__09768__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15190_ net1256 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08670__C team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14141_ net1084 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11353_ _06358_ _06638_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\] net756 net732 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__a22o_1
X_14072_ net1195 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11284_ _06786_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__inv_2
X_13023_ _06273_ net233 _07443_ net978 _07542_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__o221a_1
X_10235_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\] net835 net815 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1000 _04264_ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_4
Xfanout1011 _03014_ vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_89_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1022 _00012_ vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__buf_2
X_10166_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\] net832 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\]
+ _05682_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__a221o_1
Xfanout1033 _04428_ vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09940__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1044 _04245_ vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1055 team_02_WB.instance_to_wrap.busy_o vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__buf_2
Xfanout1066 _00018_ vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__buf_2
XFILLER_0_83_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1077 net1079 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_4
X_10097_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\] net737 net721 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__a22o_1
X_14974_ net1257 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
Xfanout1088 net1199 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_2
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1099 net1103 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_4
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16713_ net1272 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
X_13925_ net1204 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
XANTENNA__08900__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13856_ net1228 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
X_16644_ clknet_leaf_100_wb_clk_i _02763_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08618__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12807_ _07234_ _07231_ _06124_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13787_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\]
+ _03275_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16575_ clknet_leaf_99_wb_clk_i _00001_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10449__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13252__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10999_ _06447_ _06510_ net369 vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15526_ clknet_leaf_43_wb_clk_i _01666_ _00334_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12738_ net379 _06579_ _06518_ _06484_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11979__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15457_ clknet_leaf_121_wb_clk_i _01597_ _00265_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12669_ net360 net2097 net436 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14408_ net1178 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
XANTENNA__09759__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15388_ clknet_leaf_48_wb_clk_i _01528_ _00196_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08967__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16240__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14339_ net1146 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
Xhold505 team_02_WB.instance_to_wrap.ramaddr\[3\] vssd1 vssd1 vccd1 vccd1 net1963
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold516 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap224 _03949_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_1
Xhold527 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold538 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08719__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08900_ net24 net1031 net989 net1807 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a22o_1
X_16009_ clknet_leaf_104_wb_clk_i _02149_ _00817_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09880_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\] net706 _05396_ vssd1
+ vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__a21o_1
XANTENNA__12603__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08831_ net106 net1043 net992 net1486 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09931__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1205 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _04296_ net847 _04363_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__and3_1
Xhold1227 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
X_07713_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] _03432_ _03433_ _03434_ vssd1
+ vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10829__A1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08693_ _04294_ _04319_ _04321_ _04310_ _04317_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__o311a_1
XFILLER_0_79_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13491__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12839__A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07644_ _03365_ _03366_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07575_ net2337 net189 _00017_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout343_A _07051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1085_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09314_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\] net747 net844 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10057__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__B2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09998__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11889__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15338__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09245_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\] net879 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16758__1302 vssd1 vssd1 vccd1 vccd1 _16758__1302/HI net1302 sky130_fd_sc_hd__conb_1
XFILLER_0_134_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1252_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A _06281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09176_ net542 _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08127_ _03803_ _03841_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08058_ _03757_ _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout977_A _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12513__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10020_ _05536_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__inv_2
Xinput103 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09922__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09135__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11971_ net361 net1831 net587 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13710_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] _03227_ net1240 vssd1
+ vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10922_ net407 _06435_ _06434_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10296__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14690_ net1202 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13641_ _03167_ _03181_ _03188_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__or3_1
X_10853_ net999 _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11245__A1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10048__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16360_ clknet_leaf_15_wb_clk_i _02500_ _01168_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09989__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ _03104_ _03115_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10784_ _05489_ net384 vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11799__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15311_ clknet_leaf_103_wb_clk_i _01454_ _00124_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12523_ net302 net2250 net447 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__mux2_1
XANTENNA__16263__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16291_ clknet_leaf_126_wb_clk_i _02431_ _01099_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15242_ clknet_leaf_65_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[1\]
+ _00055_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12454_ net274 net2027 net450 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__mux2_1
XANTENNA__08949__B1 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ net419 _06438_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15173_ net1241 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
X_12385_ net280 net2638 net459 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__mux2_1
X_14124_ net1082 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
X_11336_ net849 net952 net496 vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__o21a_2
XFILLER_0_61_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14055_ net1117 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
X_11267_ net373 _06535_ _06769_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12423__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13006_ team_02_WB.instance_to_wrap.top.pc\[21\] _06184_ _07525_ vssd1 vssd1 vccd1
+ vccd1 _07526_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09374__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10218_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\] net778 _05728_ _05733_
+ _05734_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__a2111oi_2
XANTENNA__09913__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10845__A2_N net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11198_ _05041_ _06600_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10451__B _04733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\] net741 net717 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\]
+ _05665_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09126__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14957_ net1147 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13473__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ net1218 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
XANTENNA__10287__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14888_ net1177 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16627_ clknet_leaf_98_wb_clk_i _02746_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13839_ net1232 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13225__A2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12433__A0 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16558_ clknet_leaf_93_wb_clk_i _02682_ _01365_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[109\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_57_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15509_ clknet_leaf_41_wb_clk_i _01649_ _00317_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_16489_ clknet_leaf_74_wb_clk_i net1601 _01297_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09030_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\] net929 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold302 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold313 team_02_WB.instance_to_wrap.ramload\[6\] vssd1 vssd1 vccd1 vccd1 net1771
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold324 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold335 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold346 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12841__B _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold357 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold368 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\] net884 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\]
+ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__a221o_1
Xhold379 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12333__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout804 _04535_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout815 _04521_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09365__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout826 net828 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_4
XANTENNA__09904__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ _05378_ _05379_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__nand2b_1
Xfanout837 net838 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__clkbuf_4
X_16882__1426 vssd1 vssd1 vccd1 vccd1 _16882__1426/HI net1426 sky130_fd_sc_hd__conb_1
Xfanout848 _04358_ vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_2
XANTENNA_fanout293_A _06791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10361__B _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net861 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08814_ net114 net1043 net993 net1772 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__a22o_1
Xhold1002 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13953__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1013 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09794_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\] net734 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a22o_1
Xhold1035 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16136__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09117__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1046 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ net848 _04365_ _04370_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__and3_4
Xhold1057 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11475__A1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10278__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _04262_ _04293_ _04294_ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__and4_4
XANTENNA__11475__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07627_ _03324_ _03327_ team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1
+ vccd1 vccd1 _03350_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout725_A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07558_ team_02_WB.instance_to_wrap.top.edg2.flip2 vssd1 vssd1 vccd1 vccd1 _03299_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_64_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12508__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10817__A _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09228_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\] net779 _04743_ _04744_
+ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13220__A1_N _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09159_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\] net893 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\]
+ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12170_ net337 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\] net465 vssd1
+ vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__mux2_1
XANTENNA__10202__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11121_ _06320_ _06339_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ _06557_ _06562_ _06561_ _06558_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_1662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10003_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\] net776 _05517_ _05519_
+ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__a211o_1
X_15860_ clknet_leaf_10_wb_clk_i _02000_ _00668_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09108__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ net1184 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
X_15791_ clknet_leaf_34_wb_clk_i _01931_ _00599_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15503__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16629__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11954_ net272 net2406 net585 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__mux2_1
X_14742_ net1096 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10905_ _06134_ net655 net495 team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] net497
+ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__a221o_1
X_14673_ net1107 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11885_ net289 net2649 net487 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16412_ clknet_leaf_66_wb_clk_i _02547_ _01220_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13624_ team_02_WB.instance_to_wrap.top.a1.row2\[27\] _03118_ _03169_ _03170_ _03175_
+ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__a2111o_1
X_10836_ _06349_ _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13555_ net1049 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] _03109_ vssd1
+ vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__and3_1
X_16343_ clknet_leaf_14_wb_clk_i _02483_ _01151_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12418__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ _04611_ _05959_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12506_ net344 net2224 net557 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__mux2_1
X_16274_ clknet_leaf_8_wb_clk_i _02414_ _01082_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13486_ team_02_WB.START_ADDR_VAL_REG\[26\] net1070 _04259_ vssd1 vssd1 vccd1 vccd1
+ net210 sky130_fd_sc_hd__a21o_1
X_10698_ team_02_WB.instance_to_wrap.top.pc\[16\] _06192_ _06214_ vssd1 vssd1 vccd1
+ vccd1 _06215_ sky130_fd_sc_hd__a21o_1
XANTENNA__10446__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15225_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[16\]
+ _00038_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12437_ net354 net2010 net455 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16829__1373 vssd1 vssd1 vccd1 vccd1 _16829__1373/HI net1373 sky130_fd_sc_hd__conb_1
XFILLER_0_65_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09595__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15156_ net1247 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
X_12368_ net339 net2275 net564 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08631__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14107_ net1156 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11319_ _06715_ _06819_ net397 vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__mux2_1
X_15087_ net1104 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
XANTENNA__10462__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12153__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ net326 net2079 net571 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__mux2_1
X_14038_ net1095 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11992__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16757__1301 vssd1 vssd1 vccd1 vccd1 _16757__1301/HI net1301 sky130_fd_sc_hd__conb_1
XFILLER_0_78_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15989_ clknet_leaf_43_wb_clk_i _02129_ _00797_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11293__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ _04216_ net1630 net850 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11457__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08461_ net1752 net1005 net981 _04163_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10680__A2 _05740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08392_ _04090_ _04092_ _04099_ _04088_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__o31a_1
XFILLER_0_64_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12836__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12328__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ net1056 _04528_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__nor2_8
XANTENNA__13948__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12852__A _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout306_A _06891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 _02588_ vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 team_02_WB.instance_to_wrap.ramaddr\[29\] vssd1 vssd1 vccd1 vccd1 net1579
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold132 team_02_WB.instance_to_wrap.top.a1.row1\[120\] vssd1 vssd1 vccd1 vccd1 net1590
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _02624_ vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _02598_ vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _02607_ vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12063__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold176 _02595_ vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1215_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 team_02_WB.instance_to_wrap.ramstore\[19\] vssd1 vssd1 vccd1 vccd1 net1645
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _07189_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_6
Xhold198 net123 vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09915_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\] net712 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15526__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 _04453_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout675_A _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout656 net657 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09846_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\] net809 net898 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\]
+ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__a221o_1
Xfanout667 net668 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_2
Xfanout678 net681 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_8
Xfanout689 _04399_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_4
X_09777_ _05292_ _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_124_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08728_ team_02_WB.instance_to_wrap.top.i_ready net1001 net790 net552 vssd1 vssd1
+ vccd1 vccd1 _04357_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15676__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08659_ net1058 net1057 vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10671__A2 _05580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11670_ _05987_ _07155_ _07150_ _05986_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10621_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] net995 vssd1 vssd1 vccd1
+ vccd1 _06138_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_137_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12238__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10547__A _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13340_ net1807 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[2\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_107_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ _06060_ _06068_ net393 vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13271_ team_02_WB.instance_to_wrap.top.pc\[24\] team_02_WB.instance_to_wrap.top.ru.state\[5\]
+ _06588_ net935 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10483_ net407 net498 _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_129_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15010_ net1229 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09577__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12222_ net1710 net288 net618 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__mux2_1
XANTENNA__16301__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input69_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13577__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12153_ net269 net2521 net462 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09329__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11104_ net379 _06606_ _06357_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__o21ba_1
XANTENNA__13125__B2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ net2557 net262 net583 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
XANTENNA__11136__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16451__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ net408 _06350_ _06400_ _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__a31o_1
X_15912_ clknet_leaf_16_wb_clk_i _02052_ _00720_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12701__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16892_ net1436 vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__buf_2
XFILLER_0_95_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15843_ clknet_leaf_127_wb_clk_i _01983_ _00651_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15774_ clknet_leaf_118_wb_clk_i _01914_ _00582_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12986_ team_02_WB.instance_to_wrap.top.pc\[9\] _05536_ vssd1 vssd1 vccd1 vccd1 _07506_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09501__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14725_ net1128 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
X_11937_ net362 net2210 net484 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__mux2_1
XANTENNA__08855__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11868_ net354 net2074 net492 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14656_ net1155 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
XANTENNA__08626__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10819_ _06331_ _06334_ net366 vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__mux2_1
X_13607_ _03289_ net1049 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] _03115_
+ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__and4_1
XANTENNA__12148__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11799_ net356 net2610 net593 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16881__1425 vssd1 vssd1 vccd1 vccd1 _16881__1425/HI net1425 sky130_fd_sc_hd__conb_1
X_14587_ net1157 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16326_ clknet_leaf_44_wb_clk_i _02466_ _01134_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13538_ _03093_ _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09280__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11987__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16257_ clknet_leaf_121_wb_clk_i _02397_ _01065_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13469_ team_02_WB.START_ADDR_VAL_REG\[9\] net1068 net1002 vssd1 vssd1 vccd1 vccd1
+ net223 sky130_fd_sc_hd__a21o_1
XFILLER_0_125_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09568__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15208_ clknet_leaf_59_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_dready _00021_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.d_ready sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput204 net204 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16188_ clknet_leaf_49_wb_clk_i _02328_ _00996_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09032__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10178__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput215 net215 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XANTENNA__15549__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11288__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15139_ net1245 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07961_ _03681_ _03683_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_71_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09700_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\] net763 net689 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\]
+ _05214_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11678__A1 _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ _03584_ _03603_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12611__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12875__B1 _07394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09740__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\] net809 net912 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09562_ _05071_ _05074_ _05076_ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__nor4_1
XFILLER_0_78_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09099__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08513_ _04171_ _04202_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09493_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\] net756 net730 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__a22o_1
XANTENNA__08846__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12847__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_A _06530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08444_ _04145_ _04146_ _04147_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08375_ _04084_ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__and2_1
XANTENNA__12058__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1165_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09271__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11897__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07676__A team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09559__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10814__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13107__B2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout420 _05716_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__clkbuf_2
Xfanout431 _07229_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11669__A1 _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout442 net445 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout453 _07222_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_4
XANTENNA__12521__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_35_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout475 _07206_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout486 _07198_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_50_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09731__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout497 _06250_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09829_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\] net706 _05344_ _05345_
+ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__a211o_1
XANTENNA__12919__A1_N net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12840_ _04842_ _06171_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16828__1372 vssd1 vssd1 vccd1 vccd1 _16828__1372/HI net1372 sky130_fd_sc_hd__conb_1
XFILLER_0_9_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12094__A1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12771_ _06942_ _07039_ _07059_ _07082_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08837__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11661__A _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11722_ net298 net2030 net603 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
X_14510_ net1114 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15490_ clknet_leaf_123_wb_clk_i _01630_ _00298_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14441_ net1102 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
X_11653_ _05336_ _05932_ _05989_ _05380_ _05559_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__o2111ai_1
XTAP_TAPCELL_ROW_29_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09798__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ _06104_ _06108_ _06120_ _06103_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a211o_1
X_14372_ net1129 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
X_11584_ net401 _06998_ _07070_ _07072_ net381 vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__o221a_1
XFILLER_0_80_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16756__1300 vssd1 vssd1 vccd1 vccd1 _16756__1300/HI net1300 sky130_fd_sc_hd__conb_1
XFILLER_0_68_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16111_ clknet_leaf_38_wb_clk_i _02251_ _00919_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13323_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] _03011_ _03010_ net1675
+ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10535_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap609 _05781_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_111_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13254_ _06415_ _02964_ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__or2_1
X_16042_ clknet_leaf_128_wb_clk_i _02182_ _00850_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ _04906_ _04908_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__or2_4
XFILLER_0_49_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12205_ net356 net2720 net577 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13185_ team_02_WB.instance_to_wrap.top.pc\[4\] net1023 _02944_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01485_ sky130_fd_sc_hd__a22o_1
X_10397_ _05690_ net505 vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12136_ net338 net2147 net468 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12431__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ net333 net1820 net472 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_97_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09722__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ net947 _06523_ _06529_ net607 vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__o211a_4
XANTENNA__09306__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16875_ net1419 vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_26_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15826_ clknet_leaf_12_wb_clk_i _01966_ _00634_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13282__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15757_ clknet_leaf_32_wb_clk_i _01897_ _00565_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08828__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ team_02_WB.instance_to_wrap.top.pc\[5\] _05695_ vssd1 vssd1 vccd1 vccd1 _07489_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_1362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10096__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14708_ net1076 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16347__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15688_ clknet_leaf_16_wb_clk_i _01828_ _00496_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14639_ net1165 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14882__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08160_ _03840_ net226 vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__and2_1
XANTENNA__09253__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11596__B1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16309_ clknet_leaf_43_wb_clk_i _02449_ _01117_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15371__CLK clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08091_ _03784_ _03810_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__xnor2_4
XANTENNA__08461__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09961__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07944_ _03602_ _03605_ _03638_ _03627_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__a31o_1
XANTENNA__12341__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07875_ _03596_ _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09614_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\] net761 net757 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\] net821 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13273__B1 _06618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ _04970_ _04991_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10809__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08427_ _04130_ _04133_ _04128_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15714__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08358_ _04056_ _04064_ _04067_ _04069_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a31o_2
XFILLER_0_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09244__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08289_ _03966_ _03979_ _03989_ _03970_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__o31ai_1
XANTENNA__12516__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10320_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\] net921 net877 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15864__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10544__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10251_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\] net760 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\]
+ _05765_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_128_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10397__A_N _05690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10182_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\] net914 net817 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\]
+ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1204 net1206 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1215 net1225 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_4
Xfanout1226 net1230 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_4
XANTENNA__12251__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1237 net1265 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_4
X_14990_ net1223 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout250 _06498_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1248 net1249 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__buf_4
Xfanout261 net263 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09704__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1259 net1260 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__buf_4
X_16880__1424 vssd1 vssd1 vccd1 vccd1 _16880__1424/HI net1424 sky130_fd_sc_hd__conb_1
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_2
Xfanout283 _06657_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
X_13941_ net1257 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
Xfanout294 _06791_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14967__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16660_ clknet_leaf_100_wb_clk_i _02779_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13872_ net1227 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15611_ clknet_leaf_127_wb_clk_i _01751_ _00419_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12823_ _04306_ _07340_ _07344_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__a21o_1
XANTENNA__13264__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16591_ clknet_leaf_99_wb_clk_i _02710_ _01384_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08684__B team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15542_ clknet_leaf_47_wb_clk_i _01682_ _00350_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12754_ _05557_ _05604_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09483__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11705_ net241 net1886 net604 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15394__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15473_ clknet_leaf_50_wb_clk_i _01613_ _00281_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ net272 net2462 net430 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14424_ net1220 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
X_11636_ net849 _06162_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__nand2_1
XANTENNA__09235__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11578__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire640 _04564_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_1
XANTENNA__12426__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14355_ net1168 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
X_11567_ _05738_ _05911_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10250__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13319__B2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13306_ net1518 net983 net964 _03002_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__a22o_1
X_10518_ _04569_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold709 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
X_14286_ net1114 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
X_11498_ team_02_WB.instance_to_wrap.top.pc\[8\] net973 _06991_ net1001 vssd1 vssd1
+ vccd1 vccd1 _06992_ sky130_fd_sc_hd__a22o_1
Xmax_cap428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_2
X_13237_ _02958_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16025_ clknet_leaf_18_wb_clk_i _02165_ _00833_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10449_ _04630_ _04652_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10002__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__B1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13168_ _07009_ net232 _02928_ net977 _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__o221a_1
X_12119_ net268 net2200 net466 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
XANTENNA__12161__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ _07519_ _02872_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07660_ _03380_ _03382_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16858_ net1402 vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_2
XANTENNA__10856__A2 _06365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15809_ clknet_leaf_121_wb_clk_i _01949_ _00617_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_07591_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__nand2_1
X_16789_ net1333 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XANTENNA__15737__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08594__B net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09330_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\] net883 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a22o_1
XANTENNA__10069__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09474__A2 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09261_ _04714_ _04733_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08212_ _03897_ _03922_ _03928_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_56_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11018__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09192_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\] net742 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\]
+ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__a221o_1
XANTENNA__15887__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09226__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ _03852_ _03861_ _03856_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_12_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12230__A1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12336__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10241__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ _03764_ _03787_ _03791_ _03794_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_86_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16827__1371 vssd1 vssd1 vccd1 vccd1 _16827__1371/HI net1371 sky130_fd_sc_hd__conb_1
XANTENNA__13956__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12860__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1128_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09934__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout490_A _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 team_02_WB.instance_to_wrap.ramstore\[9\] vssd1 vssd1 vccd1 vccd1 net1472
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _04326_ _04492_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_32_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold25 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[16\] vssd1 vssd1
+ vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 net183 vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 net176 vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03636_ _03611_ vssd1 vssd1
+ vccd1 vccd1 _03650_ sky130_fd_sc_hd__o21bai_1
Xhold58 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ net1516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 team_02_WB.instance_to_wrap.top.a1.data\[10\] vssd1 vssd1 vccd1 vccd1 net1527
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout755_A _04375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14787__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07858_ _03578_ _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07789_ _03507_ _03509_ _03499_ _03501_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout922_A _04513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09528_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\] net762 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09465__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10539__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09459_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\] net814 net911 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12470_ net355 net2416 net452 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11421_ net424 _06473_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__nand2_1
XANTENNA__12246__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10555__A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140_ net1147 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
XANTENNA__10232__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08670__D team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11352_ _06104_ _06851_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08025__A team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10303_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\] net708 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a22o_1
X_14071_ net1173 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11283_ _06263_ _06785_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _07540_ _07541_ net230 vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_1372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input51_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\] net811 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\]
+ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1001 _04263_ vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1012 net1013 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10165_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\] net828 net816 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10290__A _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1023 net1025 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__buf_2
Xfanout1034 _04428_ vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1045 _04173_ vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
Xfanout1056 team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1 vccd1
+ vccd1 net1056 sky130_fd_sc_hd__buf_4
X_10096_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\] net765 net741 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__a22o_1
XANTENNA__13485__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1067 _00018_ vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_4
X_14973_ net1248 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_4
XANTENNA_output138_A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1089 net1097 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_4
XFILLER_0_136_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16712_ net1271 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XANTENNA__10299__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ net1216 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12929__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16643_ clknet_leaf_100_wb_clk_i net1696 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_13855_ net1222 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12806_ _07323_ _07324_ _07322_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16574_ clknet_leaf_99_wb_clk_i _00000_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_13786_ _03276_ _03277_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__nor2_1
X_10998_ _06314_ _06325_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__or2_1
XANTENNA__09456__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15525_ clknet_leaf_32_wb_clk_i _01665_ _00333_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12737_ _07260_ _06924_ _07259_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__and3b_1
XFILLER_0_123_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15456_ clknet_leaf_108_wb_clk_i _01596_ _00264_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12668_ net355 net2159 net436 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14407_ net1102 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12156__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ net945 _07104_ _07106_ net605 vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__o211a_1
X_15387_ clknet_leaf_126_wb_clk_i _01527_ _00195_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10465__A _04885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ net338 net2538 net441 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14338_ net1205 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
Xhold506 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap225 _03936_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold517 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11995__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold528 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ net1082 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16008_ clknet_leaf_16_wb_clk_i _02148_ _00816_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_41_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08830_ net117 net1042 net992 net1633 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a22o_1
Xhold1206 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1217 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] vssd1 vssd1 vccd1 vccd1
+ net2675 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\] net774 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a22o_1
Xhold1228 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1239 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13476__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ _03433_ _03434_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__and2_1
X_08692_ net1057 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] net1059 vssd1
+ vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07643_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] _03334_ _03360_ vssd1 vssd1
+ vccd1 vccd1 _03366_ sky130_fd_sc_hd__or3_1
XANTENNA__13228__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07574_ team_02_WB.instance_to_wrap.top.pad.count\[0\] team_02_WB.instance_to_wrap.top.pad.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__and2b_1
XFILLER_0_76_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09447__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\] net739 net715 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12855__A _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09244_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\] net826 net891 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\]
+ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1078_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16065__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09175_ net972 _04691_ net545 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__o21ai_4
XANTENNA__12066__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1245_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ _03842_ _03843_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10214__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09080__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08057_ _03734_ _03756_ _03736_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09907__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__A1 _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput104 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08959_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\] net781 net753 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__a22o_1
XANTENNA__09135__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11970_ net354 net1943 net587 vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09686__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10921_ _06302_ _06306_ net365 vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08894__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13219__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10852_ _06272_ _06367_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__nand2_1
X_13640_ team_02_WB.instance_to_wrap.top.a1.row2\[15\] _03103_ _03165_ _03117_ team_02_WB.instance_to_wrap.top.a1.row1\[63\]
+ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__a32o_1
XANTENNA__09438__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10783_ _06297_ _06298_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__or2_1
X_13571_ net1047 _03103_ _03113_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ clknet_leaf_65_wb_clk_i _01453_ _00123_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12522_ net294 net2431 net449 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__mux2_1
X_16290_ clknet_leaf_124_wb_clk_i _02430_ _01098_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input99_A wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[0\]
+ _00054_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12453_ net288 net1950 net452 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__mux2_1
XANTENNA__14980__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10205__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11404_ net423 _06451_ _06900_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__o21ai_2
X_15172_ net1243 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
X_12384_ net270 net1924 net458 vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11335_ _06194_ net654 _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] _06835_
+ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__a221o_1
X_14123_ net1202 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12704__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07594__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11266_ net378 _06539_ _06639_ _06534_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__o22a_1
X_14054_ net1089 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10217_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\] net766 net718 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__a22o_1
X_13005_ _07460_ _07524_ vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11197_ _06117_ _06696_ _06699_ _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_118_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10148_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\] net773 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14956_ net1079 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
X_10079_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\] net823 net819 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\]
+ _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__a221o_1
XANTENNA__08629__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ net1204 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14887_ net1112 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16626_ clknet_leaf_100_wb_clk_i _02745_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13838_ net1232 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
X_16826__1370 vssd1 vssd1 vccd1 vccd1 _16826__1370/HI net1370 sky130_fd_sc_hd__conb_1
XFILLER_0_130_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16088__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16557_ clknet_leaf_94_wb_clk_i _02681_ _01364_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_13769_ _03265_ _03266_ net961 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15051__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15508_ clknet_leaf_12_wb_clk_i _01648_ _00316_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16488_ clknet_leaf_71_wb_clk_i net1504 _01296_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15439_ clknet_leaf_38_wb_clk_i _01579_ _00247_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14890__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09601__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold303 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold314 team_02_WB.instance_to_wrap.ramaddr\[17\] vssd1 vssd1 vccd1 vccd1 net1772
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15925__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12614__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold369 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\] net912 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout805 net808 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout816 _04521_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_2
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_8
X_09862_ _05355_ _05376_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout838 _04470_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_4
Xfanout849 _04325_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_2
Xhold1003 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ net115 net1044 net991 net1500 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__a22o_1
X_09793_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\] net762 net722 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\]
+ _05309_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__a221o_1
Xhold1014 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1025 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1047 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _04302_ net931 _04359_ _04368_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1058 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09668__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08675_ _04298_ _04299_ _04300_ _04303_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__and4_1
XFILLER_0_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1195_A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07626_ team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] _03324_ _03327_ vssd1 vssd1
+ vccd1 vccd1 _03349_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07557_ net1057 vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout718_A _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09840__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09227_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\] net691 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09158_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\] net921 net877 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13202__A2_N _02955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09053__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08109_ _03824_ _03825_ _03820_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08800__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\] net914 net809 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\]
+ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a221o_1
XANTENNA__12524__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10833__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14305__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11120_ net398 _06511_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold870 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold881 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _06151_ _06152_ _06233_ net974 vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__o31a_1
Xhold892 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10002_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\] net716 net708 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\]
+ _05518_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15136__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14810_ net1184 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
X_15790_ clknet_leaf_27_wb_clk_i _01930_ _00598_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09659__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ net1187 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11953_ net290 net2078 net587 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16230__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10904_ net975 _06417_ _06418_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__and3_1
X_14672_ net1110 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08973__A team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11884_ net277 net2594 net488 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__mux2_1
X_16411_ clknet_leaf_67_wb_clk_i _02546_ _01219_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13623_ _03132_ _03172_ _03173_ _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ net546 net397 vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_101_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16342_ clknet_leaf_52_wb_clk_i _02482_ _01150_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13554_ _03107_ _03108_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__nor2_2
XANTENNA__09292__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766_ net2213 net243 net643 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__mux2_1
XANTENNA__16380__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09831__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12505_ net350 net1909 net559 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__mux2_1
X_16273_ clknet_leaf_50_wb_clk_i _02413_ _01081_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10697_ _06195_ _06212_ _06213_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__a21oi_1
X_13485_ team_02_WB.START_ADDR_VAL_REG\[25\] net1068 net1002 vssd1 vssd1 vccd1 vccd1
+ net209 sky130_fd_sc_hd__a21o_1
XFILLER_0_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15224_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[15\]
+ _00037_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_12436_ net356 net2356 net454 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12942__B _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15155_ net1244 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12434__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ net330 net1959 net563 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__mux2_1
XANTENNA__14215__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14106_ net1184 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _06771_ _06818_ net371 vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__mux2_1
X_15086_ net1236 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
X_12298_ net323 net2496 net571 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14037_ net1215 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
X_11249_ _06502_ _06639_ _06752_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09898__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15988_ clknet_leaf_10_wb_clk_i _02128_ _00796_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire519_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14939_ net1157 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08460_ _04157_ _04162_ _04158_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16609_ clknet_leaf_80_wb_clk_i _02728_ _01402_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08391_ net1617 net1005 net981 _04100_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a22o_1
XANTENNA__12609__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09283__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09822__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10129__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09012_ net1056 _04295_ _04297_ net951 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__and4_4
XFILLER_0_66_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09035__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12852__B _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold100 _02564_ vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold111 team_02_WB.instance_to_wrap.ramstore\[16\] vssd1 vssd1 vccd1 vccd1 net1569
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12344__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold122 team_02_WB.instance_to_wrap.ramload\[15\] vssd1 vssd1 vccd1 vccd1 net1580
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__A0 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold133 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16103__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold144 team_02_WB.instance_to_wrap.ramstore\[7\] vssd1 vssd1 vccd1 vccd1 net1602
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 team_02_WB.instance_to_wrap.top.a1.row1\[11\] vssd1 vssd1 vccd1 vccd1 net1613
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 team_02_WB.START_ADDR_VAL_REG\[28\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold177 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _02581_ vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _02619_ vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13964__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09914_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\] net752 net708 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__a22o_1
X_16736__1282 vssd1 vssd1 vccd1 vccd1 _16736__1282/HI net1282 sky130_fd_sc_hd__conb_1
Xfanout602 _07189_ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_4
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1110_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1208_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 _04453_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_1
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\] net914 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__a22o_1
Xfanout657 _06123_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout570_A _07217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 _06038_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_4
Xfanout679 net681 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_4
XANTENNA__16253__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09776_ net610 _05290_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_124_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _04328_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__inv_2
XANTENNA__10120__A2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07609_ team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] _03331_ vssd1 vssd1 vccd1
+ vccd1 _03332_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08589_ net43 net42 net45 net44 vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__or4_2
XANTENNA__12519__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ team_02_WB.instance_to_wrap.top.pc\[29\] _06134_ vssd1 vssd1 vccd1 vccd1
+ _06137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09274__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10547__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09813__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10551_ net366 _06063_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10039__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13270_ net1707 net985 net966 _02984_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a22o_1
X_10482_ _05833_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__or2_1
XANTENNA__11908__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12221_ net1795 net279 net617 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12254__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10563__A _04631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10187__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ net260 net2725 net463 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11103_ _06610_ _06611_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12083_ net1893 net266 net583 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15911_ clknet_leaf_29_wb_clk_i _02051_ _00719_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11034_ net408 _06544_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16891_ net1435 vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__buf_2
XANTENNA__11687__A2 _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12884__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__A2 _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15842_ clknet_leaf_122_wb_clk_i _01982_ _00650_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07591__B team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09176__A_N net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15620__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ clknet_leaf_51_wb_clk_i _01913_ _00581_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11439__A2 _06931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ _07484_ _07504_ _07482_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_103_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08304__A2 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ net1127 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11936_ net352 net2634 net484 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10111__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14655_ net1183 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11867_ net359 net2640 net490 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__mux2_1
XANTENNA__12429__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ team_02_WB.instance_to_wrap.top.a1.row1\[19\] _03111_ _03116_ team_02_WB.instance_to_wrap.top.a1.row1\[123\]
+ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10818_ _06332_ _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nand2_1
X_14586_ net1167 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ net341 net1829 net596 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
XANTENNA__09804__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16325_ clknet_leaf_33_wb_clk_i _02465_ _01133_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13537_ _03072_ _03078_ _03082_ _03075_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_82_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10749_ team_02_WB.instance_to_wrap.top.pc\[22\] team_02_WB.instance_to_wrap.top.pc\[21\]
+ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16256_ clknet_leaf_106_wb_clk_i _02396_ _01064_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13468_ team_02_WB.START_ADDR_VAL_REG\[8\] _04260_ vssd1 vssd1 vccd1 vccd1 net222
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13281__A1_N _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15207_ clknet_leaf_59_wb_clk_i net1016 _00020_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.i_ready
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12419_ net277 net2177 net456 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16187_ clknet_leaf_126_wb_clk_i _02327_ _00995_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12164__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10473__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13399_ team_02_WB.instance_to_wrap.ramload\[28\] net1012 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[28\] sky130_fd_sc_hd__and2_1
Xoutput205 net205 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_23_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput216 net216 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15138_ net1243 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16276__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07960_ _03656_ _03673_ _03678_ _03682_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__o2bb2a_1
X_15069_ net1258 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
XANTENNA__12324__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07891_ _03612_ _03613_ _03608_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a21o_1
XANTENNA__08597__B _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\] net904 net889 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a22o_1
XANTENNA__10350__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09561_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\] net829 net894 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\]
+ _05077_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08512_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[6\] net980 vssd1 vssd1 vccd1
+ vccd1 _04203_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09492_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\] net768 _05000_ _05001_
+ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10102__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12847__B _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ _04146_ _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__nor2_1
XANTENNA__12339__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11243__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08374_ _04072_ _04075_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13959__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1158_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12074__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10169__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout785_A _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08782__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16805__1349 vssd1 vssd1 vccd1 vccd1 _16805__1349/HI net1349 sky130_fd_sc_hd__conb_1
XANTENNA__11118__A1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout432 _07229_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout443 net445 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout454 net457 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_126_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout465 _07213_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout476 _07206_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09828_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\] net782 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a22o_1
Xfanout487 _07198_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_4
XFILLER_0_119_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10341__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09759_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\] net822 net907 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15793__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12770_ _07112_ _07136_ _07261_ _07271_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__a41o_1
XANTENNA__09495__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13291__B2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11721_ net310 net2387 net603 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__mux2_1
XANTENNA__11661__B _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12249__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10558__A _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16149__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14440_ net1176 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
X_11652_ _04482_ _04488_ _04565_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__or3_2
XFILLER_0_7_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10603_ _04569_ _06110_ net662 _04568_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__a221o_1
X_14371_ net1133 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11583_ net388 _07071_ net392 vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12773__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16110_ clknet_leaf_8_wb_clk_i _02250_ _00918_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input81_A wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13322_ _04174_ _03010_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10534_ _06047_ _06050_ net365 vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16041_ clknet_leaf_120_wb_clk_i _02181_ _00849_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16299__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11389__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13253_ team_02_WB.instance_to_wrap.ramaddr\[30\] net986 net966 _02972_ vssd1 vssd1
+ vccd1 vccd1 _01449_ sky130_fd_sc_hd__a22o_1
X_10465_ _04885_ _04905_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ net343 net2695 net580 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__mux2_1
X_10396_ net506 _05690_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nand2b_1
X_13184_ net228 _02941_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12135_ net330 net1892 net467 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
XANTENNA__08698__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__A1 _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12066_ net326 net1862 net472 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11017_ net975 _06524_ _06527_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_105_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16874_ net1418 vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_105_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10332__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15825_ clknet_leaf_21_wb_clk_i _01965_ _00633_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15756_ clknet_leaf_15_wb_clk_i _01896_ _00564_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ _05695_ team_02_WB.instance_to_wrap.top.pc\[5\] vssd1 vssd1 vccd1 vccd1 _07488_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09486__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13282__B2 _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14707_ net1168 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
X_11919_ net291 net1894 net484 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12159__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15687_ clknet_leaf_26_wb_clk_i _01827_ _00495_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12899_ _07372_ _07418_ _07373_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_64_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14638_ net1114 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16735__1281 vssd1 vssd1 vccd1 vccd1 _16735__1281/HI net1281 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_60_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15516__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13585__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14569_ net1109 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11596__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ clknet_leaf_12_wb_clk_i _02448_ _01116_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_08090_ _03784_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_67_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16239_ clknet_leaf_36_wb_clk_i _02379_ _01047_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15666__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08764__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12622__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__and3b_2
XFILLER_0_76_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07943_ _03631_ _03665_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07874_ _03558_ _03566_ _03589_ _03561_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_121_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10323__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09613_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\] net762 net742 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\] net786 _05055_ _05059_
+ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13273__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12069__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09475_ net971 _04990_ net543 vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_138_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08426_ _04106_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_134_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08357_ _04050_ _04051_ _04057_ _04068_ _04044_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__a32oi_1
XFILLER_0_62_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout700_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16441__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08288_ _03962_ _03988_ _03979_ _03970_ _03966_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11339__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11002__A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\] net732 net728 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\]
+ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a221o_1
XANTENNA__09401__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10181_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\] net922 net906 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12532__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1205 net1206 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__buf_4
XFILLER_0_100_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1216 net1225 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__buf_4
Xfanout1227 net1230 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__buf_2
XFILLER_0_100_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1238 net1239 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__buf_4
Xfanout240 _06424_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
Xfanout251 net254 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_2
Xfanout1249 net1250 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_4
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout273 _06740_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_2
X_13940_ net1257 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11511__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout284 net287 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_2
Xfanout295 _06791_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_92_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09180__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ net1231 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15610_ clknet_leaf_118_wb_clk_i _01750_ _00418_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12822_ _04305_ _07340_ _07344_ team_02_WB.instance_to_wrap.top.a1.state\[2\] vssd1
+ vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16590_ clknet_leaf_98_wb_clk_i _02709_ _01383_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09468__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15541_ clknet_leaf_43_wb_clk_i _01681_ _00349_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12753_ _05513_ _05904_ _05929_ _07276_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__or4_1
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08140__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11704_ _04291_ net645 _07188_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__or3_4
X_15472_ clknet_leaf_40_wb_clk_i _01612_ _00280_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12684_ net289 net1753 net432 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ net1172 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ _07119_ _07121_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11578__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14354_ net1121 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
Xwire630 _05121_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_1
XFILLER_0_4_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11566_ net375 _06898_ _07055_ _06695_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__a211o_1
XANTENNA__09640__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13305_ team_02_WB.instance_to_wrap.top.pc\[7\] net1051 _07007_ net933 vssd1 vssd1
+ vccd1 vccd1 _03002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10517_ _04589_ _04608_ _04611_ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__a22oi_1
X_14285_ net1154 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11497_ _06257_ _06990_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_113_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16024_ clknet_leaf_19_wb_clk_i _02164_ _00832_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13236_ team_02_WB.instance_to_wrap.top.d_ready _03308_ _04268_ _04346_ vssd1 vssd1
+ vccd1 vccd1 _02958_ sky130_fd_sc_hd__or4_1
X_10448_ _04462_ _05963_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12442__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ net228 _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10379_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\] net809 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12118_ net260 net2668 net466 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13098_ _07464_ _07465_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11058__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11591__A1_N net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12049_ net256 net1896 net471 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10305__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16314__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09171__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16857_ net1401 vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_2
XFILLER_0_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15808_ clknet_leaf_106_wb_clk_i _01948_ _00616_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_07590_ team_02_WB.instance_to_wrap.top.a1.state\[2\] _03313_ vssd1 vssd1 vccd1 vccd1
+ _03315_ sky130_fd_sc_hd__nand2_1
X_16788_ net1332 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
XANTENNA__09459__B1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15739_ clknet_leaf_126_wb_clk_i _01879_ _00547_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ net538 _04775_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16804__1348 vssd1 vssd1 vccd1 vccd1 _16804__1348/HI net1348 sky130_fd_sc_hd__conb_1
XFILLER_0_111_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08211_ _03922_ _03923_ _03897_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09191_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\] net758 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12617__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11521__S net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08142_ _03854_ _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09631__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08073_ _03722_ _03763_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12352__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1023_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__B _06970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] _04330_ net651 team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout483_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[6\] vssd1 vssd1 vccd1 vccd1
+ net1473 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 team_02_WB.instance_to_wrap.top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 net1484
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold37 team_02_WB.instance_to_wrap.top.a1.data\[2\] vssd1 vssd1 vccd1 vccd1 net1495
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03611_ _03637_ vssd1 vssd1
+ vccd1 vccd1 _03649_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_97_1650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold48 team_02_WB.instance_to_wrap.top.a1.data\[11\] vssd1 vssd1 vccd1 vccd1 net1506
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_02_WB.START_ADDR_VAL_REG\[4\] vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__A2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07857_ _03545_ _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07788_ _03507_ _03509_ _03499_ _03501_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_49_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09527_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\] net718 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout915_A _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09458_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\] net834 net891 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\]
+ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09870__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08409_ _04115_ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__nand2_1
XANTENNA__12527__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ _04886_ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_95_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11420_ _05928_ net661 net658 _05420_ _06916_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__a221o_1
XANTENNA__08425__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09622__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11351_ net419 _06348_ _06850_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15981__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10302_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\] net764 net728 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__a22o_1
X_14070_ net1095 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
X_11282_ team_02_WB.instance_to_wrap.top.pc\[17\] _06262_ vssd1 vssd1 vccd1 vccd1
+ _06785_ sky130_fd_sc_hd__nor2_1
X_13021_ _07445_ _07538_ _07539_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__and3_1
XANTENNA__09925__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\] net916 net807 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__a22o_1
XANTENNA__12262__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15211__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16337__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\] net812 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\]
+ _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_89_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1002 _04259_ vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__buf_2
Xfanout1013 _03014_ vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08041__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1024 net1025 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__buf_2
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_2
Xfanout1046 _04171_ vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__buf_2
Xfanout1057 team_02_WB.instance_to_wrap.top.a1.instruction\[13\] vssd1 vssd1 vccd1
+ vccd1 net1057 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10095_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\] net842 _05609_ _05611_
+ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a211o_1
X_14972_ net1257 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
XANTENNA__09689__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1068 net1070 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_2
Xfanout1079 net1199 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_4
X_13923_ net1221 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
XANTENNA__09153__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16711_ net1270 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08900__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16642_ clknet_leaf_102_wb_clk_i _02761_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13854_ net1228 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ _04423_ _07328_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_18_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16573_ clknet_leaf_94_wb_clk_i _02697_ _01380_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_13785_ net2714 _03275_ net960 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10997_ net668 _06508_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15524_ clknet_leaf_1_wb_clk_i _01664_ _00332_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12736_ _06823_ _06851_ _06873_ _06901_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08915__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12945__B _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15455_ clknet_leaf_111_wb_clk_i _01595_ _00263_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12437__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12667_ net358 net2176 net434 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14406_ net1075 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11618_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04347_ net952 _07105_ vssd1
+ vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15386_ clknet_leaf_121_wb_clk_i _01526_ _00194_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09613__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12598_ net331 net2373 net440 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__mux2_1
XANTENNA__08967__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14337_ net1211 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11549_ net421 _06666_ _07038_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold507 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold518 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold529 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ net1148 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16007_ clknet_leaf_26_wb_clk_i _02147_ _00815_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13219_ net626 net937 net1018 net1663 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12172__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ net1173 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire549_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10931__C1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1207 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15704__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08760_ net848 _04364_ _04370_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1218 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07711_ _03302_ net425 _03398_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09144__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08691_ net1057 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _04320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07642_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] _03360_ _03334_ vssd1 vssd1
+ vccd1 vccd1 _03365_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07573_ net2660 net190 _00017_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09312_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\] net759 net751 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\]
+ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09852__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09243_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\] net907 vssd1 vssd1
+ vccd1 vccd1 _04760_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12347__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13032__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09174_ _04684_ _04690_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__nor2_2
XFILLER_0_127_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__inv_2
XANTENNA__13967__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1140_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15234__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__A2 _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__A team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _03734_ _03756_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__xor2_2
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout698_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12082__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10391__A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11175__C1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__A2 _04608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09383__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput105 wbs_we_i vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XANTENNA__15384__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\] net777 net712 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\]
+ _04474_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__a221o_1
XANTENNA__09135__A2 _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07909_ _03622_ _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__and2_1
X_08889_ net6 net1029 net987 net1713 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10920_ net392 _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ team_02_WB.instance_to_wrap.top.pc\[30\] _06271_ vssd1 vssd1 vccd1 vccd1
+ _06367_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ net1047 net1050 _03290_ _03103_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__and4b_1
X_10782_ _05534_ net402 vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__nor2_1
XANTENNA__09843__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12765__B _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12521_ net284 net2560 net448 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12257__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15240_ clknet_leaf_70_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[31\]
+ _00053_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12452_ net276 net2392 net450 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11403_ net423 _06450_ _06900_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__o21a_1
X_15171_ net1241 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12383_ net261 net2076 net459 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ net1142 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11334_ net999 _06834_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15727__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14053_ net1128 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11265_ _05980_ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__xnor2_1
X_13004_ _07461_ _07523_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__nor2_1
X_10216_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\] net674 _05729_ _05732_
+ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a211o_1
XANTENNA__09374__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11196_ _05041_ net665 _06700_ _06105_ _06701_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16803__1347 vssd1 vssd1 vccd1 vccd1 _16803__1347/HI net1347 sky130_fd_sc_hd__conb_1
X_10147_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\] net789 net745 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\]
+ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__a221o_1
XANTENNA__15877__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09126__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14955_ net1200 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
X_10078_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\] net924 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a22o_1
X_13906_ net1217 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
XANTENNA__10141__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14886_ net1074 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
XANTENNA__08885__B2 team_02_WB.instance_to_wrap.ramload\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_76_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13837_ net1232 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16625_ clknet_leaf_97_wb_clk_i _02744_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16556_ clknet_leaf_92_wb_clk_i _02680_ _01363_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_13768_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] _03263_
+ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09834__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15507_ clknet_leaf_53_wb_clk_i _01647_ _00315_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12719_ _06713_ _06741_ _06781_ _07242_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__nand4_1
X_16487_ clknet_leaf_72_wb_clk_i net1566 _01295_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12167__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13699_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\] _03221_ vssd1 vssd1 vccd1
+ vccd1 _03222_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15438_ clknet_leaf_8_wb_clk_i _01578_ _00246_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_wire499_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15369_ clknet_leaf_76_wb_clk_i _01509_ _00182_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[28\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_83_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold304 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 _02611_ vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold326 team_02_WB.START_ADDR_VAL_REG\[12\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold337 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold348 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09930_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\] net835 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a22o_1
Xhold359 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16652__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout806 net808 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__buf_4
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09365__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout817 _04520_ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_8
X_09861_ _05355_ _05376_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout828 _04512_ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_4
XFILLER_0_123_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout839 net842 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__buf_6
X_08812_ net116 net1043 net992 net1496 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a22o_1
XANTENNA__12630__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1004 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\] net766 net750 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a22o_1
Xhold1015 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1026 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08743_ _04302_ net847 _04364_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__and3_4
Xhold1037 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1059 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08325__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A _06686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ team_02_WB.instance_to_wrap.top.a1.instruction\[4\] net1061 _04301_ _04302_
+ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__and4_1
XFILLER_0_95_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07625_ _03324_ _03327_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12866__A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1188_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ team_02_WB.instance_to_wrap.Ren vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__inv_2
XANTENNA__09825__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12077__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1296_A team_02_WB.instance_to_wrap.ramstore\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_91_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09226_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\] net711 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__a22o_1
XANTENNA__16182__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09157_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\] net929 net901 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08108_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09088_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\] net863 net856 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13137__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08039_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03744_ _03750_ vssd1 vssd1
+ vccd1 vccd1 _03761_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold860 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net1000 _06560_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__nor2_1
Xhold893 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10001_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\] net784 net756 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a22o_1
XANTENNA__10371__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09108__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14740_ net1076 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11952_ net276 net2166 net585 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _06136_ _06137_ _06239_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14671_ net1115 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
X_11883_ net280 net2504 net488 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ clknet_leaf_66_wb_clk_i _02545_ _01218_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08973__B net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13622_ team_02_WB.instance_to_wrap.top.a1.row1\[3\] _03119_ _03126_ team_02_WB.instance_to_wrap.top.a1.row2\[3\]
+ _03159_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ net546 net372 vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09816__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16525__CLK clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16341_ clknet_leaf_50_wb_clk_i _02481_ _01149_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13553_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__nand2b_1
X_10765_ net947 _06124_ _06276_ net608 vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__o211a_2
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12504_ net360 net1940 net559 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16272_ clknet_leaf_39_wb_clk_i _02412_ _01080_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13484_ team_02_WB.START_ADDR_VAL_REG\[24\] _04260_ vssd1 vssd1 vccd1 vccd1 net208
+ sky130_fd_sc_hd__and2_1
X_10696_ team_02_WB.instance_to_wrap.top.pc\[16\] _06192_ vssd1 vssd1 vccd1 vccd1
+ _06213_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15223_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[14\]
+ _00036_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_12435_ net343 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\] net456 vssd1
+ vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09595__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15154_ net1244 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12366_ net334 net1812 net563 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14105_ net1137 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11317_ net521 net406 _06065_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__a21o_1
X_15085_ net1235 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
X_12297_ net319 net2230 net569 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__mux2_1
X_14036_ net1076 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
X_11248_ net373 _06503_ _06506_ net377 vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12450__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11179_ net946 _06679_ _06685_ net608 vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__o211a_2
XANTENNA__09325__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16055__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15987_ clknet_leaf_57_wb_clk_i _02127_ _00795_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13300__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10114__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14938_ net1182 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
XANTENNA__11311__C1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14869_ net1216 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16608_ clknet_leaf_80_wb_clk_i _02727_ _01401_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_08390_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__inv_2
XANTENNA__09807__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16539_ clknet_leaf_93_wb_clk_i _02666_ _01346_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09995__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09011_ _04295_ _04297_ net951 vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__nand3_4
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12625__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold101 team_02_WB.instance_to_wrap.top.a1.row1\[112\] vssd1 vssd1 vccd1 vccd1 net1559
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold112 _02578_ vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold123 team_02_WB.instance_to_wrap.top.a1.row1\[8\] vssd1 vssd1 vccd1 vccd1 net1581
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 team_02_WB.instance_to_wrap.ramstore\[12\] vssd1 vssd1 vccd1 vccd1 net1592
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold145 _02569_ vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 team_02_WB.instance_to_wrap.top.a1.row1\[3\] vssd1 vssd1 vccd1 vccd1 net1614
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 net155 vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09338__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold178 team_02_WB.START_ADDR_VAL_REG\[30\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\] net732 _05427_ _05429_
+ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout603 _07189_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_8
Xhold189 net112 vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout396_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout647 _04452_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12360__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\] net855 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\]
+ _05360_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__a221o_1
XANTENNA__14141__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout658 net660 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1103_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10353__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 _05965_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_4
X_09775_ net610 _05290_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout563_A _07219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ _04344_ _04349_ _04354_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_55_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10105__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09510__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] net997 vssd1 vssd1 vccd1
+ vccd1 _04286_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_16_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout730_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07608_ _03324_ _03328_ team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1
+ vccd1 vccd1 _03331_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08588_ net104 net71 net105 vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ net391 _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__or2_1
X_16802__1346 vssd1 vssd1 vccd1 vccd1 _16802__1346/HI net1346 sky130_fd_sc_hd__conb_1
XFILLER_0_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09209_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\] net886 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12535__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481_ net389 _05876_ _05995_ _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12220_ net2266 net280 net617 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09577__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10563__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08785__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ net265 net1873 net463 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11102_ net416 _06053_ net382 _06101_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__a22o_1
XANTENNA__09329__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12082_ net2011 net258 net583 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold690 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11136__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15910_ clknet_leaf_42_wb_clk_i _02050_ _00718_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11033_ net369 _06478_ _06543_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12270__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16890_ net1434 vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__buf_2
XANTENNA__11687__A3 _04608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15841_ clknet_leaf_122_wb_clk_i _01981_ _00649_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15772_ clknet_leaf_47_wb_clk_i _01912_ _00580_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _07486_ _07503_ _07485_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08984__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09501__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14723_ net1145 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
X_11935_ net356 net2621 net482 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14654_ net1191 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
X_11866_ net341 net2367 net493 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13605_ net2207 net962 _03157_ net1065 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__o211a_1
X_10817_ _05103_ net404 vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__or2_1
XANTENNA__08068__A2 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14585_ net1137 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13061__A2 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11797_ net337 net2728 net596 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__mux2_1
X_13536_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] _03061_ _03092_ _03095_
+ net1067 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__o221a_1
X_16324_ clknet_leaf_1_wb_clk_i _02464_ _01132_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10748_ team_02_WB.instance_to_wrap.top.pc\[20\] _06264_ vssd1 vssd1 vccd1 vccd1
+ _06265_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16255_ clknet_leaf_87_wb_clk_i _02395_ _01063_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13467_ team_02_WB.START_ADDR_VAL_REG\[7\] net1069 net1003 vssd1 vssd1 vccd1 vccd1
+ net221 sky130_fd_sc_hd__a21o_1
XANTENNA__12445__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10679_ net994 _05785_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ clknet_leaf_74_wb_clk_i _01418_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.debounce
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12418_ net281 net2013 net456 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09568__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16186_ clknet_leaf_118_wb_clk_i _02326_ _00994_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13398_ net2755 net1012 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[27\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput206 net206 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput217 net217 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ net1247 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
X_12349_ net267 net2666 net561 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ net1262 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15057__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ net1133 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12180__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07890_ _03575_ _03609_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__xor2_1
XANTENNA__10335__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15445__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09740__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire629_A _05289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15207__D net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09560_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\] net801 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08511_ team_02_WB.instance_to_wrap.top.a1.data\[6\] net958 vssd1 vssd1 vccd1 vccd1
+ _04202_ sky130_fd_sc_hd__or2_1
X_09491_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\] net720 _05005_ _05006_
+ _05007_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_76_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08700__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08442_ _04135_ _04138_ _04142_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08373_ _04078_ _04080_ _04082_ _04076_ _04075_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__o311a_1
XFILLER_0_110_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout311_A _06840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08988__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12355__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1053_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout409_A _05809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09559__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08767__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1161_A team_02_WB.instance_to_wrap.ramaddr\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16220__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13975__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1220_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout680_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 net401 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_2
XFILLER_0_111_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout778_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _05715_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_2
XANTENNA__12090__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout433 _07229_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_6
XANTENNA__10326__B1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout455 net457 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_4
Xfanout466 net469 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09192__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout477 _07206_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
X_09827_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\] net738 net730 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09731__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 _07198_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_8
XANTENNA_fanout945_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15938__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\] net903 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08709_ net651 net932 _04337_ _04286_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_69_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09689_ net968 _05205_ _04497_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10839__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11720_ net303 net2494 net603 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11651_ net666 _07127_ _07136_ _06583_ _07131_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__o221a_1
XFILLER_0_83_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13043__A2 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11054__A1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ net547 _06117_ _04567_ net659 vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_65_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09798__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14370_ net1207 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
X_11582_ _06040_ _06045_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13321_ net1063 _04180_ _04231_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__or3_2
X_10533_ _06048_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12265__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10574__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ clknet_leaf_18_wb_clk_i _02180_ _00848_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13252_ team_02_WB.instance_to_wrap.top.pc\[30\] net1054 _02968_ _02971_ vssd1 vssd1
+ vccd1 vccd1 _02972_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input74_A wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ _04885_ _04905_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__nor2_1
XANTENNA__08044__A team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12203_ net339 net2471 net579 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183_ net977 _07397_ _02942_ _07066_ net232 vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__o32a_1
X_10395_ _05738_ _05911_ _05736_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12134_ net333 net2287 net467 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
XANTENNA__09970__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08698__B net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10317__A0 _05785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ net323 net1637 net472 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09183__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ _06147_ net655 net495 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] net497
+ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__a221o_1
XANTENNA__09722__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16873_ net1417 vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_105_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15824_ clknet_leaf_40_wb_clk_i _01964_ _00632_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12967_ team_02_WB.instance_to_wrap.top.pc\[6\] _05671_ vssd1 vssd1 vccd1 vccd1 _07487_
+ sky130_fd_sc_hd__xnor2_1
X_15755_ clknet_leaf_114_wb_clk_i _01895_ _00563_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13282__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14706_ net1123 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
XANTENNA__10096__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ net279 net1839 net483 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15686_ clknet_leaf_44_wb_clk_i _01826_ _00494_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12898_ _05271_ _06197_ _07417_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_64_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11849_ net282 net1926 net491 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
X_14637_ net1147 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11045__A1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14568_ net1175 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16307_ clknet_leaf_52_wb_clk_i _02447_ _01115_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13519_ _03074_ _03076_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12175__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14499_ net1134 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XANTENNA__08461__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16238_ clknet_leaf_27_wb_clk_i _02378_ _01046_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16169_ clknet_leaf_104_wb_clk_i _02309_ _00977_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08991_ net943 _04503_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__and3_1
XANTENNA__09961__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07942_ _03634_ _03637_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07873_ _03556_ _03586_ _03587_ _03591_ _03595_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__o311ai_4
XTAP_TAPCELL_ROW_121_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13019__B _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16801__1345 vssd1 vssd1 vccd1 vccd1 _16801__1345/HI net1345 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_3_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11520__A2 _07007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09612_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\] net712 net676 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\]
+ _05128_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09543_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\] net770 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout261_A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13273__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_A _07069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09474_ net971 _04990_ net544 vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04119_ _04125_ _04118_ vssd1
+ vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__o31a_1
XFILLER_0_59_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12874__A _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1170_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _04055_ _04058_ _04050_ _04051_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_24_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08287_ _03966_ _04001_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12085__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout895_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11339__A2 _06830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10180_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\] net825 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15760__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1212 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__clkbuf_4
Xfanout1217 net1225 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__clkbuf_4
Xfanout1228 net1229 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__buf_4
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout241 _06282_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09165__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1239 net1250 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__buf_4
XANTENNA__09704__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout252 net254 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
Xfanout263 _06595_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_2
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_2
Xfanout285 net287 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
Xfanout296 net299 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
X_13870_ net1231 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16116__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ _03318_ _07342_ _07339_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__a21o_1
XANTENNA__13264__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10078__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ _05938_ _05952_ _05958_ _07275_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__or4_1
X_15540_ clknet_leaf_13_wb_clk_i _01680_ _00348_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11275__B2 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08039__A team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11703_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] _04333_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__or3b_2
X_15471_ clknet_leaf_38_wb_clk_i _01611_ _00279_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12683_ net276 net1983 net431 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08981__B net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ net1093 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
X_11634_ net656 _07112_ _07120_ net795 vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11578__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14353_ net1106 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
Xwire620 _07215_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11565_ net392 _06979_ _07054_ net381 vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__o211a_1
Xwire631 net632 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13304_ net1549 net986 net967 _03001_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__a22o_1
X_10516_ _05966_ _06032_ _05967_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a21boi_1
XANTENNA__10250__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14284_ net1073 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11496_ team_02_WB.instance_to_wrap.top.pc\[8\] _06256_ vssd1 vssd1 vccd1 vccd1 _06990_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13235_ net1054 team_02_WB.instance_to_wrap.top.ru.state\[0\] net985 vssd1 vssd1
+ vccd1 vccd1 _02957_ sky130_fd_sc_hd__o21ba_2
X_16023_ clknet_leaf_14_wb_clk_i _02163_ _00831_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10447_ _04462_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10002__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13166_ _07486_ _07503_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10378_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\] net914 _05893_ _05894_
+ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a211o_1
X_12117_ net264 net2365 net466 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__mux2_1
X_13097_ net1027 _02871_ net1024 team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1
+ vccd1 vccd1 _01500_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09156__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ net249 net2633 net470 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16856_ net1400 vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15807_ clknet_leaf_86_wb_clk_i _01947_ _00615_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16787_ net1331 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
X_13999_ net1115 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
XANTENNA__10069__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ clknet_leaf_121_wb_clk_i _01878_ _00546_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15669_ clknet_leaf_43_wb_clk_i _01809_ _00477_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15070__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11802__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08210_ net2214 net1007 net982 _03927_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XANTENNA__11018__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09190_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\] net770 _04703_ _04704_
+ _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a2111o_1
XANTENNA__15633__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08141_ _03849_ _03859_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08072_ _03790_ _03792_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__nor2_1
XANTENNA__10241__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12633__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09395__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08412__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap997 _04275_ vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] net790 vssd1 vssd1 vccd1
+ vccd1 _04491_ sky130_fd_sc_hd__or2_2
XFILLER_0_23_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 team_02_WB.instance_to_wrap.ramstore\[25\] vssd1 vssd1 vccd1 vccd1 net1474
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09147__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold27 _00010_ vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03636_ vssd1 vssd1 vccd1
+ vccd1 _03648_ sky130_fd_sc_hd__xnor2_2
Xhold38 team_02_WB.instance_to_wrap.ramaddr\[19\] vssd1 vssd1 vccd1 vccd1 net1496
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_02_WB.instance_to_wrap.top.a1.data\[5\] vssd1 vssd1 vccd1 vccd1 net1507
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout476_A _07206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ _03544_ net329 vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07787_ _03507_ _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16289__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout643_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09526_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\] net766 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\] net806 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout810_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11712__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ _04108_ _04111_ _04102_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09388_ net968 _04904_ _04497_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08339_ _04022_ _04038_ _04027_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10232__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11350_ net374 _06631_ _06849_ net383 vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10301_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\] net740 net676 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a22o_1
X_11281_ _06215_ _06216_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12543__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13020_ _07445_ _07538_ _07539_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09386__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\] net831 net924 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\]
+ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10571__B net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11159__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\] net901 net881 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__a22o_1
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1014 team_02_WB.instance_to_wrap.top.ru.next_iready vssd1 vssd1 vccd1 vccd1
+ net1014 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10940__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1025 _07348_ vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__buf_2
XANTENNA__09138__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1036 _04428_ vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__buf_2
XANTENNA_input37_A gpio_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 team_02_WB.instance_to_wrap.top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1
+ net1047 sky130_fd_sc_hd__clkbuf_2
X_10094_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\] net769 net677 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\]
+ _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__a221o_1
XANTENNA__09689__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14971_ net1257 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
Xfanout1058 net1059 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13485__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15506__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1069 net1070 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_2
X_16710_ net1269 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13922_ net1219 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
XANTENNA__10299__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16641_ clknet_leaf_102_wb_clk_i _02760_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_13853_ net1226 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
X_12804_ _05835_ _05876_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__xnor2_1
X_16572_ clknet_leaf_93_wb_clk_i net1770 _01379_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13784_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] _03275_
+ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__and2_1
X_10996_ net424 _06504_ _06507_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__o21a_1
XANTENNA__15656__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15523_ clknet_leaf_2_wb_clk_i _01663_ _00331_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12735_ _06943_ _06963_ _06982_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12666_ net343 net2355 net437 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__mux2_1
X_15454_ clknet_leaf_114_wb_clk_i _01594_ _00262_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14405_ net1094 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
X_11617_ net1001 net973 team_02_WB.instance_to_wrap.top.pc\[2\] vssd1 vssd1 vccd1
+ vccd1 _07105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15385_ clknet_leaf_17_wb_clk_i _01525_ _00193_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12597_ net335 net2017 net440 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__mux2_1
X_16800__1344 vssd1 vssd1 vccd1 vccd1 _16800__1344/HI net1344 sky130_fd_sc_hd__conb_1
XFILLER_0_108_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11548_ net421 _06673_ _07038_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__o21ai_1
X_14336_ net1151 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12961__B _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold508 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap227 _03788_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_1
XANTENNA__12453__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14267_ net1159 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
Xhold519 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11479_ team_02_WB.instance_to_wrap.top.pc\[9\] net973 _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\]
+ _06973_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap539_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16006_ clknet_leaf_44_wb_clk_i _02146_ _00814_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13218_ net629 net936 net1020 net1744 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09377__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09916__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198_ net1138 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
XANTENNA__07927__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13149_ net228 _02913_ _02914_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09129__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1208 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13476__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] _03398_ net425 vssd1 vssd1
+ vccd1 vccd1 _03433_ sky130_fd_sc_hd__or3b_1
X_08690_ _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08352__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire611_A _05270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07641_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] _03360_ vssd1 vssd1 vccd1
+ vccd1 _03364_ sky130_fd_sc_hd__xnor2_2
X_16839_ net1383 vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_2
XFILLER_0_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07572_ _03310_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09301__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09311_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\] net771 net735 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a22o_1
XANTENNA__16581__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12628__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09242_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\] net822 net919 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\]
+ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09173_ _04686_ _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__or3_1
XANTENNA__13125__A1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08124_ _03778_ _03805_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10214__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12871__B _05828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ _03720_ _03772_ _03773_ _03715_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__12363__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1133_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09907__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13164__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11175__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10391__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout760_A _04374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\] net737 net689 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout858_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ _03626_ _03629_ _03630_ _03628_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_93_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08888_ net7 net1031 net989 net2098 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a22o_1
XANTENNA__09540__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07839_ _03521_ _03553_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08894__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10850_ _06132_ _06240_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09509_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\] net884 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12538__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ _05579_ net384 vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ net275 net1919 net446 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12451_ net283 net2225 net451 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11402_ net374 _06691_ _06899_ net380 vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__o22a_1
XANTENNA__10205__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15170_ net1242 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
X_12382_ net265 net2313 net459 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11402__B2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14121_ net1112 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11333_ team_02_WB.instance_to_wrap.top.pc\[15\] _06261_ vssd1 vssd1 vccd1 vccd1
+ _06834_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12273__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14052_ net1130 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11264_ _05211_ _06016_ _05208_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13003_ _07462_ _07522_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__nor2_1
XANTENNA__13893__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\] net786 _05730_ _05731_
+ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08031__B1 _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ _05040_ net659 _06113_ _05038_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08987__A team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\] net761 net709 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10077_ _05587_ _05589_ _05591_ _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__or4_1
X_14954_ net1139 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09531__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ net1252 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
X_14885_ net1085 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
X_16624_ clknet_leaf_96_wb_clk_i _02743_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13836_ net1234 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08926__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16555_ clknet_leaf_92_wb_clk_i _02679_ _01362_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
X_13767_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] _03263_
+ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__and2_1
XANTENNA__12448__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10757__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979_ _06144_ _06145_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15506_ clknet_leaf_3_wb_clk_i _01646_ _00314_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12718_ _06805_ _06828_ _07241_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__and3_1
X_16486_ clknet_leaf_71_wb_clk_i net1521 _01294_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13698_ net1240 _03220_ _03221_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__nor3_1
XANTENNA__10476__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15437_ clknet_leaf_21_wb_clk_i _01577_ _00245_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12649_ net282 net2005 net435 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15368_ clknet_leaf_82_wb_clk_i _01508_ _00181_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09062__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold305 team_02_WB.instance_to_wrap.ramstore\[24\] vssd1 vssd1 vccd1 vccd1 net1763
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ net1111 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12183__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold316 team_02_WB.instance_to_wrap.top.a1.row1\[57\] vssd1 vssd1 vccd1 vccd1 net1774
+ sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ clknet_leaf_67_wb_clk_i _01443_ _00112_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold327 team_02_WB.instance_to_wrap.top.a1.row2\[26\] vssd1 vssd1 vccd1 vccd1 net1785
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold349 team_02_WB.instance_to_wrap.ramload\[2\] vssd1 vssd1 vccd1 vccd1 net1807
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09860_ _05356_ _05376_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__and2_1
Xfanout807 net808 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_8
Xfanout818 _04520_ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_4
Xfanout829 net832 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08573__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15821__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ net118 net1044 net991 net1598 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a22o_1
X_09791_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\] net730 net710 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\]
+ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__a221o_1
Xhold1005 team_02_WB.instance_to_wrap.ramload\[29\] vssd1 vssd1 vccd1 vccd1 net2463
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _04296_ net848 _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__and3_4
Xhold1027 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08673_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__and2_2
XANTENNA__08876__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15971__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07624_ _03328_ _03346_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10683__A2 _05785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09521__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07555_ team_02_WB.instance_to_wrap.Wen vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout341_A _07051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12358__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout439_A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09225_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\] net750 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\]
+ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1250_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12882__A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09589__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\] net836 net800 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09053__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10199__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08107_ _03824_ _03825_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\] net798 _04591_ _04603_
+ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12093__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08800__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08038_ _03744_ _03750_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1
+ vccd1 vccd1 _03760_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold850 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout975_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold872 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11699__A1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold894 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10000_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\] net736 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__a22o_1
XANTENNA__09761__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09989_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\] net920 net900 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11951_ net282 net2301 net586 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10902_ _06136_ _06137_ _06239_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11882_ net269 net2189 net486 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__mux2_1
X_14670_ net1164 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09431__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10833_ net546 net369 vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__nor2_1
X_13621_ team_02_WB.instance_to_wrap.top.a1.row1\[59\] _03117_ _03123_ team_02_WB.instance_to_wrap.top.a1.row2\[43\]
+ _03158_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_120_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13073__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12268__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09816__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16340_ clknet_leaf_12_wb_clk_i _02480_ _01148_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10764_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _06278_ _06280_ _04334_
+ team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__o311a_1
X_13552_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] net1048 vssd1 vssd1 vccd1
+ vccd1 _03107_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09292__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13888__A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12503_ net355 net1918 net559 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__mux2_1
X_16271_ clknet_leaf_38_wb_clk_i _02411_ _01079_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13483_ team_02_WB.START_ADDR_VAL_REG\[23\] net1070 net1003 vssd1 vssd1 vccd1 vccd1
+ net207 sky130_fd_sc_hd__a21o_1
XFILLER_0_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10695_ _06198_ _06209_ _06211_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11900__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15222_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[13\]
+ _00035_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_12434_ net338 net2302 net457 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__mux2_1
XANTENNA__09044__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12365_ net327 net2362 net563 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__mux2_1
X_15153_ net1249 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14104_ net1193 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
X_11316_ _05988_ _06816_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__xnor2_1
X_15084_ net1253 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12296_ net312 net1913 net569 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14035_ net1165 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ net421 _06750_ _06355_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__a21boi_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09606__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net999 _06683_ _06684_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10129_ _05627_ net649 net968 vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__mux2_2
X_15986_ clknet_leaf_11_wb_clk_i _02126_ _00794_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09504__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13300__A1 team_02_WB.instance_to_wrap.ramaddr\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13300__B2 _02999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14937_ net1139 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14868_ net1076 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16607_ clknet_leaf_80_wb_clk_i _02726_ _01400_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_13819_ net1226 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__inv_2
XANTENNA__12178__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14799_ net1116 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07818__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16538_ clknet_leaf_93_wb_clk_i _02665_ _01345_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[61\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09283__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16469_ clknet_leaf_93_wb_clk_i net1583 _01277_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
X_09010_ _04295_ net951 vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__nand2_1
XANTENNA__11810__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09035__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold102 team_02_WB.instance_to_wrap.top.a1.row1\[113\] vssd1 vssd1 vccd1 vccd1 net1560
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold113 net185 vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07597__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10050__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold124 net107 vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold135 _02574_ vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold146 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold157 net160 vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _02586_ vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\] net756 net845 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\]
+ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__a221o_1
XANTENNA__12641__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout604 _07189_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_2
XANTENNA__09743__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\] net890 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__a22o_1
Xfanout659 net660 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_2
XANTENNA_fanout291_A _06712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09774_ _05271_ _05290_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_124_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ net651 net932 _04351_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _04274_ _04279_ _04280_ net976 vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07607_ _03324_ _03328_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08587_ _04244_ _04247_ _04248_ net1055 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__o22a_1
XANTENNA__12088__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15717__CLK clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09274__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11081__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11720__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09208_ _04718_ _04720_ _04722_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ _05996_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__inv_2
XANTENNA__15867__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09139_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\] net733 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\]
+ _04655_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12150_ net256 net1828 net463 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__mux2_1
XANTENNA__09982__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11101_ net424 _06069_ net413 vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12081_ net1941 net250 net581 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
XANTENNA__12551__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold680 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ net390 _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15840_ clknet_leaf_107_wb_clk_i _01980_ _00648_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ clknet_leaf_126_wb_clk_i _01911_ _00579_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _03295_ _05671_ _07502_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_107_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14722_ net1206 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15163__A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934_ net342 net2222 net485 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15397__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14653_ net1084 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
X_11865_ net339 net1954 net493 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_107_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13604_ team_02_WB.instance_to_wrap.top.a1.row2\[26\] _03118_ _03150_ _03156_ vssd1
+ vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__a211o_1
X_10816_ net525 net404 vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__nand2_1
X_14584_ net1215 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11796_ net330 net2022 net595 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16323_ clknet_leaf_125_wb_clk_i _02463_ _01131_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13535_ _03076_ _03084_ _03093_ _03094_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__or4_1
XANTENNA__11072__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10747_ team_02_WB.instance_to_wrap.top.pc\[19\] team_02_WB.instance_to_wrap.top.pc\[18\]
+ _06263_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10280__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16254_ clknet_leaf_113_wb_clk_i _02394_ _01062_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10678_ team_02_WB.instance_to_wrap.top.pc\[15\] _06194_ vssd1 vssd1 vccd1 vccd1
+ _06195_ sky130_fd_sc_hd__nand2_1
X_13466_ team_02_WB.START_ADDR_VAL_REG\[6\] net1068 net1002 vssd1 vssd1 vccd1 vccd1
+ net220 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_11_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08346__A2_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15205_ clknet_leaf_78_wb_clk_i net1463 _00019_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.edg2.flip2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12417_ net270 net2474 net454 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__mux2_1
X_16185_ clknet_leaf_17_wb_clk_i _02325_ _00993_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13397_ team_02_WB.instance_to_wrap.ramload\[26\] net1012 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[26\] sky130_fd_sc_hd__and2_1
XFILLER_0_84_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput207 net207 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput218 net218 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
X_15136_ net1230 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12348_ net258 net1936 net562 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11780__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16022__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15067_ net1258 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
XANTENNA__12461__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net238 net1801 net569 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__mux2_1
XANTENNA__14242__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ net1205 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire524_A _05186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15969_ clknet_leaf_121_wb_clk_i _02109_ _00777_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08510_ _04201_ net1613 _04186_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15073__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09490_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\] net772 net728 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08441_ _04135_ _04142_ _04138_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a21oi_2
XANTENNA__13037__B1 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08372_ _04080_ _04082_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08464__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12636__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13321__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10023__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12371__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1213_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _05808_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_2
XANTENNA__09716__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout412 _05763_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout423 net424 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout434 net437 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout445 _07225_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout456 net457 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_35_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\] net726 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\]
+ _05337_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_35_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout467 net469 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_8
Xfanout478 net481 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_35_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout489 _07198_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_4
X_09757_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\] net834 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\]
+ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a221o_1
XANTENNA__13276__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout938_A _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11715__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ _04271_ _04336_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09688_ _05198_ _05201_ _05202_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__or4_4
XFILLER_0_55_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09495__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08639_ net1062 net1060 _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__or3_4
XFILLER_0_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11650_ net424 _06797_ _07134_ _07135_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__inv_2
X_11581_ net365 _07033_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__nor2_1
XANTENNA__12546__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13320_ net1486 net985 net966 _03009_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__a22o_1
XANTENNA__10262__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10532_ _05579_ net402 vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10574__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16045__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13251_ _06365_ _02965_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__or2_1
X_10463_ _05167_ _05168_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__and2b_2
XFILLER_0_122_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10014__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09955__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ net332 net2162 net579 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__mux2_1
X_13182_ _07388_ _07395_ _07396_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__and3_1
X_10394_ _05906_ _05909_ _05783_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input67_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10565__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ net325 net2156 net467 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
XANTENNA__12281__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15158__A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10590__A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14062__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09707__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ net317 net2129 net470 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11015_ net1000 _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_109_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16872_ net1416 vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__buf_2
XFILLER_0_99_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout990 net991 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
X_15823_ clknet_leaf_38_wb_clk_i _01963_ _00631_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13267__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15754_ clknet_leaf_130_wb_clk_i _01894_ _00562_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12966_ team_02_WB.instance_to_wrap.top.pc\[7\] _05627_ vssd1 vssd1 vccd1 vccd1 _07486_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__09486__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ net1106 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11917_ net282 net2064 net483 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ clknet_leaf_34_wb_clk_i _01825_ _00493_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _07374_ _07375_ _07416_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14636_ net1080 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ net270 net2577 net490 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14567_ net1117 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12456__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11779_ net262 net2744 net594 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ clknet_leaf_6_wb_clk_i _02446_ _01114_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13518_ _03077_ _03078_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14498_ net1210 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16237_ clknet_leaf_24_wb_clk_i _02377_ _01045_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13449_ _03052_ _03053_ _03041_ _03048_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_45_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_75_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10005__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11202__C1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16168_ clknet_leaf_19_wb_clk_i _02308_ _00976_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15119_ net1104 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12191__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__and3b_2
XFILLER_0_80_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16099_ clknet_leaf_13_wb_clk_i _02239_ _00907_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_07941_ _03641_ _03662_ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15562__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _03592_ _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08921__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\] net784 net736 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09542_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\] net742 _05044_ _05058_
+ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09473_ _04980_ _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_138_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout254_A _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08424_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04125_ vssd1 vssd1 vccd1
+ vccd1 _04131_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_138_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09229__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12874__B _05781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ _04051_ _04065_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__xor2_2
XFILLER_0_74_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12366__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1163_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ _03962_ _03988_ _03979_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09937__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout790_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08799__B _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A _04536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15905__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1207 net1209 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_4
Xfanout1218 net1219 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__buf_4
Xfanout1229 net1230 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__buf_4
Xfanout231 _07333_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
Xfanout242 _06282_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
Xfanout253 net254 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout264 net267 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_2
XANTENNA__14610__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 _06740_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08912__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout297 net299 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlymetal6s2s_1
X_09809_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\] net886 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__a22o_1
XANTENNA__08912__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13249__B1 _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12820_ _03318_ _07342_ _07339_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09468__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11275__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12751_ _04780_ _05933_ _07272_ _07274_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__or4_1
XANTENNA__08140__A2 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11702_ net2562 net346 net642 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15470_ clknet_leaf_26_wb_clk_i _01610_ _00278_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12682_ net281 net2202 net431 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ net1185 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ net422 _06774_ _07111_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__o21a_1
XANTENNA__08428__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11180__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10235__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15435__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14352_ net1091 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_8
Xwire621 _05713_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_2
X_11564_ net407 _07053_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__or2_1
Xwire632 _05079_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09640__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ team_02_WB.instance_to_wrap.top.pc\[8\] net1051 _06989_ net933 vssd1 vssd1
+ vccd1 vccd1 _03001_ sky130_fd_sc_hd__a22o_2
X_10515_ _04695_ _06031_ net542 _04692_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_108_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11495_ net671 _06976_ _06988_ net673 _06987_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__a221o_2
XFILLER_0_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14283_ net1151 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
X_16022_ clknet_leaf_48_wb_clk_i _02162_ _00830_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13234_ net1055 team_02_WB.instance_to_wrap.top.ru.state\[2\] net1022 _00011_ vssd1
+ vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a211o_2
XFILLER_0_21_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10446_ _04464_ _04467_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__nand2_2
XFILLER_0_126_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10377_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\] net886 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\]
+ _05885_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a221o_1
X_13165_ _07404_ _07406_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12116_ net257 net1986 net468 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__mux2_1
X_13096_ _06735_ net233 _02868_ net978 _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12047_ net253 net1910 net473 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12959__B _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16855_ net1399 vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_122_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15806_ clknet_leaf_118_wb_clk_i _01946_ _00614_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16786_ net1330 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13998_ net1095 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
XANTENNA__09459__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15737_ clknet_leaf_112_wb_clk_i _01877_ _00545_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12949_ team_02_WB.instance_to_wrap.top.pc\[16\] _06194_ vssd1 vssd1 vccd1 vccd1
+ _07469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15668_ clknet_leaf_12_wb_clk_i _01808_ _00476_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11018__A2 _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14619_ net1184 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12186__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15599_ clknet_leaf_34_wb_clk_i _01739_ _00407_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08140_ net2240 net1007 net982 net226 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10226__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10777__A1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09631__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07642__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08071_ _03769_ _03791_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_126_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15928__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09919__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08973_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] net791 vssd1 vssd1 vccd1
+ vccd1 _04490_ sky130_fd_sc_hd__nor2_8
XANTENNA__13479__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold17 _02587_ vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07924_ _03615_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__xor2_2
Xhold28 team_02_WB.instance_to_wrap.ramaddr\[0\] vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold39 _02613_ vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12869__B _05828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] _03575_ _03576_ _03577_ vssd1
+ vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout371_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A _07211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09243__B net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07786_ _03473_ _03497_ _03508_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12885__A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09456_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\] net826 net883 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\]
+ _04972_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_26_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09870__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _04102_ _04108_ _04111_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__nand3_1
XANTENNA__12096__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout803_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ _04897_ _04900_ _04902_ _04903_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_95_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10217__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08338_ _04021_ _04048_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__xnor2_4
XANTENNA__09083__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09622__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08269_ _03919_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08830__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10300_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\] net841 _05813_ _05814_
+ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_105_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ net952 _06782_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10231_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\] net876 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12390__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\] net807 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\]
+ _05678_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_89_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1004 _04259_ vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1015 team_02_WB.instance_to_wrap.top.ru.next_iready vssd1 vssd1 vccd1 vccd1
+ net1015 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_89_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1026 _07338_ vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_4
X_10093_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\] net744 net729 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__a22o_1
Xfanout1037 net1038 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
X_14970_ net1247 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
Xfanout1048 team_02_WB.instance_to_wrap.top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1
+ net1048 sky130_fd_sc_hd__clkbuf_2
Xfanout1059 team_02_WB.instance_to_wrap.top.a1.instruction\[12\] vssd1 vssd1 vccd1
+ vccd1 net1059 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09689__A2 _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ net1218 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
XANTENNA__08897__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ clknet_leaf_102_wb_clk_i _02759_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13852_ net1229 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ team_02_WB.instance_to_wrap.top.i_ready net235 vssd1 vssd1 vccd1 vccd1 _07327_
+ sky130_fd_sc_hd__nand2_1
X_16749__1293 vssd1 vssd1 vccd1 vccd1 _16749__1293/HI net1293 sky130_fd_sc_hd__conb_1
X_16571_ clknet_leaf_92_wb_clk_i _02695_ _01378_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13783_ _03275_ net960 _03274_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__and3b_1
XANTENNA__12795__A _06102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08992__B team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10995_ net378 _06505_ _06506_ net373 vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__o22a_1
XANTENNA__11903__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15522_ clknet_leaf_123_wb_clk_i _01662_ _00330_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07889__A team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12734_ _06284_ _07257_ _06414_ _06035_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_84_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15453_ clknet_leaf_49_wb_clk_i _01593_ _00261_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12665_ net338 net1915 net437 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14404_ net1127 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
XANTENNA__10208__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11616_ _07095_ _07096_ _07103_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__o21ai_4
XANTENNA__09074__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15384_ clknet_leaf_51_wb_clk_i _01524_ _00192_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10759__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ net328 net2117 net440 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__mux2_1
XANTENNA__11956__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09613__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14335_ net1183 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11420__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11547_ _06087_ _06870_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08821__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09609__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold509 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ net1186 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11478_ net998 _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16005_ clknet_leaf_32_wb_clk_i _02145_ _00813_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13217_ _05250_ net936 net1020 net1479 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_81_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10429_ _05042_ _05945_ _05038_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14197_ net1215 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13148_ _07480_ _07481_ _07508_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13079_ team_02_WB.instance_to_wrap.top.pc\[22\] net1024 _02856_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1209 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08888__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ _03332_ _03360_ _03362_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__a21oi_1
X_16838_ net1382 vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_2
XFILLER_0_117_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07571_ net37 net36 net35 net34 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__nor4_2
XFILLER_0_18_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16769_ net1313 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15081__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09310_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\] net775 _04825_ _04826_
+ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a211o_1
XANTENNA__11813__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09852__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09241_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\] net915 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15750__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09172_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\] net819 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\]
+ _04673_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a221o_1
XANTENNA__09065__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _03778_ _03805_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08812__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12644__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08054_ _03774_ _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13164__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11175__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10922__A1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\] net701 _04472_ vssd1
+ vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__a21o_1
X_07907_ _03593_ _03624_ _03594_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__a21o_1
X_08887_ net8 net1029 net987 net1580 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout753_A _04376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07838_ _03559_ _03560_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15280__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout920_A _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07769_ _03449_ _03477_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__xor2_1
XANTENNA__11723__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09508_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\] net835 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\]
+ _05024_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10780_ _06288_ _06295_ net396 vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__mux2_2
XANTENNA__09843__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09439_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\] net774 net731 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a22o_1
XANTENNA__10339__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13232__A1_N net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ net270 net2055 net451 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11401_ _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08803__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ net258 net2412 net459 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__mux2_1
XANTENNA__12554__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14120_ net1177 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
X_11332_ net849 _04354_ _06154_ _06832_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__a31o_2
X_14051_ net1130 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11263_ net2697 net284 net643 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13002_ team_02_WB.instance_to_wrap.top.pc\[19\] _06188_ _07521_ vssd1 vssd1 vccd1
+ vccd1 _07522_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10214_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\] net774 net710 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__a22o_1
X_11194_ net421 _06693_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__nand2_1
X_10145_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\] net713 net697 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\]
+ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14953_ net1102 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
X_10076_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] net807 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\]
+ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13904_ net1253 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
X_14884_ net1132 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
XANTENNA__10141__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16623_ clknet_leaf_97_wb_clk_i _02742_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_13835_ net1252 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
XANTENNA__15773__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16554_ clknet_leaf_96_wb_clk_i _02678_ _01361_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13766_ _03263_ _03264_ net961 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__and3b_1
XANTENNA__09295__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ net952 _06490_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__nand2_1
XANTENNA__13091__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15505_ clknet_leaf_51_wb_clk_i _01645_ _00313_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12717_ _06844_ _06882_ _06895_ _07240_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__and4_1
X_16485_ clknet_leaf_71_wb_clk_i _02620_ _01293_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13697_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\]
+ _03217_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15436_ clknet_leaf_25_wb_clk_i _01576_ _00244_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16129__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12648_ net268 net2573 net434 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_109_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15367_ clknet_leaf_82_wb_clk_i _01507_ _00180_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12464__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12579_ net259 net2248 net439 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10773__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14318_ net1113 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15298_ clknet_leaf_82_wb_clk_i _01442_ _00111_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold306 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold317 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13146__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14249_ net1101 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout808 _04534_ vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__buf_4
Xfanout819 _04520_ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_8
X_08810_ net119 net1041 net992 net1703 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a22o_1
XANTENNA__11808__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\] net786 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__a22o_1
Xhold1006 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1017 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08741_ team_02_WB.instance_to_wrap.top.a1.instruction\[16\] net931 team_02_WB.instance_to_wrap.top.a1.instruction\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__and3b_2
Xhold1028 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1039 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
X_08672_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] team_02_WB.instance_to_wrap.top.a1.instruction\[6\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] team_02_WB.instance_to_wrap.top.a1.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__and4_1
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07623_ team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] _03326_ _03330_ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07554_ team_02_WB.instance_to_wrap.top.pc\[6\] vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09286__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09825__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09224_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\] net771 net755 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09038__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09155_ _04656_ _04661_ _04671_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__nor3_2
XANTENNA__12374__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10199__A2 _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08106_ _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09086_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\] net822 net813 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\]
+ _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08037_ _03741_ _03757_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__xnor2_2
X_16748__1292 vssd1 vssd1 vccd1 vccd1 _16748__1292/HI net1292 sky130_fd_sc_hd__conb_1
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11148__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold840 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold851 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15646__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold862 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold884 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout870_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout968_A _04496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ _05498_ _05500_ _05502_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_129_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10371__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08939_ net1001 net996 _04347_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or3_2
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11950_ net268 net2703 net585 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11320__B2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net952 _06415_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__nand2_1
X_11881_ net263 net2721 net488 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
XANTENNA__12549__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13620_ team_02_WB.instance_to_wrap.top.a1.row2\[35\] _03125_ _03128_ team_02_WB.instance_to_wrap.top.a1.row1\[107\]
+ _03171_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_120_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10832_ net410 _06347_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_120_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09816__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13551_ net1047 team_02_WB.instance_to_wrap.top.a1.row2\[12\] _03103_ _03104_ vssd1
+ vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__and4b_1
X_10763_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ _04334_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ net358 net2282 net557 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09029__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16270_ clknet_leaf_26_wb_clk_i _02410_ _01078_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13482_ team_02_WB.START_ADDR_VAL_REG\[22\] _04260_ vssd1 vssd1 vccd1 vccd1 net206
+ sky130_fd_sc_hd__and2_1
XFILLER_0_125_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input97_A wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10694_ _06195_ _06210_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__nand2_1
X_15221_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[12\]
+ _00034_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12433_ net332 net2168 net455 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__mux2_1
XANTENNA__12284__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16421__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15152_ net1247 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
X_12364_ net323 net2730 net563 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14103_ net1172 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
X_11315_ _05295_ _06015_ _05291_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__a21oi_1
X_15083_ net1262 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12295_ net305 net1870 net569 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14034_ net1118 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11246_ _06515_ _06748_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__o21bai_2
XANTENNA__09201__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11177_ net974 _06681_ _06682_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10128_ _05629_ _05640_ _05642_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__nor4_1
XFILLER_0_78_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15985_ clknet_leaf_50_wb_clk_i _02125_ _00793_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13300__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14936_ net1186 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
X_10059_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\] net712 _05573_ _05575_
+ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_19_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10114__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11311__B2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12459__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14867_ net1169 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13818_ net1224 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__inv_2
X_16606_ clknet_leaf_80_wb_clk_i _02725_ _01399_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09268__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14798_ net1114 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
XANTENNA__09807__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16537_ clknet_leaf_93_wb_clk_i _02664_ _01344_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11614__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] _03251_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16468_ clknet_leaf_77_wb_clk_i _02603_ _01276_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15419_ clknet_leaf_1_wb_clk_i _01559_ _00227_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12194__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16399_ clknet_leaf_65_wb_clk_i _02534_ _01207_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15669__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09440__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold103 team_02_WB.instance_to_wrap.ramstore\[31\] vssd1 vssd1 vccd1 vccd1 net1561
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold114 team_02_WB.START_ADDR_VAL_REG\[9\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold125 _02604_ vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12327__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold136 team_02_WB.instance_to_wrap.top.a1.row1\[115\] vssd1 vssd1 vccd1 vccd1 net1594
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 team_02_WB.START_ADDR_VAL_REG\[6\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold158 _02591_ vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09911_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\] net760 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__a22o_1
Xhold169 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1
+ net1627 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12878__A1 _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_4
Xfanout616 net619 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__buf_6
X_09842_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\] net918 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\]
+ _05358_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__a221o_1
XANTENNA__10353__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13038__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ net970 net628 net543 vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _04276_ _04277_ _04352_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_124_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10105__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ net1060 _04283_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__nor2_1
XANTENNA__12369__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1193_A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11273__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07606_ _03324_ _03328_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__and2_1
XANTENNA__09259__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08586_ team_02_WB.instance_to_wrap.wb.curr_state\[0\] _04246_ _04243_ vssd1 vssd1
+ vccd1 vccd1 _04248_ sky130_fd_sc_hd__o21a_1
XANTENNA__13055__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10397__B net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12802__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16444__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout716_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08482__A1 _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09207_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\] net817 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\]
+ _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12566__A0 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09138_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\] net744 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08785__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09069_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\] net738 net711 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14613__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11100_ _06607_ _06608_ net418 vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12080_ net1782 net252 net584 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__mux2_1
Xhold670 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold681 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09734__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11031_ _06073_ _06075_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07745__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13663__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15770_ clknet_leaf_118_wb_clk_i _01910_ _00578_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _07488_ _07501_ _07487_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_107_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13294__B2 _02996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ net1214 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
X_11933_ net340 net2151 net485 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12279__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10588__A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ net1149 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11864_ net330 net2261 net492 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13603_ _03132_ _03152_ _03154_ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__or4_1
XFILLER_0_71_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10815_ net521 net385 _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a21o_1
X_14583_ net1173 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11795_ net335 net1792 net595 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__mux2_1
XANTENNA__11911__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16322_ clknet_leaf_123_wb_clk_i _02462_ _01130_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13534_ _03072_ _03086_ _03081_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__a21oi_1
X_10746_ team_02_WB.instance_to_wrap.top.pc\[17\] _06262_ vssd1 vssd1 vccd1 vccd1
+ _06263_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16253_ clknet_leaf_51_wb_clk_i _02393_ _01061_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13465_ team_02_WB.START_ADDR_VAL_REG\[5\] net1069 net1003 vssd1 vssd1 vccd1 vccd1
+ net219 sky130_fd_sc_hd__a21o_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10677_ net790 _05693_ _06127_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__o22a_2
XFILLER_0_109_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15204_ clknet_leaf_78_wb_clk_i team_02_WB.instance_to_wrap.top.edg2.button_i net1067
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.edg2.flip1 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11212__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12416_ net263 net2565 net456 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16184_ clknet_leaf_22_wb_clk_i _02324_ _00992_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13396_ net1659 net1012 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[25\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09422__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput208 net208 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
X_15135_ net1230 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XANTENNA__08776__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12347_ net248 net2615 net561 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput219 net219 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__15961__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15066_ net1258 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12278_ net244 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\] net570 vssd1
+ vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__mux2_1
XANTENNA__08521__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14017_ net1214 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
X_11229_ team_02_WB.instance_to_wrap.top.pc\[18\] _06263_ team_02_WB.instance_to_wrap.top.pc\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap514_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10335__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11532__A1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16317__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09489__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15968_ clknet_leaf_107_wb_clk_i _02108_ _00776_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14919_ net1122 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
XANTENNA__12189__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15899_ clknet_leaf_127_wb_clk_i _02039_ _00707_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ _04131_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08371_ _04067_ _04073_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__xor2_2
XFILLER_0_129_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11821__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15491__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09661__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09413__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08767__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12652__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14433__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout402 net403 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
Xfanout413 net414 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 _05715_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout435 net437 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11523__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1206_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10326__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 net449 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_6
XFILLER_0_96_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 _07221_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_4
X_09825_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\] net734 net843 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a22o_1
XANTENNA__09192__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout479 net481 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09756_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\] net915 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__a22o_1
X_08707_ net1058 _04277_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09687_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\] net834 net814 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\]
+ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12099__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08638_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04265_ vssd1 vssd1 vccd1
+ vccd1 _04267_ sky130_fd_sc_hd__or2_2
XFILLER_0_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15834__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08569_ _02813_ _04230_ _04180_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11731__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10600_ _04459_ _06114_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__or2_4
XFILLER_0_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ net2450 net356 net642 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09652__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10531_ _05624_ net384 vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13250_ net1573 net985 net966 _02970_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ net528 _05166_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_111_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12201_ net335 net2000 net579 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12562__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13181_ _07492_ _07499_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__xor2_1
X_10393_ _05783_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__nand2_2
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12132_ net324 net2384 net467 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12063_ net313 net2220 net470 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11014_ _06269_ _06525_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__or2_1
XANTENNA__09183__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16871_ net1415 vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__buf_2
XANTENNA__12798__A _07321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout980 _04177_ vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout991 _04427_ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__buf_2
X_15822_ clknet_leaf_27_wb_clk_i _01962_ _00630_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ clknet_leaf_119_wb_clk_i _01893_ _00561_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12965_ _05627_ team_02_WB.instance_to_wrap.top.pc\[7\] vssd1 vssd1 vccd1 vccd1 _07485_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_0_73_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ net268 net2664 net482 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__mux2_1
X_14704_ net1076 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
X_15684_ clknet_leaf_3_wb_clk_i _01824_ _00492_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09891__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12896_ _07415_ _07376_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_64_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14635_ net1150 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ net263 net2700 net491 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ net1090 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
X_11778_ net265 net2583 net594 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13517_ team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__or4b_2
X_16305_ clknet_leaf_23_wb_clk_i _02445_ _01113_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10729_ team_02_WB.instance_to_wrap.top.pc\[31\] _06244_ vssd1 vssd1 vccd1 vccd1
+ _06246_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14497_ net1158 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16236_ clknet_leaf_21_wb_clk_i _02376_ _01044_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13448_ _03038_ _02763_ _03051_ _02768_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11202__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ clknet_leaf_27_wb_clk_i _02307_ _00975_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12472__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ team_02_WB.instance_to_wrap.ramload\[8\] net1010 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[8\] sky130_fd_sc_hd__and2_1
XFILLER_0_109_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10781__A _05579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15118_ net1104 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09347__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16098_ clknet_leaf_123_wb_clk_i _02238_ _00906_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15707__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15049_ net1195 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
X_07940_ _03645_ _03647_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor2_1
XANTENNA__10308__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_wire634_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07871_ _03555_ _03570_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15084__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11816__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ _05123_ _05126_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_121_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15857__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09541_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\] net710 _05056_ _05057_
+ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_30_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09472_ _04982_ _04984_ _04986_ _04988_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_138_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ _04126_ _04129_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12647__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14428__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout247_A _06372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ _04051_ _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09634__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08285_ _03995_ _03996_ _03974_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__or3b_2
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12382__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14163__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout783_A _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10952__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15387__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16632__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1208 net1209 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_2
Xfanout1219 net1220 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_4
Xfanout232 net235 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
XANTENNA__09165__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout243 _06282_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
Xfanout254 _06466_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_2
Xfanout265 net267 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11726__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net279 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout287 _06766_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_2
X_09808_ _05318_ _05320_ _05322_ _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__or4_1
XANTENNA__08912__A2 _04200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout298 net299 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10180__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_104_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09739_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\] net743 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\]
+ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _05123_ _05167_ _05207_ _07273_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10483__A1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11701_ net605 _07184_ _07186_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__and3_2
XANTENNA__12557__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12681_ net269 net1996 net430 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__mux2_1
XANTENNA__13242__A _06490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14420_ net1090 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
X_11632_ net666 net377 _06534_ _07116_ _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_13_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14351_ net1111 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire611 _05270_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_2
X_11563_ _07015_ _07052_ net365 vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire622 net623 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__buf_1
XFILLER_0_68_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13302_ net2169 net984 net965 _03000_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__a22o_1
Xwire633 _05035_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10514_ _05968_ _06030_ _05969_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14282_ net1156 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11494_ _05559_ _05924_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__xnor2_1
X_16021_ clknet_leaf_42_wb_clk_i _02161_ _00829_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13233_ net1055 team_02_WB.instance_to_wrap.top.ru.state\[4\] net1461 vssd1 vssd1
+ vccd1 vccd1 _00011_ sky130_fd_sc_hd__a21o_1
XANTENNA__12292__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10445_ net838 _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13164_ team_02_WB.instance_to_wrap.top.pc\[8\] net1023 _02927_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01489_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10376_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\] net829 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12115_ net250 net2253 net466 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13095_ net229 _02869_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nand2_1
XANTENNA__09156__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12046_ net237 net2227 net470 vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__mux2_1
XANTENNA__11499__B1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16854_ net1398 vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__B1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10710__A2 _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15805_ clknet_leaf_51_wb_clk_i _01945_ _00613_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16785_ net1329 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
X_13997_ net1140 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15736_ clknet_leaf_53_wb_clk_i _01876_ _00544_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12948_ _07467_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10474__A1 _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12467__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ net507 _05671_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__nand2_1
X_15667_ clknet_leaf_54_wb_clk_i _01807_ _00475_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10776__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14618_ net1167 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15598_ clknet_leaf_8_wb_clk_i _01738_ _00406_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14549_ net1214 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10777__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08070_ _03765_ _03787_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__nor2_2
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15079__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16219_ clknet_leaf_127_wb_clk_i _02359_ _01027_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09395__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08972_ _04482_ _04488_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14711__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ _03618_ _03637_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__and2_1
XANTENNA__09147__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold18 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[3\] vssd1 vssd1 vccd1 vccd1
+ net1476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 _02594_ vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07854_ _03304_ net329 _03543_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10162__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10701__A2 _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07785_ _03471_ net364 _03472_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16035__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09524_ _05038_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09855__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09455_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\] net927 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12377__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08406_ _04113_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16185__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09386_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\] net911 net898 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\]
+ _04888_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11414__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ _04046_ _04049_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08268_ _03945_ _03948_ _03957_ _03960_ _03935_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__a41o_1
XANTENNA_fanout998_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08199_ _03910_ _03867_ _03905_ _03913_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10230_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\] net819 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\]
+ _05746_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__a221o_1
XANTENNA__09386__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\] net905 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 net1006 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_4
Xfanout1016 team_02_WB.instance_to_wrap.top.ru.next_iready vssd1 vssd1 vccd1 vccd1
+ net1016 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09138__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1027 _07338_ vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
X_10092_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\] net725 net846 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__a22o_1
Xfanout1038 _04245_ vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1049 net1050 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08346__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10153__A0 _05625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ net1149 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08897__B2 team_02_WB.instance_to_wrap.ramload\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13851_ net1224 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ net998 net552 _07232_ _07235_ _07325_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_35_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13782_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ _03271_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__and3_1
X_16570_ clknet_leaf_92_wb_clk_i _02694_ _01377_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09846__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ _06310_ _06335_ net393 vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09310__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15521_ clknet_leaf_121_wb_clk_i _01661_ _00329_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12733_ _06427_ _06603_ _07256_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__or3_1
XFILLER_0_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12287__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15452_ clknet_leaf_46_wb_clk_i _01592_ _00260_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12664_ _07013_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\] net436 vssd1
+ vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__mux2_1
X_14403_ net1146 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
X_11615_ net669 _07098_ _07099_ net666 _07102_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15383_ clknet_leaf_116_wb_clk_i _01523_ _00191_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12595_ net321 net2549 net438 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14334_ net1191 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
X_11546_ net394 _06960_ _07036_ net381 vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08821__B2 team_02_WB.instance_to_wrap.ramaddr\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13158__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14265_ net1132 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11477_ team_02_WB.instance_to_wrap.top.pc\[9\] _06257_ vssd1 vssd1 vccd1 vccd1 _06972_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_55_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16004_ clknet_leaf_0_wb_clk_i _02144_ _00812_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13216_ net1569 net1021 net938 _05205_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10428_ _05082_ _05944_ _05081_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09377__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14196_ net1091 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13147_ _07480_ _07481_ _07508_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__or3_1
X_10359_ _05869_ _05875_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__nor2_4
XANTENNA__14531__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09129__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ net979 _07429_ _02854_ _02855_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__o31ai_1
XANTENNA__11366__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12029_ net312 net1879 net474 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10144__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16837_ net1381 vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07570_ team_02_WB.instance_to_wrap.top.pad.count\[1\] team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__and2_1
X_16768_ net1312 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_18_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09301__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15719_ clknet_leaf_27_wb_clk_i _01859_ _00527_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12197__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16699_ net1266 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_53_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09240_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\] net834 net903 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\]
+ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09171_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\] net827 net861 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\]
+ _04687_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08122_ _03815_ _03816_ _03801_ _03803_ _03807_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08053_ _03731_ _03768_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12660__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1021_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1119_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08955_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\] net708 net693 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout579_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ _03596_ _03597_ _03624_ _03587_ _03586_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13057__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ net9 net1029 net987 net1653 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__o22a_1
XANTENNA__15425__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07837_ _03525_ _03534_ _03527_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09540__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout746_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ _03442_ _03486_ _03487_ _03440_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__a22o_1
XANTENNA__09828__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09507_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\] net892 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07699_ _03392_ _03421_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout913_A _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09438_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\] net743 _04953_ _04954_
+ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09369_ _04885_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13214__A2_N net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11400_ _06794_ _06897_ net395 vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12380_ net249 net2160 net458 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11331_ net849 _06161_ _06248_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14050_ net1210 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
XANTENNA__09359__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11262_ net946 _06759_ _06765_ net606 vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__o211a_2
XFILLER_0_127_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13001_ _07463_ _07520_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__and2b_1
X_10213_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\] net706 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__a22o_1
XANTENNA__12570__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11193_ _06037_ _06698_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10374__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input42_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\] net729 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a22o_1
XANTENNA__11694__B _07137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13312__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14952_ net1175 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
XANTENNA__10126__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\] net831 net900 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__a22o_1
X_13903_ net1252 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
XANTENNA__11874__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09531__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14883_ net1147 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
XANTENNA__11914__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15182__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16622_ clknet_leaf_97_wb_clk_i _02741_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13834_ net1234 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
X_13765_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _03264_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16553_ clknet_leaf_97_wb_clk_i _02677_ _01360_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_10977_ _06122_ _06482_ _06489_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__a21oi_4
XANTENNA__13091__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15504_ clknet_leaf_41_wb_clk_i _01644_ _00312_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12716_ _06929_ _07239_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16484_ clknet_leaf_67_wb_clk_i net1657 _01292_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
X_13696_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] _03217_ net1658 vssd1 vssd1
+ vccd1 vccd1 _03220_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12647_ net262 net2737 net435 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15435_ clknet_leaf_117_wb_clk_i _01575_ _00243_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15366_ clknet_leaf_59_wb_clk_i _01506_ _00179_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[25\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_87_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12578_ _06498_ net2270 net438 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10773__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11529_ _05649_ _06110_ net661 _05647_ _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__a221o_1
X_14317_ net1132 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
X_15297_ clknet_leaf_76_wb_clk_i _01441_ _00110_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold307 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 team_02_WB.instance_to_wrap.top.a1.row2\[12\] vssd1 vssd1 vccd1 vccd1 net1776
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ net1175 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
Xhold329 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12480__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14179_ net1130 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
XANTENNA__10365__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15448__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 net812 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__buf_6
XFILLER_0_42_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09770__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16769__1313 vssd1 vssd1 vccd1 vccd1 _16769__1313/HI net1313 sky130_fd_sc_hd__conb_1
XANTENNA__13303__B1 _06989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ _04302_ net931 _04358_ _04368_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__and4_1
Xhold1007 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10117__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1029 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08671_ net1056 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] team_02_WB.instance_to_wrap.top.a1.instruction\[26\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 _04300_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_94_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11824__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__or2_2
XANTENNA__15092__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16710__1269 vssd1 vssd1 vccd1 vccd1 _16710__1269/HI net1269 sky130_fd_sc_hd__conb_1
XFILLER_0_117_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07603__A team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11617__A0 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07553_ team_02_WB.instance_to_wrap.top.pc\[12\] vssd1 vssd1 vccd1 vccd1 _03294_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\] net683 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12655__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout327_A _06975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1069_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\] net704 _04662_ _04663_
+ _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09589__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08105_ _03796_ _03821_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__xor2_2
X_09085_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\] net878 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1236_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08036_ _03741_ _03743_ _03751_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_9_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold830 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold841 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout696_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold852 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold863 team_02_WB.instance_to_wrap.top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net2321
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12390__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10356__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold885 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16373__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09761__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09987_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\] net928 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\]
+ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout863_A _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ _04268_ _04346_ _04283_ net1000 vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08869_ net1055 team_02_WB.instance_to_wrap.wb.prev_BUSY_O net1030 vssd1 vssd1 vccd1
+ vccd1 _04431_ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10900_ net838 _06376_ _06414_ net669 _06412_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__o221a_2
XANTENNA__11734__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11880_ net266 net2656 net488 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11608__B1 _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ net398 _06346_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11084__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] net1048 vssd1 vssd1 vccd1
+ vccd1 _03105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10762_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] _04334_ vssd1 vssd1 vccd1
+ vccd1 _06279_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12501_ net343 net2617 net560 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__mux2_1
X_13481_ team_02_WB.START_ADDR_VAL_REG\[21\] net1070 net1003 vssd1 vssd1 vccd1 vccd1
+ net205 sky130_fd_sc_hd__a21o_1
X_10693_ team_02_WB.instance_to_wrap.top.pc\[15\] _06194_ vssd1 vssd1 vccd1 vccd1
+ _06210_ sky130_fd_sc_hd__or2_1
XANTENNA__12565__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15220_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[11\]
+ _00033_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12432_ net333 net2040 net454 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__mux2_1
XANTENNA__11689__B _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15151_ net1247 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
X_12363_ net319 net1805 net563 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14102_ net1096 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
X_11314_ net1699 net301 net641 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
X_15082_ net1252 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12294_ net296 net1755 net570 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14033_ net1118 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
XANTENNA__11909__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11245_ net414 _06513_ _06748_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_120_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14081__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10347__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09752__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ team_02_WB.instance_to_wrap.top.pc\[21\] _06265_ vssd1 vssd1 vccd1 vccd1
+ _06683_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08960__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15740__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\] net835 net896 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\]
+ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a221o_1
X_15984_ clknet_leaf_39_wb_clk_i _02124_ _00792_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11847__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14935_ net1172 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
X_10058_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\] net764 _05560_ _05574_
+ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11311__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14866_ net1123 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15890__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16605_ clknet_leaf_81_wb_clk_i _02724_ _01398_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_13817_ net1224 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__inv_2
X_14797_ net1156 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16893__1437 vssd1 vssd1 vccd1 vccd1 _16893__1437/HI net1437 sky130_fd_sc_hd__conb_1
X_16536_ clknet_leaf_93_wb_clk_i _02663_ _01343_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13748_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] _03251_ net949 vssd1
+ vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_57_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12475__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16467_ clknet_leaf_77_wb_clk_i net1550 _01275_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10784__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13679_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\] _03198_ vssd1 vssd1 vccd1
+ vccd1 _03210_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13160__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13293__A1_N _06883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15418_ clknet_leaf_118_wb_clk_i _01558_ _00226_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16398_ clknet_leaf_65_wb_clk_i _02533_ _01206_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11378__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08779__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15349_ clknet_leaf_86_wb_clk_i _01489_ _00162_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_79_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold104 _02593_ vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 team_02_WB.instance_to_wrap.ramaddr\[31\] vssd1 vssd1 vccd1 vccd1 net1573
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10050__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09991__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold126 team_02_WB.instance_to_wrap.top.a1.row1\[122\] vssd1 vssd1 vccd1 vccd1 net1584
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold137 team_02_WB.START_ADDR_VAL_REG\[31\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11819__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 team_02_WB.instance_to_wrap.top.a1.row2\[0\] vssd1 vssd1 vccd1 vccd1 net1606
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15087__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09910_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\] net768 net740 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold159 team_02_WB.instance_to_wrap.top.a1.row2\[18\] vssd1 vssd1 vccd1 vccd1 net1617
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12878__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10950__C net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout606 net608 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_4
Xfanout617 net619 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_8
X_09841_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\] net926 net922 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a22o_1
XANTENNA__09743__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _05274_ _05284_ _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__nor4_2
X_08723_ net1061 _04266_ _04289_ _04346_ _04269_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_52_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08654_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] team_02_WB.instance_to_wrap.top.a1.instruction\[6\]
+ _04262_ net1062 vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_55_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10678__B _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] _03325_ _03322_ team_02_WB.instance_to_wrap.top.a1.dataIn\[24\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1 vccd1 _03328_
+ sky130_fd_sc_hd__o2111ai_4
X_08585_ net1 _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__nand2_1
XANTENNA__09259__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout444_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13055__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1186_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12385__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout709_A _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09206_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\] net906 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__a22o_1
XANTENNA__15613__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09137_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\] net749 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09068_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\] net727 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\]
+ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__a221o_1
XANTENNA__09982__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout980_A _04177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08019_ _03740_ _03741_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__nor2_1
XANTENNA__11729__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10329__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net383 _06537_ _06538_ _06540_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__a31o_1
Xhold682 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A2 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12981_ _07490_ _07500_ _07489_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_107_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13294__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13245__A _06365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14720_ net1210 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
X_11932_ _07013_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] net484 vssd1
+ vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10588__B _04464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11863_ net333 net1811 net492 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
X_14651_ net1160 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10814_ _05231_ net384 vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nor2_1
X_13602_ team_02_WB.instance_to_wrap.top.a1.row1\[2\] _03119_ _03122_ team_02_WB.instance_to_wrap.top.a1.row2\[10\]
+ _03149_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__a221o_1
X_11794_ net325 net1859 net595 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux2_1
X_14582_ net1096 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16321_ clknet_leaf_121_wb_clk_i _02461_ _01129_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13533_ _03075_ _03077_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__nor2_1
XANTENNA__12295__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10745_ team_02_WB.instance_to_wrap.top.pc\[16\] team_02_WB.instance_to_wrap.top.pc\[15\]
+ _06261_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16768__1312 vssd1 vssd1 vccd1 vccd1 _16768__1312/HI net1312 sky130_fd_sc_hd__conb_1
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13464_ team_02_WB.START_ADDR_VAL_REG\[4\] _04260_ vssd1 vssd1 vccd1 vccd1 net218
+ sky130_fd_sc_hd__and2_1
X_16252_ clknet_leaf_47_wb_clk_i _02392_ _01060_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10280__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ net994 _05740_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ net266 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\] net456 vssd1
+ vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__mux2_1
X_15203_ net1261 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13395_ team_02_WB.instance_to_wrap.ramload\[24\] net1012 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[24\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16183_ clknet_leaf_125_wb_clk_i _02323_ _00991_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15134_ net1230 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
X_12346_ net251 net1775 net564 vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput209 net209 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_0_49_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15065_ net1257 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_116_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12277_ net242 net1978 net572 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14016_ net1210 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09186__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ _06221_ _06222_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16724__1279 vssd1 vssd1 vccd1 vccd1 _16724__1279/HI net1279 sky130_fd_sc_hd__conb_1
X_11159_ _06405_ _06665_ net415 vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15967_ clknet_leaf_86_wb_clk_i _02107_ _00775_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10099__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14918_ net1083 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
XANTENNA__11296__A1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15898_ clknet_leaf_121_wb_clk_i _02038_ _00706_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14849_ net1211 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08370_ _04073_ _04079_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15636__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09110__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16519_ clknet_leaf_5_wb_clk_i _02653_ _01326_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08464__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10023__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__B2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09716__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 net406 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_2
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout425 _03427_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout436 net437 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_6
XANTENNA__11523__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout447 net449 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_8
X_09824_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\] net758 _05340_ vssd1
+ vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1101_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout458 _07220_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_8
Xfanout469 _07211_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12888__B _05536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09755_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\] net895 net939 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout561_A _07219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13276__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16411__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout659_A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ _04308_ _04330_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__or2_1
XANTENNA__11287__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09686_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\] net907 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08637_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04265_ vssd1 vssd1 vccd1
+ vccd1 _04266_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout826_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07998__A team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08568_ team_02_WB.instance_to_wrap.top.a1.row1\[60\] _04235_ _04225_ vssd1 vssd1
+ vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09101__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08499_ team_02_WB.instance_to_wrap.top.a1.data\[9\] net958 _04193_ vssd1 vssd1 vccd1
+ vccd1 _04194_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10530_ _06045_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__nor2_1
XANTENNA__10262__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10461_ net528 _05166_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12200_ net327 net2540 net579 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10014__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ net1026 _02940_ net1025 team_02_WB.instance_to_wrap.top.pc\[5\] vssd1 vssd1
+ vccd1 vccd1 _01486_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09955__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ net415 net609 vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12131_ net319 net2419 net467 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09168__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ net305 net2322 net470 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
Xhold490 team_02_WB.instance_to_wrap.ramload\[7\] vssd1 vssd1 vccd1 vccd1 net1948
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16892__1436 vssd1 vssd1 vccd1 vccd1 _16892__1436/HI net1436 sky130_fd_sc_hd__conb_1
XANTENNA__15509__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ team_02_WB.instance_to_wrap.top.pc\[26\] _06268_ vssd1 vssd1 vccd1 vccd1
+ _06525_ sky130_fd_sc_hd__nor2_1
XANTENNA__11514__A2 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16870_ net1414 vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout970 net972 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_4
X_15821_ clknet_leaf_33_wb_clk_i _01961_ _00629_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13267__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16091__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15752_ clknet_leaf_16_wb_clk_i _01892_ _00560_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12964_ _07482_ _07483_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09340__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
X_14703_ net1115 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
X_11915_ net260 net2489 net483 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ clknet_leaf_125_wb_clk_i _01823_ _00491_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _07377_ _07380_ _07413_ _06205_ _05356_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__a32o_1
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11922__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15190__A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ net1180 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
X_11846_ net265 net2588 net491 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11777_ net259 net2101 net593 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux2_1
X_14565_ net1087 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16304_ clknet_leaf_39_wb_clk_i _02444_ _01112_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10728_ _06244_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__inv_2
X_13516_ team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__or4b_2
XANTENNA__10253__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A_N team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14496_ net1158 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16235_ clknet_leaf_117_wb_clk_i _02375_ _01043_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10659_ net995 _05442_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13447_ _03038_ _02763_ _03051_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11202__A1 _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10005__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16166_ clknet_leaf_43_wb_clk_i _02306_ _00974_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13378_ team_02_WB.instance_to_wrap.ramload\[7\] net1010 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[7\] sky130_fd_sc_hd__and2_1
XANTENNA__11202__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10781__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15117_ net1103 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ net312 net1664 net565 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__mux2_1
X_16097_ clknet_leaf_117_wb_clk_i _02237_ _00905_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09159__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15048_ net1201 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07870_ _03554_ _03570_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09540_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\] net782 net750 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12466__A0 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_84_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09331__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\] net919 net863 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\]
+ _04987_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14709__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08422_ _04121_ _04125_ _04114_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_138_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12769__A1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08353_ _04046_ _04049_ _04058_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_28_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08284_ _03974_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12663__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout407_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16839__1383 vssd1 vssd1 vccd1 vccd1 _16839__1383/HI net1383 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_93_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13194__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1149_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09937__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout776_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1209 net1212 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_4
Xfanout233 net235 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_2
Xfanout244 _06372_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
Xfanout255 _03703_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16767__1311 vssd1 vssd1 vccd1 vccd1 _16767__1311/HI net1311 sky130_fd_sc_hd__conb_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout266 net267 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09570__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09807_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\] net825 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\]
+ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__a221o_1
XANTENNA__15801__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 net279 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout288 net291 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13249__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ _03305_ net255 vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__xnor2_1
Xfanout299 _06865_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_104_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09738_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\] net747 net739 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09322__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09669_ _05180_ _05182_ _05184_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nor4_2
XANTENNA__08381__A_N team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15951__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] _04347_ net953 _07185_ vssd1
+ vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__a211o_1
X_12680_ net260 net2507 net431 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__mux2_1
XANTENNA__10483__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__A1 _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11631_ net671 _07117_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08428__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10235__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ _06290_ _06292_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14350_ net1138 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16723__1278 vssd1 vssd1 vccd1 vccd1 _16723__1278/HI net1278 sky130_fd_sc_hd__conb_1
XFILLER_0_0_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire612 net613 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire623 _05689_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_1
XFILLER_0_110_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire634 net635 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_2
X_10513_ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__inv_2
X_13301_ team_02_WB.instance_to_wrap.top.pc\[9\] net1051 _06970_ net933 vssd1 vssd1
+ vccd1 vccd1 _03000_ sky130_fd_sc_hd__a22o_2
XFILLER_0_134_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14281_ net1109 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
X_11493_ _06985_ _06986_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13232_ net648 net937 net1019 net1538 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a2bb2o_1
X_16020_ clknet_leaf_12_wb_clk_i _02160_ _00828_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input72_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10444_ _04569_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__xor2_1
XANTENNA__13185__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15331__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16457__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13077__A1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ net228 _02926_ _02925_ _02923_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10375_ _05887_ _05888_ _05890_ _05891_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12114_ net252 net1787 net468 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_1
X_16746__1291 vssd1 vssd1 vccd1 vccd1 _16746__1291/HI net1291 sky130_fd_sc_hd__conb_1
XFILLER_0_62_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13094_ _07463_ _07520_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13488__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12045_ net245 net2171 net471 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11499__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09561__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16853_ net1397 vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15804_ clknet_leaf_45_wb_clk_i _01944_ _00612_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12448__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16784_ net1328 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_66_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13996_ net1071 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
XANTENNA__13645__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15735_ clknet_leaf_14_wb_clk_i _01875_ _00543_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12947_ team_02_WB.instance_to_wrap.top.pc\[16\] _06194_ vssd1 vssd1 vccd1 vccd1
+ _07467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15666_ clknet_leaf_3_wb_clk_i _01806_ _00474_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12878_ _05695_ net499 _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_115_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10776__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14617_ net1140 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
X_11829_ net336 net1966 net591 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__mux2_1
X_15597_ clknet_leaf_24_wb_clk_i _01737_ _00405_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10226__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14548_ net1089 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12483__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14479_ net1111 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XANTENNA__10792__A _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07577__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16218_ clknet_leaf_120_wb_clk_i _02358_ _01026_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09919__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16149_ clknet_leaf_41_wb_clk_i _02289_ _00957_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15824__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\] net756 _04483_ _04485_
+ _04487_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__a2111o_2
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13479__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15095__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11827__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07922_ _03639_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold19 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[5\] vssd1 vssd1 vccd1 vccd1
+ net1477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09552__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__A _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ _03304_ _03543_ net329 vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__nand3_1
XANTENNA__15974__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07784_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] _03506_ _03504_ _03503_ vssd1
+ vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09523_ _05016_ _05036_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12658__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13343__A team_02_WB.instance_to_wrap.ramload\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09454_ _04970_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1099_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15204__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11662__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08405_ _04090_ _04112_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__xnor2_1
X_09385_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\] net810 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\]
+ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16891__1435 vssd1 vssd1 vccd1 vccd1 _16891__1435/HI net1435 sky130_fd_sc_hd__conb_1
XFILLER_0_136_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10217__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _04019_ _04038_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_95_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11414__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09083__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15354__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ _03963_ _03982_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08830__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08198_ _03909_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout893_A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12914__A1 _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10160_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\] net884 _04550_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\]
+ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__a221o_1
XANTENNA__09791__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1007 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__buf_2
XFILLER_0_41_1642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1017 team_02_WB.instance_to_wrap.top.ru.next_iready vssd1 vssd1 vccd1 vccd1
+ net1017 sky130_fd_sc_hd__clkbuf_2
X_10091_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\] net785 _05606_ _05607_
+ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a211o_1
Xfanout1028 _07337_ vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_4
Xfanout1039 net1040 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__buf_2
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09543__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08897__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13850_ net1224 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12801_ _07324_ _07323_ _07322_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13781_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\]
+ _03269_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\] vssd1
+ vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__a31o_1
XANTENNA__12568__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ _06328_ _06341_ net409 vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__mux2_1
XANTENNA__11102__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15520_ clknet_leaf_109_wb_clk_i _01660_ _00328_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12732_ _06485_ _07255_ _06647_ _06660_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_35_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15451_ clknet_leaf_127_wb_clk_i _01591_ _00259_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12663_ net334 net2068 net436 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__mux2_1
X_14402_ net1205 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
X_11614_ _05832_ net664 _07100_ net837 _07101_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__o221a_1
XANTENNA__10208__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15382_ clknet_leaf_35_wb_clk_i _01522_ _00190_ vssd1 vssd1 vccd1 vccd1 team_02_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09074__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12594_ net317 net2683 net438 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14333_ net1086 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11545_ net394 _07035_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__nand2_1
XANTENNA__08821__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14264_ net1193 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
XANTENNA__15847__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11476_ net945 _06970_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11169__B1 _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16003_ clknet_leaf_125_wb_clk_i _02143_ _00811_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08513__C _04203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ _05127_ _05943_ _05123_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__o21ba_1
X_13215_ net2756 _00012_ net938 _05164_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14195_ net1167 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09782__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\] net681 _05871_ _05873_
+ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_46_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13146_ team_02_WB.instance_to_wrap.top.pc\[11\] net1023 _02912_ vssd1 vssd1 vccd1
+ vccd1 _01492_ sky130_fd_sc_hd__a21o_1
XANTENNA__15997__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13077_ net230 _02853_ _06653_ net234 vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__o2bb2a_1
X_10289_ _05795_ _05800_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__nor3_2
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09534__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ net307 net1938 net474 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08888__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16836_ net1380 vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_2
XANTENNA__15227__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12986__B _05536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16838__1382 vssd1 vssd1 vccd1 vccd1 _16838__1382/HI net1382 sky130_fd_sc_hd__conb_1
XFILLER_0_88_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12478__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ net1311 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
X_13979_ net1156 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15718_ clknet_leaf_49_wb_clk_i _01858_ _00526_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16698_ net138 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15377__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15649_ clknet_leaf_121_wb_clk_i _01789_ _00457_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\] net917 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a22o_1
XANTENNA__09065__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08121_ _03815_ _03816_ _03801_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16766__1310 vssd1 vssd1 vccd1 vccd1 _16766__1310/HI net1310 sky130_fd_sc_hd__conb_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08812__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ _03718_ _03772_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11130__B net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09773__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10383__A1 _04422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08954_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\] net789 net721 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07905_ net316 _03597_ _03626_ _03587_ _03586_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_138_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08885_ net10 net1032 _04431_ team_02_WB.instance_to_wrap.ramload\[17\] vssd1 vssd1
+ vccd1 vccd1 _02545_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout474_A _07206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16722__1277 vssd1 vssd1 vccd1 vccd1 _16722__1277/HI net1277 sky130_fd_sc_hd__conb_1
X_07836_ _03525_ _03527_ _03535_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_93_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16152__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13085__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ _03474_ _03489_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout641_A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout739_A _04379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09506_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\] net916 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\]
+ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07698_ _03378_ _03387_ _03395_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09437_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\] net751 net703 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__a22o_1
X_16745__1290 vssd1 vssd1 vccd1 vccd1 _16745__1290/HI net1290 sky130_fd_sc_hd__conb_1
XFILLER_0_13_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout906_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ _04878_ _04884_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__nor2_4
XANTENNA__09056__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08319_ _04006_ _04029_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nand2_1
X_09299_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\] net830 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\]
+ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__a221o_1
XANTENNA__08803__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11330_ _06198_ _06209_ _06211_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__nand3_1
XANTENNA__10071__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11261_ net974 _06760_ _06764_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10212_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\] net738 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__a22o_1
X_13000_ _07464_ _07519_ _07465_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09764__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _06432_ _06639_ _06697_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10143_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\] net721 _05652_ _05653_
+ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13248__A _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09516__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13312__B2 _03005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input35_A gpio_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14951_ net1105 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
X_10074_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\] net815 net908 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\]
+ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a221o_1
XANTENNA__11323__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ net1261 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
XANTENNA__10677__A2 _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14882_ net1161 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
X_16621_ clknet_leaf_98_wb_clk_i _02740_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13833_ net1233 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
XANTENNA__12298__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16552_ clknet_leaf_93_wb_clk_i _02676_ _01359_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[111\]
+ sky130_fd_sc_hd__dfstp_1
X_13764_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _03263_ sky130_fd_sc_hd__and3_1
XANTENNA__09295__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08077__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10976_ net673 _06469_ _06485_ net672 _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15503_ clknet_leaf_34_wb_clk_i _01643_ _00311_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12715_ _06969_ _07238_ _06988_ _06949_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__or4b_1
XFILLER_0_6_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16483_ clknet_leaf_67_wb_clk_i net1610 _01291_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
X_13695_ net2134 _03217_ _03219_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14807__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11930__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15434_ clknet_leaf_130_wb_clk_i _01574_ _00242_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12646_ net265 net2500 net435 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15365_ clknet_leaf_83_wb_clk_i _01505_ _00178_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[24\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12577_ net252 net2283 net441 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ net1072 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11528_ _05648_ _06116_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15296_ clknet_leaf_76_wb_clk_i _01440_ _00109_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold308 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16025__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold319 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
X_14247_ net1101 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
X_11459_ net945 _06950_ _06954_ net605 vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__o211a_2
XANTENNA__09755__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ net1207 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13129_ _07375_ _07376_ _07415_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a21oi_1
XANTENNA__16175__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16890__1434 vssd1 vssd1 vccd1 vccd1 _16890__1434/HI net1434 sky130_fd_sc_hd__conb_1
XANTENNA__09507__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13303__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1019 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1
+ net2477 sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] team_02_WB.instance_to_wrap.top.a1.instruction\[29\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] team_02_WB.instance_to_wrap.top.a1.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__and4_1
XFILLER_0_108_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07621_ team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] _03337_ vssd1 vssd1 vccd1
+ vccd1 _03344_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16819_ net1363 vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__buf_2
X_07552_ team_02_WB.instance_to_wrap.top.pc\[30\] vssd1 vssd1 vccd1 vccd1 _03293_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11617__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12001__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09286__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14717__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11840__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09222_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\] net775 _04737_ _04738_
+ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09038__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\] net781 _04666_ _04667_
+ _04669_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_1_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08104_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] _03821_ _03822_ vssd1 vssd1
+ vccd1 vccd1 _03824_ sky130_fd_sc_hd__or3_1
XANTENNA__11141__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__A0 _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09084_ _04595_ _04597_ _04598_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__or4_1
XFILLER_0_114_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08035_ _03743_ _03751_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput80 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
Xhold820 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12671__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1131_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput91 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
Xhold831 team_02_WB.instance_to_wrap.ramaddr\[22\] vssd1 vssd1 vccd1 vccd1 net2289
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09746__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold842 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold886 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_A _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold897 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09986_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\] net827 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a22o_1
X_08937_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04293_ _04334_ vssd1
+ vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and3_1
XANTENNA__10108__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10108__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08868_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _04430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07819_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] _03532_ _03533_ vssd1 vssd1
+ vccd1 vccd1 _03542_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08799_ net1 _04245_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10830_ net390 _06345_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_120_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09277__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10761_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ _04334_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11750__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12500_ net337 net2402 net560 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13480_ team_02_WB.START_ADDR_VAL_REG\[20\] _04260_ vssd1 vssd1 vccd1 vccd1 net204
+ sky130_fd_sc_hd__and2_1
XANTENNA__09029__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10692_ _06201_ _06206_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12431_ net325 net2083 net455 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13230__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10044__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09985__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15150_ net1247 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ net312 net2031 net561 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14101_ net1187 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
X_11313_ net946 _06807_ _06814_ net606 vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__o211a_4
X_16837__1381 vssd1 vssd1 vccd1 vccd1 _16837__1381/HI net1381 sky130_fd_sc_hd__conb_1
X_15081_ net1263 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
XANTENNA__12581__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12293_ net308 net2609 net571 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16198__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09737__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ net411 _06747_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__nor2_1
X_14032_ net1076 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
XANTENNA__09201__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ _06180_ net654 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] net496
+ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\] net929 net811 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__a22o_1
X_15983_ clknet_leaf_38_wb_clk_i _02123_ _00791_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13297__B1 _06931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10057_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\] net780 net776 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__a22o_1
X_14934_ net1093 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ net1118 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
XANTENNA__13049__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13425__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08519__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16604_ clknet_leaf_91_wb_clk_i _02723_ _01397_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_13816_ net1222 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10130__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09268__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14796_ net1072 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16535_ clknet_leaf_93_wb_clk_i _02662_ _01342_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_13747_ _03251_ net950 _03250_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__and3b_1
XFILLER_0_57_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10959_ _06051_ _06060_ net392 vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13441__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16466_ clknet_leaf_89_wb_clk_i net1519 _01274_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_2
X_13678_ _03206_ _03209_ net1241 vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10784__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15417_ clknet_leaf_17_wb_clk_i _01557_ _00225_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12629_ net2303 net328 net555 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__mux2_1
X_16397_ clknet_leaf_65_wb_clk_i _02532_ _01205_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13275__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11232__C1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09976__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15415__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15348_ clknet_leaf_85_wb_clk_i _01488_ _00161_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_83_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09440__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12491__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold105 team_02_WB.START_ADDR_VAL_REG\[16\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ clknet_leaf_72_wb_clk_i _01423_ _00092_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold116 team_02_WB.START_ADDR_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold127 team_02_WB.instance_to_wrap.ramstore\[22\] vssd1 vssd1 vccd1 vccd1 net1585
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold138 team_02_WB.instance_to_wrap.ramstore\[6\] vssd1 vssd1 vccd1 vccd1 net1596
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09728__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 team_02_WB.instance_to_wrap.top.a1.row1\[123\] vssd1 vssd1 vccd1 vccd1 net1607
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15565__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout607 net608 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
X_09840_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__a22o_1
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__buf_8
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09771_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\] net899 net856 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\]
+ _05275_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__a221o_1
XANTENNA__13288__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13213__A2_N net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11835__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] team_02_WB.instance_to_wrap.top.a1.instruction\[6\]
+ _04262_ net1062 vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07604_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] _03325_ team_02_WB.instance_to_wrap.top.a1.dataIn\[24\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1 vccd1 _03327_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10040__A _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08584_ team_02_WB.instance_to_wrap.wb.curr_state\[2\] team_02_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__or2_1
XANTENNA__09259__A2 _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13228__A2_N net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08467__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12666__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1081_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1179_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10274__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09205_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\] net797 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\]
+ _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout604_A _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10026__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09967__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ _04630_ _04651_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\] net702 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08018_ _03696_ _03708_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold650 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout973_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold672 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold694 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09969_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\] net740 _05484_ _05485_
+ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__a211o_1
XANTENNA__13279__B1 _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12980_ _07492_ _07499_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__nand2_1
XANTENNA__09498__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ net334 net2449 net484 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10588__C _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14650_ net1180 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11862_ net328 net2173 net492 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13601_ team_02_WB.instance_to_wrap.top.a1.row1\[10\] _03110_ _03128_ team_02_WB.instance_to_wrap.top.a1.row1\[106\]
+ _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__a221o_1
X_10813_ _06319_ _06327_ net408 vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__mux2_1
X_14581_ net1215 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
XANTENNA__08458__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12576__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11793_ net322 net2544 net595 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16320_ clknet_leaf_106_wb_clk_i _02460_ _01128_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13532_ _03091_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10744_ team_02_WB.instance_to_wrap.top.pc\[14\] _06260_ vssd1 vssd1 vccd1 vccd1
+ _06261_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16251_ clknet_leaf_127_wb_clk_i _02391_ _01059_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13463_ team_02_WB.START_ADDR_VAL_REG\[3\] net1069 net1004 vssd1 vssd1 vccd1 vccd1
+ net217 sky130_fd_sc_hd__a21o_1
XANTENNA__13203__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ net790 _05669_ _06127_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__o22a_4
X_15202_ net1259 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ net258 net2475 net456 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09958__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16182_ clknet_leaf_63_wb_clk_i _02322_ _00990_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13394_ net2761 net1012 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[23\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09422__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15188__A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15133_ net1247 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
X_12345_ net237 net2316 net561 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15064_ net1258 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
X_12276_ _04291_ net647 _07190_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__or3_4
XFILLER_0_65_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14015_ net1189 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11227_ net952 _06731_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11158_ _06544_ _06663_ net397 vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10109_ _05580_ _05625_ net551 vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__mux2_1
X_15966_ clknet_leaf_117_wb_clk_i _02106_ _00774_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11089_ _06597_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__inv_2
XANTENNA__09489__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14917_ net1128 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15897_ clknet_leaf_18_wb_clk_i _02037_ _00705_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16213__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14848_ net1158 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08449__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12486__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14779_ net1157 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13171__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ clknet_leaf_37_wb_clk_i _02652_ _01325_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10256__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16363__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09661__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16449_ clknet_leaf_63_wb_clk_i net1586 _01257_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09413__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15098__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11220__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07609__A team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_2
Xfanout415 _05762_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08924__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout437 _07228_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_4
X_09823_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\] net762 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\]
+ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a221o_1
XANTENNA__08924__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_6
Xfanout459 _07220_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_A _05901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ net610 vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08705_ _04308_ _04329_ net650 vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__or3_2
X_09685_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\] net802 net863 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\]
+ _05189_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout554_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ team_02_WB.instance_to_wrap.top.a1.instruction\[2\] team_02_WB.instance_to_wrap.top.a1.instruction\[3\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[0\] team_02_WB.instance_to_wrap.top.a1.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__or4bb_2
X_16836__1380 vssd1 vssd1 vccd1 vccd1 _16836__1380/HI net1380 sky130_fd_sc_hd__conb_1
XFILLER_0_136_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12236__A1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout721_A _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12396__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ _04180_ _04234_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout819_A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10247__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13081__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11995__A0 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08498_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[9\] net980 vssd1 vssd1 vccd1
+ vccd1 _04193_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09652__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08860__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10460_ _05975_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_115_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09404__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09119_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\] net866 vssd1 vssd1
+ vccd1 vccd1 _04636_ sky130_fd_sc_hd__and2_1
X_10391_ net412 net609 vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12130_ net313 net1818 net466 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12061_ net298 net2234 net471 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold480 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11012_ _06148_ _06234_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_70_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout960 _03261_ vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08391__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15820_ clknet_leaf_20_wb_clk_i _01960_ _00628_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout971 net972 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_2
Xfanout982 _03320_ vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 _04427_ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15751_ clknet_leaf_27_wb_clk_i _01891_ _00559_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12963_ team_02_WB.instance_to_wrap.top.pc\[8\] _05583_ vssd1 vssd1 vccd1 vccd1 _07483_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1180 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1191 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
X_14702_ net1096 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
X_11914_ net264 net1868 net483 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ clknet_leaf_124_wb_clk_i _01822_ _00490_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_68_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _07380_ _07413_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_83_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09891__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12227__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14633_ net1112 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11845_ net257 net1856 net490 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14564_ net1130 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
X_11776_ net248 net2071 net593 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09643__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16303_ clknet_leaf_34_wb_clk_i _02443_ _01111_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13515_ _03072_ _03075_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10727_ _06168_ _06243_ _06167_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__a21o_2
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14495_ net1170 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
XANTENNA__08851__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16234_ clknet_leaf_129_wb_clk_i _02374_ _01042_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13446_ _03036_ _03048_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10658_ team_02_WB.instance_to_wrap.top.pc\[23\] _04494_ vssd1 vssd1 vccd1 vccd1
+ _06175_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16165_ clknet_leaf_32_wb_clk_i _02305_ _00973_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11570__A2_N net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ net1771 net1010 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[6\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_11_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10589_ net546 net390 net405 vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__or3_1
X_15116_ net1108 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
X_12328_ net306 net1857 net565 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16096_ clknet_leaf_106_wb_clk_i _02236_ _00904_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_15047_ net1220 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12259_ net300 net2378 net574 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08906__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15949_ clknet_leaf_32_wb_clk_i _02089_ _00757_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09470_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\] net907 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09882__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08421_ _04117_ _04126_ _04123_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_138_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15753__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10229__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12769__A2 _07177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08352_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04059_ _04061_ _04062_ vssd1
+ vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__o211a_1
XANTENNA__09095__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09634__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08842__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08283_ _03952_ _03994_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11729__A0 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1044_A _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10952__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1211_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout234 net235 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
Xfanout245 _06372_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout769_A _04372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 _06530_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_2
Xfanout267 _06564_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
X_09806_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\] net910 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_2
X_07998_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] net255 vssd1 vssd1 vccd1 vccd1
+ _03721_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10180__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout289 net291 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_104_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\] net787 net783 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout936_A _02955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09668_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\] net767 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\]
+ _05169_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09873__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08619_ net76 net1530 net955 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__mux2_1
X_09599_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\] net815 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11630_ _05995_ _05996_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09086__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11561_ net1961 net341 net644 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire613 _05230_ vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ team_02_WB.instance_to_wrap.ramaddr\[10\] net983 net964 _02999_ vssd1 vssd1
+ vccd1 vccd1 _01429_ sky130_fd_sc_hd__a22o_1
Xwire624 _05463_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_2
X_10512_ _04783_ _06028_ net538 _04776_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14280_ net1178 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
Xwire635 _04860_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11492_ net416 net666 _06569_ _06583_ _06983_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__o32a_1
XFILLER_0_134_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13231_ net1666 net1020 _02954_ _05855_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a22o_1
XANTENNA__13185__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10443_ _04611_ _05959_ _04609_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_116_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11196__B2 _06105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input65_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ _07484_ _07504_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_72_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10374_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\] net918 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\]
+ _05886_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10943__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12113_ net238 net1930 net466 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__mux2_1
XANTENNA__12145__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ _07424_ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12044_ net242 net1865 net472 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__mux2_1
XANTENNA__11499__A2 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16852_ net1396 vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_2
XFILLER_0_40_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10171__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout790 net791 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15803_ clknet_leaf_1_wb_clk_i _01943_ _00611_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_16783_ net1327 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13995_ net1150 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11933__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15734_ clknet_leaf_52_wb_clk_i _01874_ _00542_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12999__A2 _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ team_02_WB.instance_to_wrap.top.pc\[17\] _06192_ vssd1 vssd1 vccd1 vccd1
+ _07466_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15665_ clknet_leaf_50_wb_clk_i _01805_ _00473_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12877_ _07388_ _07395_ _07396_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08527__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14616_ net1193 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09077__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ net327 net1905 net591 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15596_ clknet_leaf_15_wb_clk_i _01736_ _00404_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09616__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14547_ net1169 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
X_11759_ net319 net2296 net599 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__mux2_1
XANTENNA__08824__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14478_ net1163 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
XANTENNA__10792__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16217_ clknet_leaf_18_wb_clk_i _02357_ _01025_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13429_ net1066 _03037_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__nand2_2
XANTENNA__16401__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap1063 net1064 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12384__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16148_ clknet_leaf_11_wb_clk_i _02288_ _00956_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16079_ clknet_leaf_38_wb_clk_i _02219_ _00887_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08970_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\] net741 net685 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\]
+ _04486_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_100_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07921_ _03605_ _03638_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07852_ _03304_ net329 vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12004__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__B _04608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10313__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10162__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
X_07783_ _03303_ net364 vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11843__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09522_ _05016_ _05037_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09855__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13343__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _04962_ _04969_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__nor2_8
XFILLER_0_133_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08404_ _04111_ _04107_ _04099_ _04092_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09068__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09384_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\] net830 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07618__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08335_ _04020_ _04038_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__or2_2
XANTENNA__12674__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08815__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1161_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1259_A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08266_ _03958_ _03960_ _03938_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16081__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08197_ _03910_ _03912_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__or2_1
XANTENNA__11178__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15649__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09240__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout886_A _04536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\] net709 net705 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1007 _03315_ vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1018 net1019 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__buf_2
XFILLER_0_41_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1029 net1030 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_2
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15799__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11350__B2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11753__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ _04355_ _07123_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13780_ net1705 _03271_ _03273_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10992_ _06502_ _06503_ net413 vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09846__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12731_ _06501_ _07254_ _06704_ _06730_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__or4b_1
XFILLER_0_74_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16859__1403 vssd1 vssd1 vccd1 vccd1 _16859__1403/HI net1403 sky130_fd_sc_hd__conb_1
XFILLER_0_13_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15450_ clknet_leaf_120_wb_clk_i _01590_ _00258_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09059__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12662_ net327 net2643 net436 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14401_ net1211 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11613_ _05831_ net660 _06113_ _05829_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_33_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08806__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15381_ clknet_leaf_83_wb_clk_i _01521_ _00189_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12584__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16424__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12593_ net313 net2179 net438 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ net1145 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
X_11544_ net388 _07033_ _07034_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ net1173 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09178__B _04694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11475_ net671 _06957_ _06969_ net673 _06968_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__a221o_1
X_16002_ clknet_leaf_123_wb_clk_i _02142_ _00810_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13214_ net630 net937 net1018 net1671 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__a2bb2o_1
Xwire498 _05828_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_2
XFILLER_0_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10426_ _05167_ _05942_ _05168_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__o21ai_1
X_14194_ net1123 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09231__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15196__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11928__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _02908_ _02911_ net1026 vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a21oi_1
X_10357_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\] net789 net745 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16815__1359 vssd1 vssd1 vccd1 vccd1 _16815__1359/HI net1359 sky130_fd_sc_hd__conb_1
XFILLER_0_57_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13076_ _07363_ _07364_ _07428_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10288_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\] net803 _05802_ _05803_
+ _05804_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_40_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12027_ net299 net2480 net476 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10144__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16835_ net1379 vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ net1182 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
X_16766_ net1310 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_73_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09837__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15717_ clknet_leaf_35_wb_clk_i _01857_ _00525_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12929_ team_02_WB.instance_to_wrap.top.pc\[28\] _06143_ vssd1 vssd1 vccd1 vccd1
+ _07449_ sky130_fd_sc_hd__nor2_1
X_16697_ net138 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_17_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15648_ clknet_leaf_118_wb_clk_i _01788_ _00456_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15579_ clknet_leaf_125_wb_clk_i _01719_ _00387_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12494__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08120_ _03838_ _03839_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__and2_1
XANTENNA__09369__A _04885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09470__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08704__C _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08051_ _03744_ _03750_ _03718_ _03732_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__a211o_1
XANTENNA__11411__B net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12357__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09773__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15941__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10383__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07617__A team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _04462_ _04463_ _04467_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__or3_4
XFILLER_0_122_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07904_ _03571_ _03600_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08884_ net11 net1032 _04431_ team_02_WB.instance_to_wrap.ramload\[18\] vssd1 vssd1
+ vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
XANTENNA__10135__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11332__A1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1007_A _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07835_ _03546_ _03550_ _03557_ _03523_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12669__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10978__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07766_ _03465_ _03488_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__and2_1
XANTENNA__09289__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09828__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\] net900 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07697_ _03403_ _03409_ _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10843__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\] net719 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout801_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\] net714 _04880_ _04882_
+ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_75_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08318_ _04000_ _04002_ _04018_ _04006_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__a31o_1
XANTENNA__15471__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09298_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\] net915 _04804_ _04805_
+ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__a211o_1
XANTENNA__09461__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08249_ _03910_ _03925_ _03953_ _03960_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__and4b_1
XFILLER_0_132_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13545__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11260_ _06188_ net654 _06763_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__a21o_1
XANTENNA__09213__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11748__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\] net762 _05717_ _05720_
+ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_63_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11191_ net373 _06437_ _06441_ net378 vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__o22a_1
XANTENNA__10374__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10142_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\] net705 _05655_ _05656_
+ _05658_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13248__B _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput190 net190 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_101_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13312__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14950_ net1073 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
X_10073_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\] net904 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__a22o_1
XANTENNA__10126__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ net1252 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881_ net1160 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
XANTENNA__12579__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13832_ net1232 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
X_16620_ clknet_leaf_98_wb_clk_i _02739_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16551_ clknet_leaf_92_wb_clk_i _02675_ _01358_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ _03064_ net961 _03262_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10975_ net668 _06477_ _06487_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__o21ai_1
X_12714_ _07025_ _07237_ _07057_ _06996_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__or4bb_1
X_15502_ clknet_leaf_10_wb_clk_i _01642_ _00310_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16482_ clknet_leaf_77_wb_clk_i net1547 _01290_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] _03217_ net1242 vssd1 vssd1
+ vccd1 vccd1 _03219_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15814__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15433_ clknet_leaf_105_wb_clk_i _01573_ _00241_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12645_ net256 net1734 net435 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15364_ clknet_leaf_82_wb_clk_i _01504_ _00177_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_12576_ net239 net2015 net438 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14315_ net1202 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
X_11527_ net417 _06636_ _06849_ net375 _07018_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15964__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15295_ clknet_leaf_89_wb_clk_i _01439_ _00108_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13536__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14246_ net1082 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold309 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09204__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11458_ team_02_WB.instance_to_wrap.top.pc\[10\] net973 _06837_ _06953_ vssd1 vssd1
+ vccd1 vccd1 _06954_ sky130_fd_sc_hd__a211o_1
XFILLER_0_106_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10409_ _05513_ _05925_ _05514_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14177_ net1214 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11389_ net998 _06887_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__nor2_1
XANTENNA__10365__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13128_ _07475_ _07512_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__13303__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13059_ _07454_ _07530_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__xnor2_1
Xhold1009 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10117__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12489__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15344__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11393__S net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ _03339_ _03342_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16818_ net1362 vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07551_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1
+ _03292_ sky130_fd_sc_hd__inv_2
X_16749_ net1293 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_18_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15494__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09221_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\] net763 net723 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12578__A0 _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\] net716 _04668_ vssd1
+ vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09443__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ _03821_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__or2_1
XANTENNA__11141__B _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\] net923 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\]
+ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14733__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08034_ _03744_ _03750_ _03733_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_13_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput70 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold810 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xinput81 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
Xhold821 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold832 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput92 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
Xhold843 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08549__A2 _04203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold854 team_02_WB.instance_to_wrap.top.a1.row2\[27\] vssd1 vssd1 vccd1 vccd1 net2312
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10356__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold887 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
X_16858__1402 vssd1 vssd1 vccd1 vccd1 _16858__1402/HI net1402 sky130_fd_sc_hd__conb_1
Xhold898 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09985_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\] net823 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\]
+ _05501_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout584_A _07209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04334_ vssd1 vssd1
+ vccd1 vccd1 _04453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08867_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _04429_ sky130_fd_sc_hd__and2_1
XANTENNA__12399__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout751_A _04376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _03532_ _03533_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1
+ vccd1 vccd1 _03541_ sky130_fd_sc_hd__a21oi_2
X_08798_ team_02_WB.instance_to_wrap.top.testpc.en_latched _04426_ vssd1 vssd1 vccd1
+ vccd1 _02627_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15837__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07749_ _03432_ _03468_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10760_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ _04334_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09682__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16814__1358 vssd1 vssd1 vccd1 vccd1 _16814__1358/HI net1358 sky130_fd_sc_hd__conb_1
X_09419_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\] net871 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a22o_1
XANTENNA__10292__A1 _05807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10691_ _06198_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12430_ net322 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\] net455 vssd1
+ vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13230__B2 _05807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ net306 net2546 net561 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15217__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100_ net1089 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11312_ _06192_ net654 _06809_ _06813_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15080_ net1252 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12292_ net300 net2195 net570 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14031_ net1113 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
X_11243_ _06630_ _06746_ net400 vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10347__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11174_ _06227_ _06680_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08960__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\] net831 net804 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\]
+ _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a221o_1
XANTENNA__16612__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15982_ clknet_leaf_10_wb_clk_i _02122_ _00790_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13297__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14933_ net1185 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
X_10056_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\] net728 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_19_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12102__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10411__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14864_ net1110 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
X_16603_ clknet_leaf_91_wb_clk_i _02722_ _01396_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13815_ net1217 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__inv_2
X_14795_ net1205 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
XANTENNA__10130__B _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13746_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\] _03019_ _03245_ vssd1
+ vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__and3_1
X_16534_ clknet_leaf_93_wb_clk_i _02661_ _01341_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_10958_ _06470_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09673__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16465_ clknet_leaf_78_wb_clk_i net1629 _01273_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13677_ _03198_ _03208_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10889_ net408 _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15416_ clknet_leaf_52_wb_clk_i _01556_ _00224_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12628_ net2486 net321 net554 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__mux2_1
X_16396_ clknet_leaf_65_wb_clk_i _02531_ _01204_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09425__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15347_ clknet_leaf_56_wb_clk_i _01487_ _00160_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08779__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12559_ net306 net1837 net442 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15278_ clknet_leaf_78_wb_clk_i _01422_ _00091_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 team_02_WB.START_ADDR_VAL_REG\[26\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 team_02_WB.instance_to_wrap.ramstore\[11\] vssd1 vssd1 vccd1 vccd1 net1575
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 _02584_ vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold139 _02568_ vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ net1216 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_78_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10292__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout608 _06281_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_2
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout619 net620 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16292__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\] net891 _05272_ _05286_
+ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__a211o_1
XANTENNA__13288__A1 team_02_WB.instance_to_wrap.ramaddr\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ _04287_ _04337_ _04342_ _04323_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1190 net1197 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08652_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] net1000 vssd1 vssd1 vccd1
+ vccd1 _04281_ sky130_fd_sc_hd__or2_2
XANTENNA__12012__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07603_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] _03325_ vssd1 vssd1 vccd1
+ vccd1 _03326_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08583_ team_02_WB.instance_to_wrap.wb.curr_state\[2\] team_02_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__nor2_4
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10040__B _05556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11851__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13460__A1 team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13351__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_A _07013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1074_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09204_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\] net922 net918 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__a22o_1
XANTENNA__09416__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09135_ net968 _04650_ _04497_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__a21o_1
XANTENNA__12682__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1241_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09066_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\] net719 net707 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\]
+ _04582_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08017_ _03675_ _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout799_A _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold640 team_02_WB.instance_to_wrap.ramload\[14\] vssd1 vssd1 vccd1 vccd1 net2098
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10329__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold651 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold673 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09195__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold684 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A _02957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09968_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\] net784 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a22o_1
XANTENNA__10930__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13279__B2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ net1489 _04441_ net930 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09899_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\] net902 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ net327 net2662 net484 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11861_ net323 net2396 net492 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XANTENNA__16015__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11761__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ team_02_WB.instance_to_wrap.top.a1.row1\[18\] _03111_ _03116_ team_02_WB.instance_to_wrap.top.a1.row1\[122\]
+ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10812_ _06327_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14580_ net1092 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
XANTENNA__09655__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ net320 net2398 net593 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13531_ _03085_ _03090_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ team_02_WB.instance_to_wrap.top.pc\[13\] team_02_WB.instance_to_wrap.top.pc\[12\]
+ _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ clknet_leaf_119_wb_clk_i _02390_ _01058_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16165__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13462_ team_02_WB.START_ADDR_VAL_REG\[2\] net1069 net1004 vssd1 vssd1 vccd1 vccd1
+ net214 sky130_fd_sc_hd__a21o_1
XANTENNA__09407__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input95_A wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ net994 _05693_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13203__B2 _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ net1261 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12413_ net248 net2651 net454 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__mux2_1
X_16181_ clknet_leaf_43_wb_clk_i _02321_ _00989_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13393_ team_02_WB.instance_to_wrap.ramload\[22\] net1012 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[22\] sky130_fd_sc_hd__and2_1
XFILLER_0_10_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12592__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15132_ net1248 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
X_12344_ net245 net2722 net562 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15063_ net1248 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
X_12275_ net344 net1971 net573 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14014_ net1191 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
X_11226_ net838 _06713_ _06730_ net670 _06729_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__o221a_2
XANTENNA__09186__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11936__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07645__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11157_ _06663_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10108_ team_02_WB.instance_to_wrap.top.a1.instruction\[26\] _04330_ net650 team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__a22o_1
X_15965_ clknet_leaf_48_wb_clk_i _02105_ _00773_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11088_ _05212_ _05980_ _06017_ _06020_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__o31a_1
X_14916_ net1126 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
X_10039_ _05537_ _05555_ net968 vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__mux2_2
XANTENNA__09894__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15896_ clknet_leaf_19_wb_clk_i _02036_ _00704_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14847_ net1170 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_125_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14778_ net1167 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09646__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16517_ clknet_leaf_35_wb_clk_i _02651_ _01324_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13729_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ _03017_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__and3_1
X_16857__1401 vssd1 vssd1 vccd1 vccd1 _16857__1401/HI net1401 sky130_fd_sc_hd__conb_1
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_128_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16448_ clknet_leaf_46_wb_clk_i net1524 _01256_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16379_ clknet_leaf_93_wb_clk_i net1492 _01187_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12007__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15682__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout405 net406 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_2
Xfanout416 net419 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11846__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09822_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\] net714 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_54_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16813__1357 vssd1 vssd1 vccd1 vccd1 _16813__1357/HI net1357 sky130_fd_sc_hd__conb_1
XANTENNA__08924__A2 _04215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout438 net441 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__clkbuf_8
Xfanout449 _07224_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09753_ _05259_ _05264_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__nor3_1
XFILLER_0_96_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16038__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08704_ _04329_ net652 _04309_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__and3b_2
XANTENNA__13130__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09684_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\] net883 _05188_ _05200_
+ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__a211o_1
XANTENNA__09885__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08635_ net1062 net1060 team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04262_
+ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_136_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12677__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout547_A _04489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16188__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08566_ _02814_ _04228_ _04226_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09637__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09101__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08497_ _04171_ _04185_ _04191_ _04192_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout714_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09118_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\] net817 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\]
+ _04634_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10390_ net412 net609 vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09049_ net547 _04565_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09168__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ net310 net2542 net473 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_1
Xhold470 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08376__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net383 _06104_ _06513_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__a31o_2
XFILLER_0_40_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10183__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout950 _03233_ vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_1
Xfanout961 _03261_ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout972 _04495_ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout983 _02956_ vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net995 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13121__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11057__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ clknet_leaf_42_wb_clk_i _01890_ _00558_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12962_ team_02_WB.instance_to_wrap.top.pc\[8\] _05583_ vssd1 vssd1 vccd1 vccd1 _07482_
+ sky130_fd_sc_hd__and2_1
Xhold1170 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15405__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09876__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09340__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11913_ net259 net2085 net483 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1181 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10486__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14701_ net1141 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1192 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12587__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15681_ clknet_leaf_124_wb_clk_i _01821_ _00489_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12893_ _07379_ _07412_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_83_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ net1177 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
X_11844_ net248 net2470 net490 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ net1145 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15555__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11775_ net253 net2710 net595 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16302_ clknet_leaf_27_wb_clk_i _02442_ _01110_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13514_ team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__or4b_2
X_10726_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] _04283_ _06169_ vssd1
+ vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14494_ net1191 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13188__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15199__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16233_ clknet_leaf_105_wb_clk_i _02373_ _01041_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13445_ _03033_ _02766_ _03049_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10657_ team_02_WB.instance_to_wrap.top.pc\[23\] _04491_ _04493_ vssd1 vssd1 vccd1
+ vccd1 _06174_ sky130_fd_sc_hd__and3_1
XANTENNA__13212__A2_N net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09197__A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13376_ team_02_WB.instance_to_wrap.ramload\[5\] net1010 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[5\] sky130_fd_sc_hd__and2_1
XFILLER_0_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16164_ clknet_leaf_3_wb_clk_i _02304_ _00972_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09800__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10588_ _04458_ _04464_ _04467_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__nand3_1
XFILLER_0_84_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12327_ net299 net2735 net566 vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__mux2_1
X_15115_ net1098 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16095_ clknet_leaf_109_wb_clk_i _02235_ _00903_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15046_ net1219 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
XANTENNA__09159__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12258_ net293 net2094 net574 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__mux2_1
X_11209_ _06091_ _06095_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__or2_1
X_12189_ net288 net2382 net577 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ clknet_leaf_20_wb_clk_i _02088_ _00756_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09867__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15879_ clknet_leaf_26_wb_clk_i _02019_ _00687_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ _04117_ _04126_ _04123_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13182__A _07388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09619__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08351_ _04061_ _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13910__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08282_ _03995_ _03996_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_15_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_93_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09398__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_93_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10952__A2 _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13357__A team_02_WB.instance_to_wrap.ramload\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10165__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_2
Xfanout246 _06372_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_2
XANTENNA__10704__A2 _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 _06530_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_1
XANTENNA__09570__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\] net813 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\]
+ _05321_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a221o_1
Xfanout268 net271 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_2
X_07997_ _03716_ _03717_ _03713_ _03714_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__o211ai_1
Xfanout279 _06686_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout664_A _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\] net723 net719 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__a22o_1
XANTENNA__09322__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09667_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\] net739 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\]
+ _05183_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__a221o_1
XANTENNA__11665__B1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout831_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15578__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_A _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ net77 net1537 net956 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12200__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _05109_ _05110_ _05112_ _05114_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__or4_1
XFILLER_0_96_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08549_ _04202_ _04203_ net653 net793 net1536 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11560_ net947 _07046_ _07050_ net607 vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__o211a_2
XFILLER_0_64_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire614 _04927_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_4
X_10511_ _05970_ _06027_ _05971_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire625 _05418_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ _05559_ net664 _06113_ _05557_ _06984_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__o221a_1
XANTENNA__11645__A2_N net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13230_ net1720 net1022 net938 _05807_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10442_ _05956_ _05958_ _04653_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11196__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _07407_ _07408_ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__a21oi_1
X_10373_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\] net902 net805 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\]
+ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_72_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12112_ net245 net2427 net468 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10943__A2 _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _07366_ _07367_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__nand2b_1
XANTENNA_input58_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12043_ _04452_ _07207_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__nand2_4
XFILLER_0_44_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10156__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16856__1400 vssd1 vssd1 vccd1 vccd1 _16856__1400/HI net1400 sky130_fd_sc_hd__conb_1
XANTENNA__16353__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16851_ net1395 vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_2
XANTENNA__09561__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout780 _04367_ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout791 _04327_ vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_85_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15802_ clknet_leaf_120_wb_clk_i _01942_ _00610_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16782_ net1326 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XANTENNA__09849__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13994_ net1142 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
XANTENNA__09313__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ clknet_leaf_41_wb_clk_i _01873_ _00541_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11656__B1 _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ team_02_WB.instance_to_wrap.top.pc\[18\] _06190_ vssd1 vssd1 vccd1 vccd1
+ _07465_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15664_ clknet_leaf_39_wb_clk_i _01804_ _00472_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12876_ _05695_ net499 vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14615_ net1174 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
X_11827_ net321 net2495 net591 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
X_15595_ clknet_leaf_115_wb_clk_i _01735_ _00403_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14546_ net1120 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
X_11758_ net315 net2278 net597 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__mux2_1
X_16812__1356 vssd1 vssd1 vccd1 vccd1 _16812__1356/HI net1356 sky130_fd_sc_hd__conb_1
XANTENNA__08824__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10709_ _06224_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11689_ _05996_ _07129_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__nand2_1
X_14477_ net1133 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16216_ clknet_leaf_54_wb_clk_i _02356_ _01024_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13428_ team_02_WB.instance_to_wrap.top.lcd.currentState\[4\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ net962 vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap1064 _03310_ vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13359_ team_02_WB.instance_to_wrap.ramload\[21\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[21\] sky130_fd_sc_hd__and2_1
X_16147_ clknet_leaf_53_wb_clk_i _02287_ _00955_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14561__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16078_ clknet_leaf_26_wb_clk_i _02218_ _00886_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07920_ _03602_ _03639_ _03641_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_36_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15029_ net1221 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XANTENNA__10147__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07851_ _03548_ _03573_ _03572_ _03550_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__09552__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10313__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15720__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13905__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_07782_ _03503_ _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09521_ _05016_ _05036_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__or2_1
XANTENNA__09390__A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11647__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09452_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\] net707 _04963_ _04966_
+ _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__a2111o_2
XANTENNA__12020__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08403_ net1725 net1005 net981 _04111_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a22o_1
XANTENNA__15870__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09383_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\] net825 _04887_ _04899_
+ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout245_A _06372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08334_ _03993_ _04045_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08815__B2 team_02_WB.instance_to_wrap.ramaddr\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ _03306_ _03974_ _03977_ _03966_ _03971_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__a311o_1
XFILLER_0_117_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1154_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13291__A1_N _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08196_ _03910_ _03912_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12690__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09565__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout781_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10138__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 _03314_ vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
Xfanout1019 _00012_ vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_1
XFILLER_0_41_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09543__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09719_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\] net877 vssd1 vssd1
+ vccd1 vccd1 _05236_ sky130_fd_sc_hd__and2_1
XANTENNA__11638__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ _06294_ _06303_ net396 vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12730_ _06555_ _07253_ _06742_ _06768_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_70_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12661_ net323 net2366 net436 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08066__A2_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11612_ _05832_ _05905_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__xnor2_1
X_14400_ net1152 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15380_ clknet_leaf_78_wb_clk_i _01520_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12592_ net307 net2023 net438 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ net388 _06997_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__nand2_1
X_14331_ net1159 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14262_ net1094 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11474_ _05925_ _06956_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16001_ clknet_leaf_124_wb_clk_i _02141_ _00809_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13213_ net631 net937 net1018 net1645 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_33_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10425_ _05207_ _05941_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__or2_1
Xwire499 net503 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14193_ net1105 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
XANTENNA__10377__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13144_ _06259_ _06932_ net232 _02910_ net977 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__o32a_1
X_10356_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\] net769 net713 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\]
+ _05872_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__a221o_1
XANTENNA__09782__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13315__B1 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_13075_ _07526_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12105__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10287_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\] net916 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__a22o_1
X_12026_ net309 net2586 net476 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
XANTENNA__09534__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11944__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16834_ net1378 vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15893__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16765_ net1309 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
X_13977_ net1132 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15716_ clknet_leaf_3_wb_clk_i _01856_ _00524_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12928_ _07446_ _07447_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__nand2_1
X_16696_ net138 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10301__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15647_ clknet_leaf_111_wb_clk_i _01787_ _00455_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16249__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12859_ net518 _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15578_ clknet_leaf_119_wb_clk_i _01718_ _00386_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10604__A1 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14529_ net1160 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15273__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ _03744_ _03750_ _03732_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10080__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10368__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09773__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07784__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13306__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07617__B team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ _04462_ _04468_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07903_ _03593_ _03625_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__nand2_2
XFILLER_0_138_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08883_ net12 net1032 _04431_ team_02_WB.instance_to_wrap.ramload\[19\] vssd1 vssd1
+ vccd1 vccd1 _02547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11854__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ _03520_ _03537_ _03554_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__nand3_1
XFILLER_0_100_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08729__A team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__B _06490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07765_ _03441_ _03486_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13354__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09504_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\] net928 net807 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\]
+ _05018_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07696_ _03414_ _03416_ _03418_ _03413_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_56_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10843__A1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09435_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\] net710 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__a22o_1
XANTENNA__12685__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\] net690 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08317_ _04020_ _04021_ _04025_ _04026_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09297_ _04809_ _04810_ _04812_ _04813_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__or4_2
XANTENNA_40 _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09994__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10071__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _03930_ _03959_ _03963_ _03940_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15766__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ _03862_ _03889_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nor2_2
XFILLER_0_63_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10210_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\] net726 _05721_ _05723_
+ _05726_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09764__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11190_ net423 _06694_ _06695_ _06358_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11571__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\] net845 net681 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\]
+ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xoutput191 net191 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XANTENNA__09516__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\] net827 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\]
+ _05588_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a221o_1
X_16811__1355 vssd1 vssd1 vccd1 vccd1 _16811__1355/HI net1355 sky130_fd_sc_hd__conb_1
XANTENNA__11764__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ net1252 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
X_14880_ net1161 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13831_ net1234 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16550_ clknet_leaf_92_wb_clk_i _02674_ _01357_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_13762_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] net2694
+ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10974_ _04734_ _06116_ _06467_ net665 _06486_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15501_ clknet_leaf_23_wb_clk_i _01641_ _00309_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08077__C _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12713_ net673 _07032_ _07079_ _07236_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__nand4_1
XFILLER_0_116_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16481_ clknet_leaf_76_wb_clk_i net1789 _01289_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12595__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13693_ _03217_ _03218_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15296__CLK clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15432_ clknet_leaf_20_wb_clk_i _01572_ _00240_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12644_ net248 net2631 net434 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12575_ net244 net2089 net439 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__mux2_1
X_15363_ clknet_leaf_82_wb_clk_i _01503_ _00176_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14314_ net1167 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11526_ net393 _06939_ _07017_ net381 vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__o211a_1
X_15294_ clknet_leaf_75_wb_clk_i _01438_ _00107_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11939__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13121__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14245_ net1093 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
X_11457_ net998 _06952_ _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1
+ vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10408_ _05558_ _05924_ _05557_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11011__A1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09755__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14176_ net1154 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11388_ _06260_ _06886_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__or2_1
XANTENNA__08963__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10339_ _05836_ _05855_ net968 vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__mux2_1
X_13127_ team_02_WB.instance_to_wrap.top.pc\[14\] net1024 _02896_ _07337_ vssd1 vssd1
+ vccd1 vccd1 _01495_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13058_ _07433_ _02838_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09507__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ net647 _07205_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__nand2_8
XFILLER_0_108_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16817_ net1361 vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__buf_2
XANTENNA__13067__A2 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16071__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07550_ net1861 vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_92_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16748_ net1292 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15639__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09140__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16679_ clknet_leaf_73_wb_clk_i _02796_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12027__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\] net737 net715 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\] net773 net713 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] _03815_ _03816_ vssd1 vssd1
+ vccd1 vccd1 _03822_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09082_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\] net890 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a22o_1
XANTENNA__10053__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08033_ _03744_ _03754_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__and2_1
XANTENNA__11849__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold800 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
Xinput60 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_1
Xinput71 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
Xhold811 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11538__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput82 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
Xinput93 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold822 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold866 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08954__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold877 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\] net924 net912 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1117_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08935_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04334_ vssd1 vssd1
+ vccd1 vccd1 _04452_ sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16414__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08866_ net1505 net1037 net1034 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07817_ _03505_ _03535_ _03538_ _03539_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__a2bb2o_1
X_08797_ team_02_WB.instance_to_wrap.top.pc\[0\] _04425_ _04357_ vssd1 vssd1 vccd1
+ vccd1 _04426_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout744_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] _03468_ _03469_ vssd1 vssd1
+ vccd1 vccd1 _03471_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09131__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16564__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07679_ _03367_ _03401_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout911_A _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09418_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\] net903 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\]
+ _04929_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__a221o_1
X_10690_ team_02_WB.instance_to_wrap.top.pc\[14\] _06197_ vssd1 vssd1 vccd1 vccd1
+ _06207_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09349_ _04865_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__inv_2
XANTENNA__13230__A2 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12360_ net297 net2595 net562 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__mux2_1
XANTENNA__10044__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09985__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] net494 _06812_ _04263_ net496
+ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__a221o_1
XANTENNA__11759__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12291_ net293 net2215 net569 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14030_ net1113 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09198__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11242_ _06745_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__inv_2
XANTENNA__09737__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11173_ _06181_ _06182_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input40_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\] net917 _05632_ _05633_
+ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a211o_1
X_15981_ clknet_leaf_33_wb_clk_i _02121_ _00789_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13297__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14932_ net1089 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
X_10055_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] net784 _05561_ _05564_
+ _05571_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09370__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ net1115 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16602_ clknet_leaf_89_wb_clk_i _02721_ _01395_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13814_ net1226 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__inv_2
X_14794_ net1143 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09122__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16533_ clknet_leaf_69_wb_clk_i net1022 _01340_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13745_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\]
+ _03245_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1
+ _03250_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10957_ net407 _06044_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15931__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16464_ clknet_leaf_77_wb_clk_i _02599_ _01272_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11480__A1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10283__A2 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13676_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _03208_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10888_ net405 _06350_ _06400_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15415_ clknet_leaf_116_wb_clk_i _01555_ _00223_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12627_ net2272 net318 net554 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__mux2_1
X_16395_ clknet_leaf_65_wb_clk_i _02530_ _01203_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11232__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10035__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15346_ clknet_leaf_85_wb_clk_i _01486_ _00159_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11232__B2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09976__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09928__A _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12558_ net296 net2136 net444 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11509_ net418 _06356_ _06607_ _07000_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_130_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15277_ clknet_leaf_74_wb_clk_i _01421_ _00090_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap542_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold107 net126 vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12489_ net294 net2516 net559 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold118 _02573_ vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09189__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold129 team_02_WB.START_ADDR_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09728__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14228_ net1077 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ net1115 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13288__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ _04328_ _04341_ _04345_ _04348_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__and4b_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15461__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1180 net1188 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__buf_4
Xfanout1191 net1197 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_4
X_08651_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] net998 vssd1 vssd1 vccd1
+ vccd1 _04280_ sky130_fd_sc_hd__nor2_4
XANTENNA__09900__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] team_02_WB.instance_to_wrap.top.a1.dataIn\[20\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1 vccd1 _03325_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08467__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11433__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10274__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09203_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\] net821 net813 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\]
+ _04719_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a221o_1
XANTENNA__14744__A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout325_A _06975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16810__1354 vssd1 vssd1 vccd1 vccd1 _16810__1354/HI net1354 sky130_fd_sc_hd__conb_1
XANTENNA_fanout1067_A _00018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ net968 _04650_ _04497_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10026__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09967__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09065_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\] net787 net779 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08016_ _03647_ _03660_ _03673_ _03645_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_113_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout694_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold663 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold685 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold696 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15804__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\] net768 net720 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__a22o_1
XANTENNA__13279__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13095__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net1045 _04209_ _04220_ net1008 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a32o_1
XANTENNA__12203__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\] net809 _05402_ _05414_
+ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__a211o_1
XANTENNA__09352__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ net145 net1040 net1035 net1479 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08418__A2_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14919__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15954__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ net320 net2192 net492 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07821__A team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ _06322_ _06326_ net370 vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__mux2_1
X_11791_ net314 net2630 net593 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08458__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13530_ _03073_ _03082_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10742_ team_02_WB.instance_to_wrap.top.pc\[11\] _06258_ vssd1 vssd1 vccd1 vccd1
+ _06259_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_81_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10673_ _06128_ _06189_ net791 _05625_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__o2bb2a_2
X_13461_ team_02_WB.START_ADDR_VAL_REG\[1\] net1068 net1002 vssd1 vssd1 vccd1 vccd1
+ net203 sky130_fd_sc_hd__a21o_1
XFILLER_0_137_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13203__A2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15200_ net1260 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
X_12412_ net251 net1833 net457 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__mux2_1
XANTENNA__09958__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16180_ clknet_leaf_10_wb_clk_i _02320_ _00988_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input88_A wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ team_02_WB.instance_to_wrap.ramload\[21\] net1012 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[21\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15334__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15131_ net1248 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
X_12343_ net241 net2002 net564 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15062_ net1259 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
X_12274_ net348 net2325 net576 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14013_ net1086 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
X_11225_ _05974_ _06599_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_75_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15484__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09591__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11156_ net391 _06662_ _06661_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13717__B _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10107_ net426 vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15964_ clknet_leaf_45_wb_clk_i _02104_ _00772_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11087_ _05948_ _05983_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12113__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08099__A team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14915_ net1130 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
X_10038_ _05540_ _05549_ _05552_ _05554_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__or4_2
X_15895_ clknet_leaf_116_wb_clk_i _02035_ _00703_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14829__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14846_ net1193 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14777_ net1129 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11989_ net285 net2426 net480 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16516_ clknet_leaf_37_wb_clk_i _02650_ _01323_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13728_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\] _03017_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__a21o_1
XANTENNA__10256__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16447_ clknet_leaf_103_wb_clk_i net1555 _01255_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13659_ net1465 net851 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11205__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10008__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16378_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[2\] _01186_
+ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15329_ clknet_leaf_46_wb_clk_i _01472_ _00142_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout406 _05900_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09582__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\] net770 net746 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a22o_1
Xfanout417 net419 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout439 net441 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_8
X_09752_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\] net715 _05266_ _05267_
+ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12023__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09334__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08703_ _04283_ net790 vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__nand2_1
X_09683_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\] net822 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\]
+ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout275_A _06740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08634_ net1062 net1060 team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04262_
+ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__and4b_2
XFILLER_0_96_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07641__A team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08565_ team_02_WB.instance_to_wrap.top.a1.row1\[63\] _04225_ _04233_ _04183_ vssd1
+ vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout442_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10247__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ team_02_WB.instance_to_wrap.top.a1.row1\[18\] _04186_ vssd1 vssd1 vccd1 vccd1
+ _04192_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12693__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout707_A _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09117_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\] net922 net910 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09048_ net972 net640 net545 vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13818__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net673 _06500_ _06501_ net672 _06521_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__a221o_1
Xhold482 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07816__A team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09573__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold493 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout940 net942 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout951 _04499_ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__buf_2
Xfanout962 _03027_ vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_4
Xfanout973 net976 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_4
Xfanout984 _02956_ vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout995 net996 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ team_02_WB.instance_to_wrap.top.pc\[10\] _05491_ vssd1 vssd1 vccd1 vccd1
+ _07481_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1160 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11772__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1171 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ net1071 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_87_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1182 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net249 net2696 net482 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__mux2_1
X_15680_ clknet_leaf_109_wb_clk_i _01820_ _00488_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1193 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ _07383_ _07411_ _07381_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__A team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14631_ net1117 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11843_ net252 net2342 net493 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11073__A _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10238__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14562_ net1205 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ net239 net1965 net593 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16301_ clknet_leaf_33_wb_clk_i _02441_ _01109_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13513_ _03072_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10725_ _03293_ _06130_ _06241_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16282__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14493_ net1084 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08851__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09478__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16232_ clknet_leaf_15_wb_clk_i _02372_ _01040_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13444_ _03028_ _03030_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10656_ team_02_WB.instance_to_wrap.top.pc\[24\] _06171_ vssd1 vssd1 vccd1 vccd1
+ _06173_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16163_ clknet_leaf_123_wb_clk_i _02303_ _00971_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13375_ team_02_WB.instance_to_wrap.ramload\[4\] net1010 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[4\] sky130_fd_sc_hd__and2_1
XANTENNA__12108__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10587_ _04458_ _04464_ _04467_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__and3_4
X_15114_ net1078 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
X_12326_ net309 net1912 net566 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16094_ clknet_leaf_113_wb_clk_i _02234_ _00902_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11947__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15045_ net1220 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
XANTENNA__12699__A0 _07051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12257_ net284 net2452 net575 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11208_ _05944_ _05974_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10734__D_N net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12188_ net278 net2066 net578 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_max_cap505_A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _04951_ _06601_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_121_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15947_ clknet_leaf_115_wb_clk_i _02087_ _00755_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15878_ clknet_leaf_42_wb_clk_i _02018_ _00686_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14829_ net1147 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XANTENNA_wire508_A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10229__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08350_ _04047_ _04058_ _04049_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_138_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11426__A1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09095__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08281_ _03975_ _03994_ _03952_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13179__B2 _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12018__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11857__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16005__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09555__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13357__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11362__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout247 _06372_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_1
X_09804_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\] net829 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__a22o_1
Xfanout258 _06530_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13639__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ _03716_ _03717_ _03713_ _03714_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__o211a_1
XANTENNA__16155__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09307__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ net612 _05251_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__nand2_1
XANTENNA__12688__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10997__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\] net755 net743 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__a22o_1
XANTENNA__11665__B2 _05556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08617_ net78 net1942 net955 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout824_A _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\] net835 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\]
+ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11417__A1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08548_ _04199_ _04200_ net653 net793 net1594 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09086__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ net1063 _04176_ _03317_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__or3b_1
XFILLER_0_33_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10510_ _04866_ _06026_ _04862_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11490_ _05558_ net658 vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire615 _04713_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_2
XFILLER_0_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire626 net627 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire637 _04732_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire648 _05898_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_2
X_10441_ _04693_ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09794__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10372_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\] net910 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__a22o_1
XANTENNA__13590__B2 team_02_WB.instance_to_wrap.top.a1.row2\[33\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13160_ net977 _07409_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12111_ net241 net1804 net468 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__mux2_1
XANTENNA__11767__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_13091_ team_02_WB.instance_to_wrap.top.pc\[20\] net1024 _02866_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12042_ _06280_ _07201_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__nor2_1
XANTENNA__09546__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold290 _02597_ vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16850_ net1394 vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_2
XFILLER_0_40_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout770 _04371_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_8
X_15801_ clknet_leaf_112_wb_clk_i _01941_ _00609_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout781 _04367_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_4
Xfanout792 _04326_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16781_ net1325 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_92_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13993_ net1101 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11105__B1 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12598__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15732_ clknet_leaf_12_wb_clk_i _01872_ _00540_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ team_02_WB.instance_to_wrap.top.pc\[18\] _06190_ vssd1 vssd1 vccd1 vccd1
+ _07464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15663_ clknet_leaf_38_wb_clk_i _01803_ _00471_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12875_ _07389_ _07393_ _07394_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11408__A1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14614_ net1093 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
X_11826_ net317 net2310 net589 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
XANTENNA__09077__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15594_ clknet_leaf_128_wb_clk_i _01734_ _00402_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14545_ net1105 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11757_ net304 net2673 net597 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__mux2_1
XANTENNA__08824__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10092__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10708_ team_02_WB.instance_to_wrap.top.pc\[20\] _06184_ vssd1 vssd1 vccd1 vccd1
+ _06225_ sky130_fd_sc_hd__xnor2_1
X_14476_ net1080 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
X_11688_ _07156_ _07161_ _07169_ _07173_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__o211a_1
XANTENNA__16028__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16215_ clknet_leaf_15_wb_clk_i _02355_ _01023_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13427_ _03036_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10639_ _04270_ _04288_ _04323_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09785__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16146_ clknet_leaf_6_wb_clk_i _02286_ _00954_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13358_ team_02_WB.instance_to_wrap.ramload\[20\] net1016 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[20\] sky130_fd_sc_hd__and2_1
XFILLER_0_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap948 _03355_ vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_1
X_12309_ _04291_ _04333_ _04452_ _06280_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__or4_2
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16077_ clknet_leaf_23_wb_clk_i _02217_ _00885_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13289_ team_02_WB.instance_to_wrap.top.pc\[15\] net1053 _06830_ net934 vssd1 vssd1
+ vccd1 vccd1 _02994_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16178__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15028_ net1204 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07850_ _03549_ _03568_ _03546_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__and3b_1
XANTENNA__10698__A2 _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07781_ _03303_ _03470_ net364 vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__nand3_1
XANTENNA__13097__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ net971 net633 net544 vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_1370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12301__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09451_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\] net723 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\]
+ _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08402_ _04102_ _04104_ _04108_ _04110_ _04097_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__a32o_4
XFILLER_0_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09382_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\] net927 net817 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\]
+ _04898_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__a221o_1
XANTENNA__09068__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08333_ _03993_ _04045_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08815__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10083__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08264_ _03972_ _03979_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08195_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout405_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1147_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09240__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13368__A team_02_WB.instance_to_wrap.ramload\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09528__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11335__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1009 _03314_ vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_2
XANTENNA_fanout774_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15545__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ _03677_ _03701_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09718_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\] net815 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\]
+ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__a221o_1
XANTENNA__11638__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12211__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15695__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ net396 _06288_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09700__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09649_ net969 _05164_ _04497_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input105_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12660_ net319 net1904 net434 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__mux2_1
XANTENNA__09059__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11611_ net377 _06502_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__or2_1
XANTENNA__08806__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13260__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12591_ net298 net2021 net439 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14330_ net1186 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
XANTENNA__10074__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ _06046_ _06048_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ net1185 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11473_ _06966_ _06967_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16000_ clknet_leaf_108_wb_clk_i _02140_ _00808_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input70_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ net633 net937 net1019 net1554 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__a2bb2o_1
X_10424_ _05212_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_55_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14192_ net1077 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
XANTENNA__09231__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13143_ _07412_ _02909_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__xnor2_1
X_10355_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\] net733 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09519__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13315__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10129__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13074_ _07458_ _07459_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__nor2_1
X_10286_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\] net920 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__a22o_1
XANTENNA__11326__B1 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12025_ net302 net2479 net476 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16833_ net1377 vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11629__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12121__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764_ net1308 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
X_13976_ net1104 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
XANTENNA__09298__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15715_ clknet_leaf_2_wb_clk_i _01855_ _00523_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12927_ team_02_WB.instance_to_wrap.top.pc\[29\] _06140_ vssd1 vssd1 vccd1 vccd1
+ _07447_ sky130_fd_sc_hd__or2_1
X_16695_ net138 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14837__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11960__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15646_ clknet_leaf_112_wb_clk_i _01786_ _00454_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12858_ net790 _04417_ _06127_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_17_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11809_ net254 net2028 net591 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15577_ clknet_leaf_17_wb_clk_i _01717_ _00385_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12789_ _06344_ _06398_ _06446_ _06477_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__and4_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14528_ net1155 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
XANTENNA__11262__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09470__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14459_ net1159 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09758__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09222__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12804__B _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15568__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16129_ clknet_leaf_119_wb_clk_i _02269_ _00937_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ _04463_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__nor2_1
XANTENNA__07617__C team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07902_ _03554_ _03570_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__or2_1
X_08882_ net14 net1030 net988 net2198 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09930__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _03555_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12031__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _03461_ _03462_ _03437_ _03441_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09289__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09503_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\] net799 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\]
+ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07695_ _03380_ _03417_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11870__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_A _07087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ _04948_ _04949_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_56_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\] net774 net710 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\]
+ _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1264_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10056__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08316_ _04028_ _04029_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__nor2_1
X_09296_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\] net918 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\]
+ _04803_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_30 _06914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16343__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09461__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08247_ _03938_ _03958_ _03960_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09749__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08178_ _03321_ _03896_ net2632 net1007 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout891_A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09213__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12206__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10140_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\] net781 net842 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
Xoutput192 net192 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_98_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10071_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\] net920 net884 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13830_ net1232 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13761_ net2726 net961 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10973_ _04778_ net662 _06484_ net796 vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_134_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14657__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11780__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15500_ clknet_leaf_25_wb_clk_i _01640_ _00308_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12712_ _07100_ _07113_ _07129_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__and3_1
XANTENNA__10295__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16480_ clknet_leaf_77_wb_clk_i net1704 _01288_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
X_13692_ net1589 _03216_ net1065 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_108_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15431_ clknet_leaf_29_wb_clk_i _01571_ _00239_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12643_ net251 net1711 net436 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ clknet_leaf_81_wb_clk_i _01502_ _00175_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12574_ net242 net2587 net440 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09452__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16721__1449 vssd1 vssd1 vccd1 vccd1 net1449 _16721__1449/LO sky130_fd_sc_hd__conb_1
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14313_ net1099 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ net407 _07016_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15293_ clknet_leaf_90_wb_clk_i _01437_ _00106_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14392__A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14244_ net1127 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
X_11456_ _06258_ _06951_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09204__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10407_ _05918_ _05923_ _05604_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o21ai_1
X_14175_ net1169 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XANTENNA__12116__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__A2 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11387_ team_02_WB.instance_to_wrap.top.pc\[12\] _06259_ team_02_WB.instance_to_wrap.top.pc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13126_ net978 _07417_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__o31ai_1
X_10338_ _05845_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_119_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10770__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13057_ net536 _06150_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10269_ _05740_ _05785_ net551 vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__mux2_1
X_12008_ _07190_ _07201_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__nor2_2
XANTENNA__09912__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16216__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16816_ net1360 vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__buf_2
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16747_ team_02_WB.instance_to_wrap.top.lcd.lcd_en vssd1 vssd1 vccd1 vccd1 net178
+ sky130_fd_sc_hd__clkbuf_1
X_13959_ net1239 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
XANTENNA__13472__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10286__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16678_ clknet_leaf_72_wb_clk_i _02795_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15629_ clknet_leaf_23_wb_clk_i _01769_ _00437_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13224__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09150_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\] net757 net677 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a22o_1
XANTENNA__09979__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ _03815_ _03816_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1
+ vccd1 vccd1 _03821_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15390__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09081_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\] net829 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\]
+ _04590_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08032_ _03711_ _03753_ _03706_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput50 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_1
XFILLER_0_4_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput61 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold801 team_02_WB.instance_to_wrap.ramload\[23\] vssd1 vssd1 vccd1 vccd1 net2259
+ sky130_fd_sc_hd__dlygate4sd3_1
Xinput72 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold812 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput83 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold834 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08403__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput94 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
Xmax_cap542 _04672_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_2
XANTENNA__12026__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold845 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold856 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\] net819 net799 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\]
+ _05499_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__a221o_1
Xhold889 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11865__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08934_ team_02_WB.instance_to_wrap.top.a1.row1\[101\] _03319_ vssd1 vssd1 vccd1
+ vccd1 _02515_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08865_ net138 _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout472_A _07208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] _03470_ _03506_ vssd1 vssd1
+ vccd1 vccd1 _03539_ sky130_fd_sc_hd__or3_1
X_08796_ _04423_ _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__and2_1
X_07747_ _03468_ _03469_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__or2_1
XANTENNA__12696__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07678_ _03393_ _03394_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] _03364_ vssd1
+ vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_32_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09682__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09417_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\] net830 net922 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\]
+ _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__a221o_1
XANTENNA__13215__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_A _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15733__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10029__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ _04863_ _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__and2b_2
XFILLER_0_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09279_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\] net703 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\]
+ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__a221o_1
XANTENNA__15101__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _06811_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07819__A team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12290_ net285 net2369 net571 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__mux2_1
XANTENNA__15883__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11241_ _06688_ _06744_ net371 vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10201__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11172_ _06677_ _06678_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16239__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ _05635_ _05636_ _05638_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__or4_1
XFILLER_0_101_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15980_ clknet_leaf_20_wb_clk_i _02120_ _00788_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14931_ net1168 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
X_10054_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\] net704 _05565_ _05567_
+ _05570_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10504__A1 _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14862_ net1113 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13813_ net1217 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__inv_2
X_16601_ clknet_leaf_97_wb_clk_i _02720_ _01394_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14793_ net1099 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16532_ clknet_leaf_59_wb_clk_i _00007_ _01339_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13744_ net2477 _03247_ _03249_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10956_ _06467_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__xor2_1
XFILLER_0_54_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09673__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16463_ clknet_leaf_72_wb_clk_i net1612 _01271_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08881__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13675_ _03206_ _03207_ net1241 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10887_ net383 _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15414_ clknet_leaf_57_wb_clk_i _01554_ _00222_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12626_ net2178 net313 net554 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__mux2_1
X_16394_ clknet_leaf_66_wb_clk_i _02529_ _01202_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09425__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15345_ clknet_leaf_84_wb_clk_i _01485_ _00158_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_12557_ net309 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\] net444 vssd1
+ vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11232__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11508_ net418 _06607_ _06608_ _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15276_ clknet_leaf_74_wb_clk_i _01420_ _00089_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12488_ net286 net2524 net559 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold108 _02622_ vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14227_ net1175 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
Xhold119 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ net945 _06931_ _06935_ net605 vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__o211a_2
XFILLER_0_125_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_max_cap535_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14850__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14158_ net1138 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13109_ team_02_WB.instance_to_wrap.top.pc\[17\] net1024 _02881_ _07337_ vssd1 vssd1
+ vccd1 vccd1 _01498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14089_ net1111 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15606__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire538_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1170 net1171 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08650_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] net1058 net997 _04277_
+ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__and4_1
Xfanout1181 net1188 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_2
Xfanout1192 net1197 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__buf_2
XFILLER_0_117_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07601_ _03322_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08581_ team_02_WB.instance_to_wrap.wb.curr_state\[0\] _04242_ vssd1 vssd1 vccd1
+ vccd1 _04243_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09664__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08872__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09202_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\] net829 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09416__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09133_ _04640_ _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__or2_4
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09064_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\] net767 _04571_ _04573_
+ _04580_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_103_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10982__A1 _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08015_ _03736_ _03734_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_128_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold620 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12184__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold642 team_02_WB.instance_to_wrap.ramaddr\[2\] vssd1 vssd1 vccd1 vccd1 net2100
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold664 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13376__A team_02_WB.instance_to_wrap.ramload\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout687_A _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold697 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09966_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\] net760 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a22o_1
XANTENNA__16531__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ net1507 _04440_ net930 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
XANTENNA__13684__B1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\] net926 net924 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\]
+ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout854_A _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16720__1448 vssd1 vssd1 vccd1 vccd1 net1448 _16720__1448/LO sky130_fd_sc_hd__conb_1
X_08848_ net146 net1040 net1036 net1569 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08779_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\] net762 net746 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10810_ _06324_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11790_ net306 net2024 net593 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__mux2_1
XANTENNA__09655__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10741_ team_02_WB.instance_to_wrap.top.pc\[10\] team_02_WB.instance_to_wrap.top.pc\[9\]
+ _06257_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13460_ team_02_WB.EN_VAL_REG net1069 net1003 _03060_ vssd1 vssd1 vccd1 vccd1 net192
+ sky130_fd_sc_hd__o31a_1
X_10672_ net994 _05669_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__nand2_1
XANTENNA__09407__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12411_ net239 net2185 net454 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13391_ team_02_WB.instance_to_wrap.ramload\[20\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[20\] sky130_fd_sc_hd__and2_1
XANTENNA__08652__B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15130_ net1248 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
X_12342_ _04292_ net647 _07193_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_11_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10973__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15061_ net1259 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12273_ net360 net2298 net575 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15629__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ net1151 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
XANTENNA__08918__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ net657 _06720_ _06728_ net796 _06725_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__o221a_1
XANTENNA__08918__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09040__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11155_ _04970_ net387 _06097_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__a21o_1
XANTENNA__13717__C net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\] net701 _05616_ _05621_
+ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a2111oi_2
X_11086_ net2453 net260 net641 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
X_15963_ clknet_leaf_127_wb_clk_i _02103_ _00771_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15779__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14914_ net1202 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
X_10037_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\] net819 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\]
+ _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__a221o_1
X_15894_ clknet_leaf_46_wb_clk_i _02034_ _00702_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09894__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14845_ net1084 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14776_ net1218 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
X_11988_ net272 net1754 net478 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09646__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13727_ net949 _03237_ _03238_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__and3_1
X_16515_ clknet_leaf_5_wb_clk_i _02649_ _01322_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08854__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10939_ net379 _06449_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14845__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16446_ clknet_leaf_103_wb_clk_i net1646 _01254_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_1
X_13658_ net1470 _04134_ net851 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12609_ net1952 net238 net554 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__mux2_1
XANTENNA__10584__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16377_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[1\] _01185_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[4\] sky130_fd_sc_hd__dfrtp_1
X_13589_ _03289_ net1047 _03142_ _03122_ team_02_WB.instance_to_wrap.top.a1.row2\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15328_ clknet_leaf_103_wb_clk_i _01471_ _00141_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15259_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[18\]
+ _00072_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_111_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09031__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout407 net409 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_2
X_09820_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\] net774 net722 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a22o_1
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12304__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10192__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\] net763 net711 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__a22o_1
X_08702_ net996 net792 vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__nor2_1
X_09682_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\] net923 net891 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__a22o_1
XANTENNA__09885__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ team_02_WB.instance_to_wrap.top.a1.instruction\[0\] team_02_WB.instance_to_wrap.top.a1.instruction\[1\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 _04262_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_102_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout268_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09098__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ _04227_ _04229_ _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09637__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08845__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08495_ team_02_WB.instance_to_wrap.top.a1.data\[10\] net958 _04190_ vssd1 vssd1
+ vccd1 vccd1 _04191_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout435_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1177_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout602_A _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09116_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\] net825 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\]
+ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09047_ _04546_ _04558_ _04561_ _04563_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__nor4_1
XFILLER_0_27_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold450 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold472 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08376__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12214__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold494 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10183__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout930 _04433_ vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_6
XFILLER_0_102_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout952 _04455_ vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_4
X_09949_ net516 _05464_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__and2_1
Xfanout963 _03027_ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout974 net976 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__clkbuf_4
Xfanout985 _02956_ vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 _04282_ vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ team_02_WB.instance_to_wrap.top.pc\[10\] _05491_ vssd1 vssd1 vccd1 vccd1
+ _07480_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09876__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11911_ net252 net1882 net484 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1161 team_02_WB.instance_to_wrap.ramaddr\[11\] vssd1 vssd1 vccd1 vccd1 net2619
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _07384_ _07410_ _07385_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__o21ba_1
Xhold1194 team_02_WB.instance_to_wrap.top.a1.row2\[33\] vssd1 vssd1 vccd1 vccd1 net2652
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ net1083 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11842_ net237 net2497 net490 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09089__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09628__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07639__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ net1209 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
XANTENNA__15301__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ net245 net2440 net594 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13512_ team_02_WB.instance_to_wrap.top.pad.keyCode\[6\] team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] team_02_WB.instance_to_wrap.top.pad.keyCode\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__or4b_1
X_16300_ clknet_leaf_20_wb_clk_i _02440_ _01108_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ _06132_ _06240_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_82_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14492_ net1146 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ clknet_leaf_29_wb_clk_i _02371_ _01039_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13443_ _03033_ _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10655_ _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16162_ clknet_leaf_122_wb_clk_i _02302_ _00970_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15451__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13374_ team_02_WB.instance_to_wrap.ramload\[3\] net1010 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[3\] sky130_fd_sc_hd__and2_1
X_10586_ net668 _06102_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nor2_1
XANTENNA__09800__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15113_ net1098 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
X_12325_ net300 net2436 net566 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__mux2_1
X_16093_ clknet_leaf_49_wb_clk_i _02233_ _00901_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15044_ net1195 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
X_12256_ net274 net2527 net573 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__mux2_1
XANTENNA__08602__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11207_ net2357 net289 net643 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12187_ net280 net1649 net578 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__mux2_1
XANTENNA__12124__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ net657 _06637_ _06642_ _06645_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__o211a_1
XANTENNA__11963__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15946_ clknet_leaf_0_wb_clk_i _02086_ _00754_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ net398 _06578_ _06575_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_30_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09867__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ clknet_leaf_32_wb_clk_i _02017_ _00685_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14828_ net1071 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09619__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08827__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14759_ net1112 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08280_ _03952_ _03975_ _03994_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_28_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13179__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16429_ clknet_leaf_65_wb_clk_i net1558 _01237_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10608__A _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09252__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16734__1458 vssd1 vssd1 vccd1 vccd1 net1458 _16734__1458/LO sky130_fd_sc_hd__conb_1
XANTENNA__12034__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10165__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 _03859_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11362__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09803_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\] net906 net805 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\]
+ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__a221o_1
Xfanout237 net240 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_2
X_07995_ _03716_ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__nor2_1
Xfanout259 _06530_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout385_A _05901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ net970 _05250_ net543 vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09665_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\] net731 net723 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\]
+ _05181_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__a221o_1
XANTENNA__15324__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ net79 net1563 net954 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
X_09596_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\] net920 net900 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08547_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.row1\[111\]
+ net794 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__mux2_1
XANTENNA__08818__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15474__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _00017_ _03317_ _04175_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__and3_2
XFILLER_0_107_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12209__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire627 _05332_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire649 _05645_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_2
X_10440_ _04630_ _04651_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10371_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\] net813 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\]
+ _05883_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12110_ net647 _07210_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_57_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ _04280_ _02864_ _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12041_ net347 net2435 net474 vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__mux2_1
Xhold280 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\] vssd1 vssd1
+ vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10156__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout760 _04374_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_6
XANTENNA__11783__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout771 _04371_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_4
X_15800_ clknet_leaf_19_wb_clk_i _01940_ _00608_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout782 _04366_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13992_ net1177 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
X_16780_ net1324 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12302__A0 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout793 _04223_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__buf_2
XANTENNA__09849__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__A team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15731_ clknet_leaf_55_wb_clk_i _01871_ _00539_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12943_ team_02_WB.instance_to_wrap.top.pc\[19\] _06188_ vssd1 vssd1 vccd1 vccd1
+ _07463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12874_ _05742_ _05781_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__xnor2_2
X_15662_ clknet_leaf_11_wb_clk_i _01802_ _00470_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11825_ net313 net1987 net589 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
X_14613_ net1215 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
XANTENNA__08809__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15593_ clknet_leaf_103_wb_clk_i _01733_ _00401_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14544_ net1076 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
X_11756_ net298 net2257 net598 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__mux2_1
XANTENNA__09482__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10707_ team_02_WB.instance_to_wrap.top.pc\[19\] _06186_ _06223_ vssd1 vssd1 vccd1
+ vccd1 _06224_ sky130_fd_sc_hd__a21oi_1
X_14475_ net1203 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11687_ _04569_ _04589_ _04608_ _07170_ _07172_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__o311a_1
XANTENNA__12119__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16214_ clknet_leaf_45_wb_clk_i _02354_ _01022_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13426_ _03289_ net962 _03035_ net1242 vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__a211o_2
X_10638_ _04272_ _04277_ net1059 vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13030__A1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11958__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16145_ clknet_leaf_50_wb_clk_i _02285_ _00953_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13357_ team_02_WB.instance_to_wrap.ramload\[19\] net1016 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[19\] sky130_fd_sc_hd__and2_1
X_10569_ net408 _06078_ _06083_ net380 vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ net344 net2044 net569 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__mux2_1
X_16076_ clknet_leaf_20_wb_clk_i _02216_ _00884_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13288_ team_02_WB.instance_to_wrap.ramaddr\[16\] net983 net964 _02993_ vssd1 vssd1
+ vccd1 vccd1 _01435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15027_ net1218 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12239_ net2165 net354 net618 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10147__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07780_ _03303_ net364 _03470_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_15929_ clknet_leaf_18_wb_clk_i _02069_ _00737_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\] net735 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08401_ _04096_ _04098_ _04094_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a21o_1
X_09381_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\] net883 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08332_ _03306_ _03990_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08734__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08263_ _03306_ _03974_ _03977_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__and3_1
XANTENNA__12029__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09225__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08194_ _03823_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11868__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13649__A _00018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1042_A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13368__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10138__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__A1 _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12532__A0 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09862__A _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12699__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout767_A _04372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ _03668_ _03699_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10801__A _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__A _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\] net916 net804 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11638__A2 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16695__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08503__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ net969 _05164_ _04497_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10310__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09579_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\] net756 _05094_ _05095_
+ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a211o_1
X_11610_ _05999_ _07097_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__nand2_1
XANTENNA__15104__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12590_ net311 net2529 net440 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09464__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11541_ _05912_ _05916_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__xor2_1
XANTENNA__10074__B2 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ net1074 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ net664 _06956_ _06965_ net656 _06958_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__o221a_1
XANTENNA__09216__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13211_ _04990_ net936 net1020 net1523 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11778__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _05935_ _05938_ _05252_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__o21a_1
X_14191_ net1111 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11574__A1 _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10377__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13142_ _07379_ _07380_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input63_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\] net785 net777 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\]
+ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09519__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11079__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13315__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ net1027 _02851_ net1024 team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1
+ vccd1 vccd1 _01504_ sky130_fd_sc_hd__a2bb2o_1
X_10285_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\] net811 net884 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\]
+ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12024_ net295 net1977 net475 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16832_ net1376 vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_2
XANTENNA__12402__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13079__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout590 net592 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16763_ net1307 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
X_13975_ net1236 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15714_ clknet_leaf_124_wb_clk_i _01854_ _00522_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12926_ team_02_WB.instance_to_wrap.top.pc\[29\] _06140_ vssd1 vssd1 vccd1 vccd1
+ _07446_ sky130_fd_sc_hd__nand2_1
X_16694_ net138 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10301__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10857__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15645_ clknet_leaf_49_wb_clk_i _01785_ _00453_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _05355_ _06205_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11808_ net238 net2238 net589 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12788_ _06508_ _06541_ _06573_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__and3_1
XANTENNA__09455__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15576_ clknet_leaf_18_wb_clk_i _01716_ _00384_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16733__1457 vssd1 vssd1 vccd1 vccd1 net1457 _16733__1457/LO sky130_fd_sc_hd__conb_1
XANTENNA__10065__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09012__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11739_ _06282_ net2032 net600 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14527_ net1176 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16145__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09207__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458_ net1184 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13409_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__or4b_1
XFILLER_0_40_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14389_ net1185 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
XANTENNA__10368__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16128_ clknet_leaf_107_wb_clk_i _02268_ _00936_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08950_ _04276_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__nand2_4
XANTENNA__13306__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16059_ clknet_leaf_127_wb_clk_i _02199_ _00867_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12514__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ _03562_ _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08881_ net15 net1032 net989 team_02_WB.instance_to_wrap.ramload\[21\] vssd1 vssd1
+ vccd1 vccd1 _02549_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07832_ _03520_ _03554_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12312__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10621__A team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ _03461_ _03462_ _03437_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09502_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\] net823 net819 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07694_ _03345_ _03347_ _03361_ _03351_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ _04928_ _04947_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout250_A _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09364_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\] net758 net730 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09446__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08315_ _04000_ _04002_ _04018_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__and3_1
X_09295_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\] net903 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\]
+ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a221o_1
XANTENNA_20 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 _06914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1257_A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _03961_ _03959_ _03932_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__mux2_2
XFILLER_0_69_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15512__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ _03888_ _03893_ _03862_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_63_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10764__C1 team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout884_A _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_100_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XANTENNA__15662__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput193 net193 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
X_10070_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\] net876 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\]
+ _05586_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12222__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10531__A _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16018__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13760_ _03065_ _03258_ _03259_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10972_ _06029_ _06467_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13481__A1 team_02_WB.START_ADDR_VAL_REG\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09685__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ _06125_ _07234_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11492__B1 _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13691_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\] _03216_ vssd1 vssd1 vccd1
+ vccd1 _03217_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15430_ clknet_leaf_44_wb_clk_i _01570_ _00238_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ net238 net1825 net434 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__mux2_1
XANTENNA__09437__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16168__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15361_ clknet_leaf_91_wb_clk_i _01501_ _00174_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_12573_ net646 _07207_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14673__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14312_ net1176 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
X_11524_ _06978_ _07015_ net365 vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__mux2_1
X_15292_ clknet_leaf_75_wb_clk_i _01436_ _00105_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08671__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14243_ net1145 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11455_ team_02_WB.instance_to_wrap.top.pc\[9\] _06257_ team_02_WB.instance_to_wrap.top.pc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10406_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__inv_2
X_14174_ net1194 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11386_ team_02_WB.instance_to_wrap.top.pc\[12\] _06205_ _06203_ vssd1 vssd1 vccd1
+ vccd1 _06885_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_123_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13125_ net229 _02893_ _06861_ net233 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08963__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10337_ _05847_ _05849_ _05851_ _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__or4_1
XFILLER_0_81_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10770__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13056_ _06560_ net234 vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10268_ team_02_WB.instance_to_wrap.top.a1.instruction\[14\] net651 _05784_ vssd1
+ vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12007_ net346 net2057 net478 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12132__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ net969 _05695_ _05714_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__o21ai_1
X_16815_ net1359 vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__buf_2
XANTENNA__14848__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11971__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16746_ net1291 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__09676__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13958_ net1239 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09140__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12909_ _07364_ _07428_ _07363_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__a21oi_1
X_16677_ clknet_leaf_72_wb_clk_i _02794_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13889_ net1253 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11272__A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15628_ clknet_leaf_10_wb_clk_i _01768_ _00436_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09428__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13224__B2 _05555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15535__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15559_ clknet_leaf_24_wb_clk_i _01699_ _00367_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08100_ _03818_ _03819_ _03799_ _03817_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\] net918 net910 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\]
+ _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08031_ _03740_ _03741_ _03743_ _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__o31a_1
Xinput40 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13199__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12307__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput51 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11538__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold802 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
Xinput62 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11211__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap510 net511 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_68_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput73 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
Xinput84 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15685__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold813 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput95 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold824 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09600__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold835 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold846 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold868 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09982_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\] net892 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a22o_1
Xhold879 team_02_WB.instance_to_wrap.top.pad.keyCode\[6\] vssd1 vssd1 vccd1 vccd1
+ net2337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12831__A _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07925__A team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08933_ net1499 _04451_ net930 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout298_A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08864_ net139 net1038 net1034 net1538 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1005_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ _03532_ _03533_ _03507_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a21oi_1
X_08795_ net549 _04422_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__nand2_1
XANTENNA__11881__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07746_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] _03461_ _03462_ vssd1 vssd1
+ vccd1 vccd1 _03469_ sky130_fd_sc_hd__and3_1
XANTENNA__09667__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09131__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07677_ _03364_ _03396_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__xor2_2
XFILLER_0_95_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08475__B team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09416_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\] net899 net875 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09419__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13215__B2 _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09347_ net532 _04861_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14493__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\] net727 net719 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08229_ _03916_ _03926_ _03918_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12217__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11240_ _06333_ _06336_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__nand2_1
XANTENNA__09198__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10960__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11171_ net838 _06658_ _06660_ net670 vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10122_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\] net921 net877 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\]
+ _05634_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__a221o_1
X_16732__1456 vssd1 vssd1 vccd1 vccd1 net1456 _16732__1456/LO sky130_fd_sc_hd__conb_1
X_14930_ net1119 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\] net788 _05568_ _05569_
+ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__a211o_1
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14861_ net1140 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11791__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16600_ clknet_leaf_97_wb_clk_i _02719_ _01393_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13812_ net1217 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14792_ net1178 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
XANTENNA__08666__A team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09658__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16531_ clknet_leaf_69_wb_clk_i net1462 _01338_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09122__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15558__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13743_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\] _03247_ net950 vssd1
+ vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__a21boi_1
X_10955_ _04777_ _05954_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16462_ clknet_leaf_78_wb_clk_i net1748 _01270_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__xnor2_1
X_10886_ net408 _06400_ _06352_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08881__B2 team_02_WB.instance_to_wrap.ramload\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15413_ clknet_leaf_39_wb_clk_i _01553_ _00221_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12625_ net2314 net306 net554 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__mux2_1
X_16393_ clknet_leaf_65_wb_clk_i _02528_ _01201_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ net302 net2294 net444 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15344_ clknet_leaf_84_wb_clk_i _01484_ _00157_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08605__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11507_ net376 _06820_ _06999_ _06084_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12127__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15275_ clknet_leaf_77_wb_clk_i _01419_ _00088_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12487_ net273 net2184 net557 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold109 net157 vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09189__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14226_ net1118 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11438_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _06833_ _06934_ vssd1 vssd1
+ vccd1 vccd1 _06935_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11966__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ net1133 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
X_11369_ _06062_ _06064_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13108_ _02878_ _02879_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__o21ai_1
X_14088_ net1176 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ _07449_ _07450_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09897__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16333__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1160 net1161 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09361__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1171 net1198 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_2
Xfanout1182 net1188 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__buf_4
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14578__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1196 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_4
X_07600_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] team_02_WB.instance_to_wrap.top.a1.dataIn\[26\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] team_02_WB.instance_to_wrap.top.a1.dataIn\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__or4_1
X_08580_ team_02_WB.instance_to_wrap.Wen team_02_WB.instance_to_wrap.Ren vssd1 vssd1
+ vccd1 vccd1 _04242_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09649__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16729_ net1453 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_49_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16483__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08872__B2 team_02_WB.instance_to_wrap.ramload\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09201_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\] net898 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\]
+ _04717_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_100_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ _04642_ _04644_ _04646_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09821__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\] net743 _04574_ _04576_
+ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_5_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12037__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ _03736_ _03734_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10982__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold610 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold621 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold632 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11876__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold643 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10780__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold654 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10195__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1
+ net2134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold698 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09965_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\] net732 _05471_ _05474_
+ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout582_A _07209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ net1045 _04206_ _04217_ net1008 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__a32o_1
XANTENNA__09888__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09896_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\] net892 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09352__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ net147 net1040 net1036 net1715 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13392__A team_02_WB.instance_to_wrap.ramload\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08778_ _04358_ _04363_ _04364_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__and3_1
XANTENNA__12500__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09104__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ _03416_ _03449_ _03451_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ team_02_WB.instance_to_wrap.top.pc\[8\] _06256_ vssd1 vssd1 vccd1 vccd1 _06257_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_32_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10671_ net791 _05580_ _06127_ _06187_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__o22a_4
XFILLER_0_14_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12410_ net246 net2658 net456 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13390_ team_02_WB.instance_to_wrap.ramload\[19\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[19\] sky130_fd_sc_hd__and2_1
XFILLER_0_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09812__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12341_ net346 net2132 net565 vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15060_ net1238 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
X_12272_ net353 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\] net575 vssd1
+ vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11786__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14011_ net1157 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11223_ _06727_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10186__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15230__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__A2 _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07565__A team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09591__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ net370 _06604_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10105_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\] net713 net697 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11085_ net607 _06589_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__and3_4
X_15962_ clknet_leaf_120_wb_clk_i _02102_ _00770_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09879__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14913_ net1207 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
X_10036_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\] net924 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15893_ clknet_leaf_43_wb_clk_i _02033_ _00701_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15380__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12410__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14844_ net1152 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
XANTENNA__08396__A team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14775_ net1174 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11987_ net289 net2012 net480 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__mux2_1
X_16514_ clknet_leaf_37_wb_clk_i _02648_ _01321_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13726_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\] _03017_ vssd1 vssd1 vccd1
+ vccd1 _03238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10938_ _05715_ _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16445_ clknet_leaf_103_wb_clk_i net1672 _01253_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10869_ net388 _06050_ _06383_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__a21oi_1
X_13657_ net1473 _04143_ net851 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12608_ net2131 net246 net553 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13060__C1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16376_ clknet_leaf_93_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[0\] _01184_
+ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09803__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ net1050 team_02_WB.instance_to_wrap.top.a1.row1\[121\] _03115_ _03290_ vssd1
+ vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_41_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15327_ clknet_leaf_104_wb_clk_i _01470_ _00140_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12539_ net345 net2492 net446 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15258_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[17\]
+ _00071_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14209_ net1209 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15189_ net1256 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire550_A _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09582__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire648_A _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 net409 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_2
Xfanout419 net420 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_103_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15723__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\] net759 net731 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09334__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ _04275_ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__or2_2
XANTENNA__09690__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ _05191_ _05193_ _05195_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08632_ net72 net1541 net956 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__mux2_1
XANTENNA__13416__S _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12320__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15873__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08563_ _03313_ net1046 vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_102_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10101__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08494_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[10\] net980 vssd1 vssd1 vccd1
+ vccd1 _04190_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout330_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1072_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16731__1455 vssd1 vssd1 vccd1 vccd1 net1455 _16731__1455/LO sky130_fd_sc_hd__conb_1
XFILLER_0_31_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09115_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\] net918 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09046_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\] net908 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\]
+ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout797_A _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold440 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10168__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10804__A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold451 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10707__A2 _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold484 team_02_WB.START_ADDR_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09573__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold495 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16779__1323 vssd1 vssd1 vccd1 vccd1 _16779__1323/HI net1323 sky130_fd_sc_hd__conb_1
XANTENNA_fanout964_A _02957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10523__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16698__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 _04515_ vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__buf_6
XANTENNA__13106__B1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout931 net932 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08781__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout942 _04532_ vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
X_09948_ net514 _05464_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__nor2_1
Xfanout953 _04455_ vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11117__C1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout964 _02957_ vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_4
Xfanout975 net976 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_2
Xfanout986 _02956_ vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\] net782 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1140 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1151 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15107__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net240 net2204 net482 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12230__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1173 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _05534_ _05537_ _07409_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1184 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 team_02_WB.instance_to_wrap.ramaddr\[28\] vssd1 vssd1 vccd1 vccd1 net2653
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ net245 net1956 net490 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13850__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11772_ net241 net2295 net596 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__mux2_1
X_14560_ net1148 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08944__A _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11840__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10723_ _06135_ _06239_ _06137_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__a21oi_1
X_13511_ team_02_WB.instance_to_wrap.top.pad.keyCode\[2\] team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] team_02_WB.instance_to_wrap.top.pad.keyCode\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__or4b_2
XFILLER_0_3_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14491_ net1184 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16230_ clknet_leaf_42_wb_clk_i _02370_ _01038_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input93_A wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10654_ _06168_ _06170_ _06167_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__a21o_2
X_13442_ _02764_ _02763_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__nor2_1
XANTENNA__13042__C1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13593__B1 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13373_ net1807 net1011 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[2\]
+ sky130_fd_sc_hd__and2_1
X_16161_ clknet_leaf_121_wb_clk_i _02301_ _00969_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10585_ net423 _06071_ net374 _06101_ _06086_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15112_ net1078 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
XANTENNA__09775__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12324_ net294 net2515 net567 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__mux2_1
X_16092_ clknet_leaf_44_wb_clk_i _02232_ _00900_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15043_ net1221 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
X_12255_ net290 net2381 net575 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10159__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12405__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206_ net946 _06705_ _06711_ net606 vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__o211a_2
X_12186_ net269 net1735 net578 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08772__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ _04951_ net665 _06643_ net796 _06644_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_125_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13648__A1 team_02_WB.instance_to_wrap.top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15896__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09316__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15945_ clknet_leaf_106_wb_clk_i _02085_ _00753_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11068_ net369 _06510_ _06577_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_121_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] _04326_ net652 _05535_
+ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_30_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12140__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10331__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15876_ clknet_leaf_2_wb_clk_i _02016_ _00684_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14827_ net1206 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14758_ net1075 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11831__A0 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13709_ _03227_ _03228_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14689_ net1208 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11280__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16428_ clknet_leaf_64_wb_clk_i net1667 _01236_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16359_ clknet_leaf_31_wb_clk_i _02499_ _01167_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12315__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09555__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08763__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\] net898 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout238 net240 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dlymetal6s2s_1
X_07994_ _03692_ net255 _03686_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__a21oi_1
Xfanout249 _06498_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09307__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ _05240_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__nor2_4
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout378_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12050__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\] net751 net735 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10322__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ net80 net1498 net956 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09595_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\] net819 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\]
+ _05111_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08546_ net1590 net793 net653 _04197_ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a22o_1
XANTENNA__08279__C1 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15619__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08477_ _04175_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout712_A _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire628 net629 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire639 _04607_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_126_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09794__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10370_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\] net817 net906 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\]
+ _05884_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_76_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12733__B _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\] net828 net808 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\]
+ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_72_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12225__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ net348 net2137 net477 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__mux2_1
XANTENNA__09546__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 team_02_WB.instance_to_wrap.top.a1.row1\[59\] vssd1 vssd1 vccd1 vccd1 net1728
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08004__A team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold281 team_02_WB.START_ADDR_VAL_REG\[23\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 team_02_WB.instance_to_wrap.top.a1.row2\[9\] vssd1 vssd1 vccd1 vccd1 net1750
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13845__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_127_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08939__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout750 _04376_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout761 _04374_ vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_4
Xfanout772 _04371_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__clkbuf_8
X_13991_ net1105 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
Xfanout783 _04366_ vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08506__B1 _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11105__A2 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout794 _04223_ vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11365__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15730_ clknet_leaf_5_wb_clk_i _01870_ _00538_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12942_ team_02_WB.instance_to_wrap.top.pc\[20\] _06186_ vssd1 vssd1 vccd1 vccd1
+ _07462_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15661_ clknet_leaf_23_wb_clk_i _01801_ _00469_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12873_ _07390_ _07392_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15299__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14612_ net1075 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11824_ net304 net2743 net589 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15592_ clknet_leaf_19_wb_clk_i _01732_ _00400_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10616__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14543_ net1115 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
X_11755_ net309 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\] net600 vssd1
+ vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10092__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ _06222_ _06221_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_1508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14474_ net1142 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11686_ _05966_ _07157_ _07171_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__nand3_1
X_16213_ clknet_leaf_42_wb_clk_i _02353_ _01021_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13425_ team_02_WB.instance_to_wrap.top.lcd.currentState\[3\] net962 vssd1 vssd1
+ vccd1 vccd1 _03035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10637_ _06153_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16144_ clknet_leaf_40_wb_clk_i _02284_ _00952_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11041__A1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13356_ team_02_WB.instance_to_wrap.ramload\[18\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[18\] sky130_fd_sc_hd__and2_1
X_10568_ net424 net413 vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09785__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__B2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08613__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13318__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12307_ net348 net2144 net571 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__mux2_1
XANTENNA__12135__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16075_ clknet_leaf_114_wb_clk_i _02215_ _00883_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13287_ team_02_WB.instance_to_wrap.top.pc\[16\] net1052 _06807_ net934 vssd1 vssd1
+ vccd1 vccd1 _02993_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10499_ _05986_ _05987_ _05989_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15026_ net1218 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09537__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12238_ net2468 net356 net616 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap510_A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12169_ net332 net2043 net464 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16730__1454 vssd1 vssd1 vccd1 vccd1 net1454 _16730__1454/LO sky130_fd_sc_hd__conb_1
XFILLER_0_21_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15928_ clknet_leaf_18_wb_clk_i _02068_ _00736_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10304__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09170__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10855__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15859_ clknet_leaf_56_wb_clk_i _01999_ _00667_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08400_ _04102_ _04104_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__and3_1
X_09380_ _04890_ _04892_ _04894_ _04896_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08331_ _04024_ _04042_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15911__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16778__1322 vssd1 vssd1 vccd1 vccd1 _16778__1322/HI net1322 sky130_fd_sc_hd__conb_1
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10083__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08262_ _03974_ _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_95_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08193_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] _03858_ vssd1 vssd1 vccd1
+ vccd1 _03911_ sky130_fd_sc_hd__or2_1
XANTENNA__12834__A _04631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13309__B1 _07046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12045__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09528__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11884__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16417__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1202_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _03668_ _03699_ _03666_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout662_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09716_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\] net928 net812 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\]
+ _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15441__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09647_ _05156_ _05160_ _05162_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__or4_4
XANTENNA__14496__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09578_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\] net728 net720 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a22o_1
X_08529_ net1046 _04214_ _04215_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13260__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10529__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11540_ _05916_ _06003_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10074__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11471_ net416 net666 _06536_ _06963_ net795 vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_59_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15120__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13210_ net1585 net1021 net938 _04946_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a22o_1
X_10422_ _05292_ _05935_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ net1138 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13141_ net791 _07332_ _07510_ _02907_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a211o_1
X_10353_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\] net757 net728 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11079__B _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13072_ _06623_ net234 _02848_ net979 _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__o221a_1
XANTENNA__09519__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input56_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\] net924 net807 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a22o_1
XANTENNA__16097__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11326__A2 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12023_ net284 net2752 net475 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
XANTENNA__11794__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16831_ net1375 vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_2
XFILLER_0_121_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13079__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _07214_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_4
Xfanout591 net592 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_8
XFILLER_0_73_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16762_ net1306 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
X_13974_ net1257 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15713_ clknet_leaf_117_wb_clk_i _01853_ _00521_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12925_ team_02_WB.instance_to_wrap.top.pc\[30\] _06134_ vssd1 vssd1 vccd1 vccd1
+ _07445_ sky130_fd_sc_hd__nand2_1
X_16693_ clknet_leaf_74_wb_clk_i _02810_ _01417_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15644_ clknet_leaf_45_wb_clk_i _01784_ _00452_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _05314_ _06200_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_17_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11807_ net246 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\] net590 vssd1
+ vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15575_ clknet_leaf_13_wb_clk_i _01715_ _00383_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12787_ _06903_ _07308_ _07309_ _07310_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__nor4_1
XFILLER_0_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14526_ net1190 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11262__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ _04291_ net645 _07190_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__or3_4
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11969__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14457_ net1139 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
X_11669_ _05271_ _05290_ _05990_ _07154_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07748__A team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13408_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\] _03019_ vssd1 vssd1 vccd1
+ vccd1 _03020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09758__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14388_ net1075 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
XANTENNA__15314__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08966__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16127_ clknet_leaf_86_wb_clk_i _02267_ _00935_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13339_ net2067 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[1\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_110_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10174__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16058_ clknet_leaf_120_wb_clk_i _02198_ _00866_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11317__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07900_ _03521_ _03553_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__and2_1
X_15009_ net1229 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ net16 net1029 net987 net2655 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_88_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07831_ _03519_ _03552_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09930__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07762_ _03481_ _03483_ _03484_ _03476_ _03461_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a32o_1
XANTENNA__09143__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\] net912 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__a22o_1
X_07693_ _03384_ _03411_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08497__A2 _04185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09432_ net614 _04947_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__nand2_2
XFILLER_0_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08518__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09363_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\] net726 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\]
+ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout243_A _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10056__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ _04000_ _04018_ _04002_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12450__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\] net910 net856 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_10 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_32 _06914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11879__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ _03929_ _03959_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_43 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1152_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12202__A0 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ _03852_ _03861_ _03889_ _03856_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08957__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1260_A team_02_WB.START_ADDR_VAL_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XANTENNA_fanout877_A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_101_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__12503__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput194 net194 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XANTENNA__09382__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11627__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10531__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15957__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _06084_ _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13481__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15115__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12710_ _04325_ _06161_ _06249_ _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__o31a_1
XFILLER_0_35_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10295__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ net1240 _03215_ _03216_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__nor3_1
XFILLER_0_6_1614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12641_ net244 net1721 net435 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10047__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15360_ clknet_leaf_90_wb_clk_i _01500_ _00173_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12572_ net345 net1852 net442 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14311_ net1101 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
XANTENNA__11789__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11523_ net426 net384 _06297_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__a21o_1
X_15291_ clknet_leaf_81_wb_clk_i _01435_ _00104_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08671__B team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16849__1393 vssd1 vssd1 vccd1 vccd1 _16849__1393/HI net1393 sky130_fd_sc_hd__conb_1
X_14242_ net1202 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
X_11454_ net669 _06937_ _06949_ net837 _06947_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ _05919_ _05920_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__nand2_1
X_14173_ net1086 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11385_ net952 _06883_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13124_ _07375_ _07416_ _07374_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10336_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\] net800 net861 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\]
+ _05852_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10267_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] net997 _04329_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__a22o_1
X_13055_ team_02_WB.instance_to_wrap.top.pc\[26\] net1025 _02836_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01507_ sky130_fd_sc_hd__a22o_1
XANTENNA__12413__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16777__1321 vssd1 vssd1 vccd1 vccd1 _16777__1321/HI net1321 sky130_fd_sc_hd__conb_1
X_12006_ net348 net2591 net481 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XANTENNA__09373__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10198_ net969 _05695_ _05714_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__o21a_2
XFILLER_0_94_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16814_ net1358 vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__buf_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09125__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16745_ net1290 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
X_13957_ net1239 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13472__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12908_ _04971_ _06180_ _07427_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15025__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10286__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16676_ clknet_leaf_72_wb_clk_i _02793_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13888_ net1256 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_128_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15627_ clknet_leaf_115_wb_clk_i _01767_ _00435_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12839_ _04802_ _06150_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__nand2_1
XANTENNA__13224__A2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15558_ clknet_leaf_42_wb_clk_i _01698_ _00366_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09979__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14509_ net1140 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
XANTENNA__16262__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15489_ clknet_leaf_121_wb_clk_i _01629_ _00297_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_08030_ net2206 net1007 net982 _03752_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput52 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_1
Xinput63 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11538__A2 _07026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_1
Xhold803 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput74 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
Xhold814 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap522 net523 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_2
Xhold825 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08403__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput85 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
Xinput96 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
Xhold836 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09693__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold847 team_02_WB.START_ADDR_VAL_REG\[27\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10210__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold858 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\] net811 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\]
+ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold869 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12499__A0 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] net1009 _04232_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10632__A team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12323__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ net150 net1039 net1035 net1666 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08102__A team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07814_ _03499_ _03536_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__xor2_2
XANTENNA__13943__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08794_ net549 _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__or2_1
XANTENNA__09116__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07745_ _03461_ _03462_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1
+ vccd1 vccd1 _03468_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout458_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07676_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] _03396_ _03397_ vssd1 vssd1
+ vccd1 vccd1 _03399_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09415_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\] net911 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13215__A2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10029__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ net532 _04861_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\] net695 _04784_ _04787_
+ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08228_ _03943_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11529__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08159_ _03865_ _03867_ _03876_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07602__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10201__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11170_ _06672_ _06675_ _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\] net905 net807 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\]
+ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12233__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09355__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\] net736 net716 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__a22o_1
XANTENNA__13151__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14860_ net1080 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09107__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ net1217 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__inv_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ net1105 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08666__B team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ clknet_leaf_69_wb_clk_i net1485 _01337_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13742_ _03247_ _03248_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__nor2_1
X_10954_ _04734_ _04778_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__or2_2
XFILLER_0_97_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16461_ clknet_leaf_74_wb_clk_i net1690 _01269_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13673_ net1644 _03206_ net1240 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a21oi_1
X_10885_ net390 _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15412_ clknet_leaf_12_wb_clk_i _01552_ _00220_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12624_ net1827 net299 net553 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16392_ clknet_leaf_91_wb_clk_i _02527_ _01200_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15343_ clknet_leaf_84_wb_clk_i _01483_ _00156_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ net292 net2307 net442 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ _06920_ _06998_ net394 vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__mux2_1
X_15274_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_read_i _00087_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.Ren sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12486_ net290 net1758 net559 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14225_ net1120 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11437_ team_02_WB.instance_to_wrap.top.pc\[11\] net973 _06933_ net1001 _06837_ vssd1
+ vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09594__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14156_ net1082 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08621__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ _06014_ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13107_ net229 _02877_ _06786_ net233 vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__o2bb2a_1
X_10319_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14087_ net1111 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XANTENNA__10452__A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11299_ net377 _06571_ _06639_ _06567_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13038_ _06460_ net234 vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11982__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 net1153 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1161 net1162 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__buf_2
Xfanout1172 net1174 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1183 net1188 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_4
Xfanout1194 net1196 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__buf_4
XANTENNA_wire426_A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09649__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14989_ net1222 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16628__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10259__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16728_ net1452 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_44_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16659_ clknet_leaf_100_wb_clk_i _02778_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08872__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09200_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\] net914 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08592__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09131_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\] net898 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\]
+ _04647_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12318__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09062_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\] net722 _04577_ _04578_
+ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_96_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08013_ _03708_ _03735_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold622 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold633 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold644 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold655 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold666 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold677 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12053__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\] net845 _05475_ _05477_
+ _05480_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a2111o_1
Xhold699 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1115_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09337__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ net1508 _04439_ net930 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
X_09895_ _05406_ _05408_ _05410_ _05411_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__or4_1
Xhold1300 team_02_WB.instance_to_wrap.ramload\[13\] vssd1 vssd1 vccd1 vccd1 net2758
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout575_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08846_ net148 net1037 net1034 net1671 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16848__1392 vssd1 vssd1 vccd1 vccd1 _16848__1392/HI net1392 sky130_fd_sc_hd__conb_1
XFILLER_0_135_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\] net766 _04388_ _04393_
+ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout742_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__A _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07728_ _03445_ _03450_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07659_ _03353_ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10670_ net994 _05625_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_81_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\] net863 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\]
+ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__a221o_1
X_16776__1320 vssd1 vssd1 vccd1 vccd1 _16776__1320/HI net1320 sky130_fd_sc_hd__conb_1
XANTENNA__12228__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12340_ net350 net2688 net568 vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12271_ net358 net2123 net573 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14010_ net1186 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11222_ net417 _06726_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__nor2_1
XANTENNA__09040__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ _04997_ _06659_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09328__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\] net781 _05617_ _05620_
+ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11084_ net975 _06593_ _06592_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15961_ clknet_leaf_17_wb_clk_i _02101_ _00769_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14679__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15525__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14912_ net1155 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
X_10035_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\] net908 _05538_ _05551_
+ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15892_ clknet_leaf_12_wb_clk_i _02032_ _00700_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08677__A _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ net1157 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11438__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ net1095 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
XANTENNA__15675__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11986_ net278 net2172 net479 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16513_ clknet_leaf_7_wb_clk_i _02647_ _01320_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13725_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\] _03017_ vssd1 vssd1 vccd1
+ vccd1 _03237_ sky130_fd_sc_hd__or2_1
XANTENNA__10110__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ net410 _06449_ _06359_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08854__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16444_ clknet_leaf_64_wb_clk_i net1716 _01252_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
X_13656_ _04153_ net851 _03196_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10868_ net365 _06055_ _06056_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__and3_1
XANTENNA__08616__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12607_ net1709 net243 net555 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16375_ clknet_leaf_96_wb_clk_i _02515_ _01183_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[101\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_45_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12138__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ team_02_WB.instance_to_wrap.top.a1.row2\[25\] _03118_ _03128_ team_02_WB.instance_to_wrap.top.a1.row1\[105\]
+ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10799_ net542 net386 _06314_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15326_ clknet_leaf_103_wb_clk_i _01469_ _00139_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12538_ net349 net2330 net449 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11977__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15257_ clknet_leaf_66_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[16\]
+ _00070_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_12469_ net357 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\] net450 vssd1
+ vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap638_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09567__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14208_ net1154 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10177__A1 _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15188_ net1256 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09031__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14139_ net1180 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout409 _05809_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_39_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09319__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13115__B2 _07337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16450__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ net1060 _04267_ net977 vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_20_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09680_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\] net919 net899 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\]
+ _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__a221o_1
XANTENNA__12601__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08631_ net83 net1543 net954 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08562_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04175_ vssd1 vssd1 vccd1
+ vccd1 _04231_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_102_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09098__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08493_ _04171_ _04185_ _04188_ _04189_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a31o_1
XANTENNA__12837__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08526__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12048__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1065_A _00018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09114_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11601__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09270__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11887__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\] net901 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1232_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09558__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold430 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\] vssd1
+ vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold441 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15548__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold485 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout910 _04523_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout921 _04515_ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout932 _04335_ vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_2
X_09947_ _05444_ net624 net969 vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__mux2_1
Xfanout943 _04501_ vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout954 _04261_ vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14499__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout957_A _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 _02957_ vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout976 _04284_ vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__buf_2
XANTENNA__12511__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout987 net988 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__buf_2
X_09878_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\] net746 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10820__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1130 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout998 net1000 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 team_02_WB.instance_to_wrap.ramload\[24\] vssd1 vssd1 vccd1 vccd1 net2599
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09730__B1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08829_ net1689 net1042 net992 team_02_WB.instance_to_wrap.ramaddr\[2\] vssd1 vssd1
+ vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
Xhold1152 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 team_02_WB.instance_to_wrap.top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 net2632
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ net243 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\] net493 vssd1
+ vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09089__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11771_ _04291_ _04333_ net646 _06280_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__or4_2
XANTENNA__13290__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08944__B _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ net1685 net1460 _03071_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10722_ team_02_WB.instance_to_wrap.top.pc\[28\] _06140_ _06238_ vssd1 vssd1 vccd1
+ vccd1 _06239_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14490_ net1180 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13441_ net1065 _03028_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__and2_1
X_10653_ team_02_WB.instance_to_wrap.top.a1.instruction\[24\] _04283_ _06169_ vssd1
+ vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14962__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16160_ clknet_leaf_113_wb_clk_i _02300_ _00968_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input86_A wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13372_ net2067 net1011 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[1\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_24_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16323__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10584_ _06093_ _06100_ net400 vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15111_ net1108 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
XANTENNA__11797__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12323_ net285 net2061 net567 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16091_ clknet_leaf_126_wb_clk_i _02231_ _00899_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09549__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15042_ net1195 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
X_12254_ net278 net1934 net573 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11205_ net974 _06710_ _06709_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__a21o_1
XANTENNA__16473__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12185_ net263 net2553 net578 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11136_ _04948_ net662 net659 _04949_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_53_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12421__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ net370 _06576_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__nand2_1
X_15944_ clknet_leaf_16_wb_clk_i _02084_ _00752_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09721__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ _04421_ _05441_ net551 vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__mux2_1
X_15875_ clknet_leaf_125_wb_clk_i _02015_ _00683_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14826_ net1142 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ net1126 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
XANTENNA__08827__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11969_ net358 net2048 net585 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13708_ net1729 _03226_ net1065 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14688_ net1158 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11280__B _06782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16427_ clknet_leaf_103_wb_clk_i net1539 _01235_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
X_13639_ net1571 net962 _03187_ net1067 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16358_ clknet_leaf_50_wb_clk_i _02498_ _01166_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09252__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15309_ clknet_leaf_64_wb_clk_i _01452_ _00122_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16289_ clknet_leaf_117_wb_clk_i _02429_ _01097_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16847__1391 vssd1 vssd1 vccd1 vccd1 _16847__1391/HI net1391 sky130_fd_sc_hd__conb_1
XFILLER_0_48_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10624__B _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09801_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\] net809 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\]
+ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09960__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 net231 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_4
X_07993_ _03686_ _03692_ net255 vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__and3_1
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_108_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13639__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09732_ _05242_ _05244_ _05246_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_108_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12331__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14112__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09663_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\] net771 _05170_ _05173_
+ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_97_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout273_A _06740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08614_ net81 team_02_WB.START_ADDR_VAL_REG\[18\] net954 vssd1 vssd1 vccd1 vccd1
+ _02646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13951__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09594_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\] net928 net908 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ net1662 net793 net653 _04194_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
XANTENNA__13272__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout440_A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__A0 _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16346__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ _04169_ _04174_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__and2_1
XANTENNA__09491__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13024__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10087__A _05579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09779__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire629 _05289_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12506__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09028_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\] net917 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_57_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold260 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1
+ net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1
+ net1729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_8
Xfanout751 _04376_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15118__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12241__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout762 net765 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_8
Xfanout773 _04371_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10550__A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ net1072 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
Xfanout784 _04366_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_6
XFILLER_0_137_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09703__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout795 net796 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_4
X_12941_ team_02_WB.instance_to_wrap.top.pc\[20\] _06186_ vssd1 vssd1 vccd1 vccd1
+ _07461_ sky130_fd_sc_hd__nor2_1
XANTENNA__14957__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15660_ clknet_leaf_25_wb_clk_i _01800_ _00468_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12872_ _07389_ _07391_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14611_ net1166 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11823_ net296 net2063 net590 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15591_ clknet_leaf_26_wb_clk_i _01731_ _00399_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08809__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14542_ net1164 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11754_ net302 net2361 net598 vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09482__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ team_02_WB.instance_to_wrap.top.pc\[19\] _06186_ vssd1 vssd1 vccd1 vccd1
+ _06222_ sky130_fd_sc_hd__xnor2_1
X_14473_ net1109 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XANTENNA__15713__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11685_ _04672_ _04692_ _05967_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16212_ clknet_leaf_11_wb_clk_i _02352_ _01020_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13424_ _03030_ _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10636_ _04344_ _04349_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__or2_1
XANTENNA__09234__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12924__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16143_ clknet_leaf_36_wb_clk_i _02283_ _00951_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13355_ team_02_WB.instance_to_wrap.ramload\[17\] net1014 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[17\] sky130_fd_sc_hd__and2_1
XFILLER_0_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11041__A2 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12416__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ net416 net412 vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__nor2_2
XFILLER_0_45_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13318__B2 _03008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12306_ net360 net1992 net571 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__mux2_1
X_16074_ clknet_leaf_130_wb_clk_i _02214_ _00882_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15863__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13286_ net1772 net986 net967 _02992_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10498_ _05991_ _06013_ _05990_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__o21a_1
X_15025_ net1213 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
X_12237_ net2554 net342 net618 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10396__A_N net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10001__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12168_ net333 net2368 net464 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16219__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ _04951_ _05947_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12151__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12099_ net1777 net327 net582 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_15927_ clknet_leaf_14_wb_clk_i _02067_ _00735_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11990__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15243__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16369__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15858_ clknet_leaf_5_wb_clk_i _01998_ _00666_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire506_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14809_ net1138 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15789_ clknet_leaf_24_wb_clk_i _01929_ _00597_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10068__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08330_ _04024_ _04035_ _04040_ _04039_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15393__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ _03952_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08192_ _03872_ _03896_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09225__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12834__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12326__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13309__B2 _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1028_A _07337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09933__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout390_A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A _07198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12061__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _03660_ _03664_ _03673_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__o21ba_1
X_09715_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\] net889 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09646_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\] net900 net799 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\]
+ _05147_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__a221o_1
XANTENNA__10846__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09577_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\] net772 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout822_A _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08528_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[2\] net980 vssd1 vssd1 vccd1
+ vccd1 _04215_ sky130_fd_sc_hd__or2_2
XANTENNA__10529__B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09464__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08459_ _03307_ _04154_ _04160_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire426 net427 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__dlymetal6s2s_1
X_11470_ net375 _06773_ _06961_ net382 _06964_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09216__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11559__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10421_ _05292_ _05936_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__or2_1
XANTENNA__12236__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10545__A _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08975__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10231__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ _07479_ _07481_ _07509_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__nor3_1
XANTENNA__08975__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10352_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\] net761 _05858_ _05861_
+ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_103_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13071_ net229 _02849_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__nand2_1
XANTENNA__13180__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__A _04694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\] net941 _05796_ _05797_
+ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ net274 net2350 net474 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__mux2_1
XANTENNA_input49_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16830_ net1374 vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_2
XANTENNA__15266__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 _07217_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_4
Xfanout581 _07209_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_8
Xfanout592 _07194_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13195__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16761_ net1305 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
X_13973_ net1255 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
XANTENNA__10298__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ team_02_WB.instance_to_wrap.top.pc\[30\] _06134_ vssd1 vssd1 vccd1 vccd1
+ _07444_ sky130_fd_sc_hd__or2_1
X_15712_ clknet_leaf_108_wb_clk_i _01852_ _00520_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_16692_ clknet_leaf_77_wb_clk_i _02809_ _01416_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08685__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16846__1390 vssd1 vssd1 vccd1 vccd1 _16846__1390/HI net1390 sky130_fd_sc_hd__conb_1
XFILLER_0_38_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15643_ clknet_leaf_128_wb_clk_i _01783_ _00451_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12855_ _05314_ _06200_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11806_ net242 net2459 net591 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15574_ clknet_leaf_48_wb_clk_i _01714_ _00382_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12786_ _06722_ _06753_ _06770_ _06802_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09455__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14525_ net1086 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
X_11737_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] _04333_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__or3b_2
XFILLER_0_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11262__A2 _06759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14456_ net1220 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
XANTENNA__13133__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11668_ _05993_ _07152_ _07153_ _05991_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__a31o_1
XANTENNA__09207__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13407_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__and2_1
X_10619_ _06135_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__inv_2
XANTENNA__12146__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ net1169 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
X_11599_ net2062 net354 net643 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16126_ clknet_leaf_109_wb_clk_i _02266_ _00934_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13338_ net1731 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[0\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_45_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10174__B _05690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11985__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16057_ clknet_leaf_111_wb_clk_i _02197_ _00865_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13269_ team_02_WB.instance_to_wrap.top.pc\[25\] net1054 net935 _02983_ vssd1 vssd1
+ vccd1 vccd1 _02984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15008_ net1229 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15609__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09915__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07830_ _03511_ _03519_ _03534_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07761_ _03453_ _03463_ _03480_ _03448_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a22o_1
XANTENNA__15759__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__inv_2
X_07692_ _03414_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ net614 _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09362_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\] net762 net734 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a22o_1
XANTENNA__09446__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08313_ _04025_ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__or2_1
X_09293_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\] net814 net863 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\]
+ _04807_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11253__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12845__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_33 _07069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ net2652 net1007 net982 _03960_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_44 _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08534__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08175_ _03888_ _03862_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12056__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1145_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10213__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11895__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XANTENNA__15289__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XANTENNA__07674__A team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09906__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XANTENNA__11713__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout772_A _04371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput195 net195 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
X_07959_ _03652_ _03655_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__and2_1
XANTENNA__13466__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09134__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ net398 _06106_ _06480_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_98_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09685__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\] net728 _05141_ _05142_
+ _05145_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_6_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12640_ net243 net2551 net436 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input103_A wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09437__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ net350 net2292 net445 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14310_ net1089 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11522_ _05649_ _06004_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__xor2_1
X_15290_ clknet_leaf_75_wb_clk_i _01434_ _00103_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08671__C team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ net1159 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
X_11453_ _05927_ _06948_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10404_ _05579_ _05603_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__or2_1
XANTENNA__10204__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14172_ net1151 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11384_ net669 _06867_ _06882_ net837 _06880_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__o221a_2
XFILLER_0_110_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13123_ _07513_ _02892_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__xnor2_1
X_10335_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\] net929 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13054_ net979 _07435_ _02834_ _02835_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__o31ai_1
X_10266_ net412 _05782_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__nand2_1
X_12005_ net362 net1764 net480 vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XANTENNA__15901__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10197_ net970 net621 vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__or2_1
X_16813_ net1357 vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16744_ net1289 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XANTENNA__14210__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ net1239 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
XANTENNA__09676__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13209__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ _07365_ _07367_ _07425_ _06184_ _05017_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__a32o_1
X_16675_ clknet_leaf_72_wb_clk_i _02792_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13887_ net1255 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12838_ net539 _06147_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__xor2_1
X_15626_ clknet_leaf_129_wb_clk_i _01766_ _00434_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09428__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15557_ clknet_leaf_35_wb_clk_i _01697_ _00365_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12769_ net664 _07177_ _07292_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14508_ net1072 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
X_15488_ clknet_leaf_109_wb_clk_i _01628_ _00296_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_14439_ net1112 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14880__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput42 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput53 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_1
XANTENNA__15431__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput64 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_1
Xmax_cap512 _05533_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09061__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput75 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
Xhold804 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16557__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput86 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
Xhold815 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09600__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold826 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xinput97 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
X_16109_ clknet_leaf_24_wb_clk_i _02249_ _00917_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold848 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12604__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09980_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\] net916 net908 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold859 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08931_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] net959 _04221_ _04173_ vssd1
+ vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_1619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15581__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08862_ net1557 net1040 net1036 team_02_WB.instance_to_wrap.ramstore\[2\] vssd1 vssd1
+ vccd1 vccd1 _02564_ sky130_fd_sc_hd__a22o_1
XANTENNA__11171__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07813_ _03532_ _03533_ _03502_ _03510_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08793_ net652 _04420_ _04421_ net792 vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_100_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07744_ _03435_ _03463_ _03464_ _03466_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09667__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07675_ _03396_ _03397_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout353_A _07087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09414_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\] net927 net810 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1095_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09419__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ _04842_ _04861_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout618_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1262_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09276_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\] net759 _04789_ _04790_
+ _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_106_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08227_ _03909_ _03915_ _03926_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08158_ _03876_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07602__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12514__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08089_ _03755_ _03786_ _03782_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__o21a_2
XFILLER_0_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10823__A _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15924__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10120_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\] net913 _04550_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10051_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\] net768 net740 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__a22o_1
XANTENNA__13151__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13810_ net1228 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14790_ net1083 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09658__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13741_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] _03245_ net950 vssd1 vssd1
+ vccd1 vccd1 _03248_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10953_ net1816 net254 net643 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10673__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16460_ clknet_leaf_74_wb_clk_i net1634 _01268_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
X_13672_ _03202_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\] _03200_ _03205_
+ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__or4bb_2
X_10884_ _06080_ _06081_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12623_ net2217 net308 net556 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__mux2_1
X_15411_ clknet_leaf_54_wb_clk_i _01551_ _00219_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16391_ clknet_leaf_92_wb_clk_i _02526_ _01199_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15342_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] _00155_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[3\] sky130_fd_sc_hd__dfrtp_1
X_12554_ net285 net1737 net443 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
XANTENNA__09291__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10976__A1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09830__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ _06959_ _06997_ net365 vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__mux2_1
X_15273_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_write_i _00086_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.Wen sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12485_ net278 net2273 net557 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__mux2_1
XANTENNA__12178__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224_ net1109 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
X_11436_ _06259_ _06932_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__nor2_1
XANTENNA__09043__B1 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14155_ net1200 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12424__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11367_ _05377_ _06013_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _07369_ _07370_ _07421_ net978 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ net792 _05442_ _05834_ net652 vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__a22oi_4
X_14086_ net1089 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11298_ _05207_ net662 net659 _05210_ _06799_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__a221o_1
XANTENNA__10452__B _04733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ _02821_ _02818_ _07349_ team_02_WB.instance_to_wrap.top.pc\[29\] vssd1 vssd1
+ vccd1 vccd1 _01510_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_123_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10249_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\] net704 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09897__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1140 net1143 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__buf_4
Xfanout1151 net1152 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__buf_4
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1162 net1198 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__clkbuf_2
Xfanout1173 net1174 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_4
XANTENNA__10900__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10900__B2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1184 net1188 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__buf_4
Xfanout1195 net1196 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11564__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14988_ net1228 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09649__A2 _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16727_ net1451 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13939_ net1257 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
XANTENNA__08857__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16869__1413 vssd1 vssd1 vccd1 vccd1 _16869__1413/HI net1413 sky130_fd_sc_hd__conb_1
X_16658_ clknet_leaf_101_wb_clk_i _02777_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08609__A0 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15609_ clknet_leaf_17_wb_clk_i _01749_ _00417_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16589_ clknet_leaf_99_wb_clk_i _02708_ _01382_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08592__B net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09130_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\] net805 net886 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09282__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10627__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09821__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09061_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\] net715 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12169__A0 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ _03694_ net255 _03680_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_128_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09034__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold601 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\] vssd1 vssd1
+ vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12842__B _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold623 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold634 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1
+ net2092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12334__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10643__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold645 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold656 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10195__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16825__1369 vssd1 vssd1 vccd1 vccd1 _16825__1369/HI net1369 sky130_fd_sc_hd__conb_1
Xhold667 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold678 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\] net788 _05478_ _05479_
+ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__a211o_1
Xhold689 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13954__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08914_ net1045 _04203_ _04214_ net1008 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout1010_A _03014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\] net870 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\]
+ _05403_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1108_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1301 team_02_WB.instance_to_wrap.ramload\[16\] vssd1 vssd1 vccd1 vccd1 net2759
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ net149 net1038 net1033 net1645 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11695__A2 _07138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout470_A _07208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08776_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\] net782 _04396_ _04398_
+ _04404_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a2111o_1
X_07727_ _03410_ net425 _03415_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08848__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14785__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout735_A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07658_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] _03349_ vssd1 vssd1 vccd1
+ vccd1 _03381_ sky130_fd_sc_hd__nand2_1
XANTENNA__15477__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout902_A _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07589_ team_02_WB.instance_to_wrap.top.a1.state\[2\] _03313_ vssd1 vssd1 vccd1 vccd1
+ _03314_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09328_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\] net915 net903 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08076__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09273__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09259_ net972 _04774_ net544 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12270_ net343 net2563 net576 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__mux2_1
X_11221_ net414 _06483_ _06717_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13235__B1_N net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12244__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12580__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16102__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11152_ _05042_ _06600_ _05039_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__o21a_1
XANTENNA__08023__A team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10103_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\] net749 _05618_ _05619_
+ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11083_ _06173_ _06231_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__xnor2_1
X_15960_ clknet_leaf_54_wb_clk_i _02100_ _00768_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09879__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ net1170 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
X_10034_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\] net892 net807 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\]
+ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__a221o_1
X_15891_ clknet_leaf_85_wb_clk_i _02031_ _00699_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ net1180 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11438__A2 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11985_ net282 net2065 net479 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14773_ net1185 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
XANTENNA_output118_A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16512_ clknet_leaf_28_wb_clk_i _02646_ _01319_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13724_ _03018_ net950 _03236_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__and3_1
X_10936_ net410 _06449_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16443_ clknet_leaf_63_wb_clk_i net1570 _01251_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10867_ _06378_ _06380_ net392 vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__mux2_1
X_13655_ net1477 net851 vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__nor2_1
XANTENNA__12419__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10728__A _06244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12606_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] net646 _06277_ _06279_
+ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__and4_1
X_16374_ clknet_leaf_47_wb_clk_i _02514_ _01182_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13060__A1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13586_ team_02_WB.instance_to_wrap.top.a1.row1\[113\] _03121_ _03124_ team_02_WB.instance_to_wrap.top.a1.row2\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13060__B2 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ _04714_ net386 vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__nor2_1
XANTENNA__09803__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11071__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ net361 net2623 net449 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
X_15325_ clknet_leaf_86_wb_clk_i _01468_ _00138_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15256_ clknet_leaf_66_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[15\]
+ _00069_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_12468_ net341 net1814 net453 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__mux2_1
XANTENNA__08632__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14207_ net1176 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
X_11419_ _06011_ net664 vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12154__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15187_ net1255 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
X_12399_ net334 net2093 net460 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ net1183 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
XANTENNA__11993__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13115__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ net1216 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
XANTENNA_wire536_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08630_ net94 net2718 net954 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08561_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04175_ vssd1 vssd1 vccd1
+ vccd1 _04230_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08492_ team_02_WB.instance_to_wrap.top.a1.row1\[19\] _04186_ vssd1 vssd1 vccd1 vccd1
+ _04189_ sky130_fd_sc_hd__and2_1
XANTENNA__10101__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12837__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_112_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12329__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09255__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09113_ _04623_ _04629_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_115_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13949__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__A _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\] net892 _04551_ _04560_
+ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a211o_1
XANTENNA__16125__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold420 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12064__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold431 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10168__A2 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1225_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold453 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold464 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold475 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold486 team_02_WB.instance_to_wrap.ramload\[31\] vssd1 vssd1 vccd1 vccd1 net1944
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout900 _04526_ vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout911 _04523_ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_4
Xhold497 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout922 _04513_ vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08781__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09946_ _05456_ _05459_ _05461_ _05462_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_70_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout933 net935 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11117__A1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 _04500_ vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__buf_2
Xfanout955 _04261_ vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_2
Xfanout966 _02957_ vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_4
Xfanout977 _04281_ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__buf_4
X_09877_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\] net690 _05382_ _05393_
+ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__a211o_1
Xhold1120 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\] vssd1 vssd1 vccd1 vccd1
+ net2578 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout988 _04432_ vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
Xhold1131 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ net1747 net1041 net990 team_02_WB.instance_to_wrap.ramaddr\[3\] vssd1 vssd1
+ vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
Xhold1153 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1175 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1 net2655
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\] net714 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11770_ net346 net2049 net597 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13290__A1 team_02_WB.instance_to_wrap.ramaddr\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09494__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13290__B2 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10721_ _06145_ _06237_ _06141_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12239__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10548__A _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13440_ _03034_ _03041_ _03042_ _03045_ _03046_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10652_ net996 _04492_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13042__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09246__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13042__B2 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13371_ net1731 net1010 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[0\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_49_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10583_ _06096_ _06099_ net371 vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15110_ net1098 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12322_ net272 net2054 net565 vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16090_ clknet_leaf_119_wb_clk_i _02230_ _00898_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input79_A wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15041_ net1204 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
X_12253_ net282 net2114 net574 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__mux2_1
XANTENNA__10159__A2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11204_ _06224_ _06225_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12184_ net267 net2336 net578 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16868__1412 vssd1 vssd1 vccd1 vccd1 _16868__1412/HI net1412 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_129_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11135_ net423 _06634_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__nand2_1
XANTENNA__08772__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12702__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11108__A1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11108__B2 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15642__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13648__A3 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11066_ _06321_ _06324_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__nor2_1
X_15943_ clknet_leaf_27_wb_clk_i _02083_ _00751_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10730__B net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ net511 vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ clknet_leaf_122_wb_clk_i _02014_ _00682_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10331__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14825_ net1099 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
XANTENNA__15792__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08627__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14756_ net1130 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
XANTENNA__09485__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ net342 net1945 net588 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16824__1368 vssd1 vssd1 vccd1 vccd1 _16824__1368/HI net1368 sky130_fd_sc_hd__conb_1
XFILLER_0_131_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13707_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\] _03226_ vssd1 vssd1 vccd1
+ vccd1 _03227_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_47_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10919_ _06293_ _06299_ net365 vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__mux2_1
XANTENNA__12149__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14687_ net1189 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
X_11899_ net338 net2290 net489 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16426_ clknet_leaf_67_wb_clk_i _02561_ _01234_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_28_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16148__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13638_ _03109_ _03113_ _03117_ team_02_WB.instance_to_wrap.top.a1.row1\[60\] _03023_
+ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_15_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11988__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16357_ clknet_leaf_35_wb_clk_i _02497_ _01165_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13569_ net1047 net1049 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] _03103_
+ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08870__B net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12792__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15308_ clknet_leaf_103_wb_clk_i _01451_ _00121_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16288_ clknet_leaf_113_wb_clk_i _02428_ _01096_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15239_ clknet_leaf_70_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[30\]
+ _00052_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09800_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\] net914 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__a22o_1
XANTENNA__08763__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07992_ _03713_ _03714_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__nand2_1
XANTENNA__12612__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout229 net231 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08598__A _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09731_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\] net826 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\]
+ _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09662_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\] net844 _05175_ _05176_
+ _05178_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10322__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ net82 net1574 net954 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
X_09593_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\] net799 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\]
+ _05105_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__a221o_1
XANTENNA__10973__A2_N net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout266_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08544_ net1584 net793 _04224_ _04191_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10086__A1 _05602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] team_02_WB.instance_to_wrap.top.a1.halfData\[2\]
+ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 _04174_
+ sky130_fd_sc_hd__nand3b_1
XANTENNA_fanout433_A _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12059__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11898__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13285__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout600_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_76_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09027_ _04516_ _04527_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11338__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15665__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold250 team_02_WB.START_ADDR_VAL_REG\[10\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold261 team_02_WB.instance_to_wrap.top.a1.row1\[56\] vssd1 vssd1 vccd1 vccd1 net1719
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 net186 vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 team_02_WB.instance_to_wrap.ramload\[9\] vssd1 vssd1 vccd1 vccd1 net1741
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold294 team_02_WB.instance_to_wrap.top.a1.row2\[3\] vssd1 vssd1 vccd1 vccd1 net1752
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12522__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 net733 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__clkbuf_8
Xfanout741 _04379_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_4
XANTENNA__08939__C _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\] net827 net823 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a22o_1
Xfanout752 _04376_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__buf_6
Xfanout763 net765 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_4
Xfanout774 net777 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_8
Xfanout785 _04366_ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08506__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout796 _06105_ vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__clkbuf_4
X_12940_ team_02_WB.instance_to_wrap.top.pc\[21\] _06184_ vssd1 vssd1 vccd1 vccd1
+ _07460_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11510__B2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12871_ _05788_ _05828_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15134__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ net1124 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
X_11822_ net308 net1674 net590 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15590_ clknet_leaf_44_wb_clk_i _01730_ _00398_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09467__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13263__B2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11274__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14541_ net1141 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
X_11753_ net295 net2645 net599 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10704_ team_02_WB.instance_to_wrap.top.pc\[18\] _06188_ _06220_ vssd1 vssd1 vccd1
+ vccd1 _06221_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ net1176 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
XANTENNA__09219__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11684_ _04781_ _05968_ _05969_ _06373_ _07158_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_37_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16211_ clknet_leaf_53_wb_clk_i _02351_ _01019_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ team_02_WB.instance_to_wrap.top.pc\[25\] _06150_ vssd1 vssd1 vccd1 vccd1
+ _06152_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ net1065 _03028_ _03031_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11577__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13354_ net1653 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[16\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16142_ clknet_leaf_8_wb_clk_i _02282_ _00950_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10566_ net369 _06079_ _06080_ _06082_ net399 vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__o311a_1
XFILLER_0_63_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11041__A3 _06549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ net355 net2239 net571 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13318__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16073_ clknet_leaf_118_wb_clk_i _02213_ _00881_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13285_ _06782_ _02959_ team_02_WB.instance_to_wrap.top.pc\[17\] net1053 vssd1 vssd1
+ vccd1 vccd1 _02992_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_121_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10497_ _05336_ _05932_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__nor2_1
XANTENNA__11329__A1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12236_ net1908 net337 net619 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__mux2_1
X_15024_ net1213 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12940__B _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ net328 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\] net464 vssd1
+ vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__mux2_1
XANTENNA__12432__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11118_ net2659 net271 net641 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12098_ net2678 net322 net581 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
X_15926_ clknet_leaf_46_wb_clk_i _02066_ _00734_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11049_ _06268_ _06559_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10304__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09170__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15857_ clknet_leaf_23_wb_clk_i _01997_ _00665_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14808_ net1194 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XANTENNA__09458__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15788_ clknet_leaf_25_wb_clk_i _01928_ _00596_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14739_ net1166 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
XANTENNA__15538__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14883__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08260_ _03925_ _03960_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16409_ clknet_leaf_66_wb_clk_i _02544_ _01217_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08191_ _03868_ _03905_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12607__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09630__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13309__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12850__B _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14123__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09217__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ _03684_ _03693_ _03697_ _03680_ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__a211o_1
XFILLER_0_96_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout383_A _06084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09714_ net612 vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__inv_2
XANTENNA__09697__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16313__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10797__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09645_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\] net835 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\]
+ _05161_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09576_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\] net841 _05090_ _05092_
+ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08527_ team_02_WB.instance_to_wrap.top.a1.data\[2\] net958 vssd1 vssd1 vccd1 vccd1
+ _04214_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16867__1411 vssd1 vssd1 vccd1 vccd1 _16867__1411/HI net1411 sky130_fd_sc_hd__conb_1
XFILLER_0_33_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout815_A _04521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ net1620 net1005 net982 _04161_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11008__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12517__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08389_ _04094_ _04096_ _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__a21oi_4
Xwire427 net428 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_59_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11559__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10420_ _05936_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09621__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10545__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10351_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\] net781 _05862_ _05864_
+ _05867_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13070_ _07457_ _07527_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__xnor2_1
X_10282_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\] net815 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\]
+ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12021_ net289 net2428 net474 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09924__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16823__1367 vssd1 vssd1 vccd1 vccd1 _16823__1367/HI net1367 sky130_fd_sc_hd__conb_1
XANTENNA__12252__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout560 _07223_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_4
Xfanout571 _07217_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_8
X_16760_ net1304 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
Xfanout582 _07209_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_4
Xfanout593 net596 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_6
X_13972_ net1255 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09152__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15711_ clknet_leaf_110_wb_clk_i _01851_ _00519_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12923_ _07441_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__xnor2_1
X_16691_ clknet_leaf_74_wb_clk_i _02808_ _01415_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08685__B team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11392__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15642_ clknet_leaf_119_wb_clk_i _01782_ _00450_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12854_ net610 _06197_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_17_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _04292_ net646 _07193_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__or3_1
X_15573_ clknet_leaf_41_wb_clk_i _01713_ _00381_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12785_ _06070_ _06313_ _06388_ net422 vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__o31a_1
XFILLER_0_51_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14524_ net1148 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
XANTENNA__09797__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11736_ net345 net2513 net601 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08905__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10470__A1 _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14455_ net1173 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
X_11667_ _05440_ _05464_ _05992_ _05376_ _05356_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__o32a_1
XANTENNA__12427__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ _03300_ _03016_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10618_ team_02_WB.instance_to_wrap.top.pc\[29\] _06134_ vssd1 vssd1 vccd1 vccd1
+ _06135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14386_ net1122 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09612__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ net945 _07083_ _07086_ net605 vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__o211a_4
XANTENNA__08206__A team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16125_ clknet_leaf_48_wb_clk_i _02265_ _00933_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08966__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13337_ net1055 team_02_WB.instance_to_wrap.top.ru.state\[2\] vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_iready sky130_fd_sc_hd__and2b_1
XFILLER_0_109_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10222__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10549_ _06064_ _06065_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16056_ clknet_leaf_19_wb_clk_i _02196_ _00864_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13268_ _06556_ _06588_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15007_ net1233 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
XANTENNA__12162__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12219_ net2646 net268 net616 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13199_ net1022 _02953_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_88_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07760_ _03457_ _03475_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__xor2_4
XFILLER_0_37_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09679__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09143__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15909_ clknet_leaf_31_wb_clk_i _02049_ _00717_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_07691_ _03372_ _03405_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__xnor2_1
X_16889_ net1433 vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__buf_2
X_09430_ net968 _04946_ _04497_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_133_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09361_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\] net746 _04867_ _04870_
+ _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_34_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08312_ _03997_ _04018_ _03999_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09292_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\] net818 net907 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\]
+ _04806_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09851__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12845__B _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _03932_ _03959_ _03929_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__a21o_2
XFILLER_0_16_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09500__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 _07069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12337__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout229_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08174_ _03892_ _03889_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09603__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08957__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13957__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12861__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1040_A _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1138_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__08709__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XANTENNA__12072__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput185 net185 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput196 net196 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XFILLER_0_100_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09382__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07958_ _03657_ _03678_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09134__A2 _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07889_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03609_ _03610_ vssd1 vssd1
+ vccd1 vccd1 _03612_ sky130_fd_sc_hd__or3_1
XFILLER_0_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\] net746 _05143_ _05144_
+ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09559_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\] net910 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\]
+ _05075_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ net360 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\] net443 vssd1
+ vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__mux2_1
XANTENNA__13208__A1_N net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09842__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16209__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11521_ net1635 net330 net643 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12247__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10556__A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08671__D team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11452_ _05468_ _05926_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__nor2_1
X_14240_ net1158 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10403_ net508 _05603_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14171_ net1157 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
X_11383_ _06014_ _06881_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15233__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10334_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\] net828 net804 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\]
+ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__a221o_1
X_13122_ _07471_ _07472_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__and2b_1
XANTENNA_input61_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13053_ net230 _02833_ _06526_ net234 vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__o2bb2a_1
X_10265_ net609 vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12004_ net352 net2624 net480 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
XANTENNA__09373__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ _05706_ _05709_ _05710_ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nor4_2
XANTENNA__15383__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16812_ net1356 vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout390 net391 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09125__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16743_ net1288 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
X_13955_ net1236 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12906_ _07367_ _07425_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__nand2_1
X_16674_ clknet_leaf_73_wb_clk_i _02791_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13209__B2 _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10140__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ net1257 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
XANTENNA__08884__B2 team_02_WB.instance_to_wrap.ramload\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_92_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15625_ clknet_leaf_104_wb_clk_i _01765_ _00433_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12837_ _04714_ _06143_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15556_ clknet_leaf_4_wb_clk_i _01696_ _00364_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12768_ _07277_ _07280_ _07281_ _07291_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__o22a_1
XANTENNA__09833__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14507_ net1200 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12157__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ net294 net2320 net602 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15487_ clknet_leaf_86_wb_clk_i _01627_ _00295_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12699_ _07051_ net2603 net433 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14438_ net1082 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput43 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11996__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput54 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
Xmax_cap502 net503 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_1
XFILLER_0_12_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput65 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap513 _05488_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_2
Xhold805 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ net1207 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
Xhold816 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xinput76 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
Xinput87 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_1
Xhold827 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xinput98 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
Xmax_cap535 net536 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16108_ clknet_leaf_10_wb_clk_i _02248_ _00916_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold838 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13145__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16039_ clknet_leaf_32_wb_clk_i _02179_ _00847_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08930_ net1512 _04449_ _04433_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16866__1410 vssd1 vssd1 vccd1 vccd1 _16866__1410/HI net1410 sky130_fd_sc_hd__conb_1
XFILLER_0_58_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09364__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08861_ net164 net1038 net1034 net1618 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07812_ _03532_ _03533_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08792_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] _04330_ net650 team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__a22o_2
XANTENNA__12620__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15876__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09116__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] _03398_ _03432_ vssd1 vssd1
+ vccd1 vccd1 _03466_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11236__S net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07674_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] _03393_ _03394_ vssd1 vssd1
+ vccd1 vccd1 _03397_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_1586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09413_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\] net895 net939 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12856__A _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1088_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ net971 net634 net543 vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16822__1366 vssd1 vssd1 vccd1 vccd1 _16822__1366/HI net1366 sky130_fd_sc_hd__conb_1
XFILLER_0_117_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\] net844 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\]
+ _04791_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12067__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1255_A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08226_ _03905_ _03914_ _03927_ _03908_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08157_ _03872_ _03873_ _03874_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__or3_2
XFILLER_0_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07602__A2 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08088_ _03801_ _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout882_A _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16651__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__C1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\] net845 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\]
+ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__a221o_1
XANTENNA__09355__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12530__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13740_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] _03245_ vssd1 vssd1 vccd1
+ vccd1 _03247_ sky130_fd_sc_hd__and2_1
XANTENNA__10122__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ net947 _06458_ _06465_ net607 vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10673__B2 _05625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13671_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] _03201_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1 _03205_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_116_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10883_ _06392_ _06393_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15410_ clknet_leaf_5_wb_clk_i _01550_ _00218_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12622_ net1712 net302 net553 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16390_ clknet_leaf_89_wb_clk_i _02525_ _01198_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15341_ clknet_leaf_79_wb_clk_i _00009_ _00154_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12553_ net275 net1853 net442 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11504_ _06049_ _06055_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_136_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16181__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15272_ clknet_leaf_70_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[31\]
+ _00085_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_134_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ net280 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\] net558 vssd1
+ vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15749__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14223_ net1115 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ team_02_WB.instance_to_wrap.top.pc\[11\] _06258_ vssd1 vssd1 vccd1 vccd1
+ _06932_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11366_ net1907 net297 net641 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
X_14154_ net1168 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
XANTENNA__09594__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10317_ _05785_ _04419_ net551 vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__mux2_1
X_13105_ _07369_ _07370_ _07421_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a21oi_1
X_14085_ net1128 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
X_11297_ _05211_ net665 vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15899__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13036_ _06422_ net234 _02820_ net978 net1028 vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__o221a_1
X_10248_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\] net756 net752 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1130 net1134 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1141 net1143 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__clkbuf_4
X_10179_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a22o_1
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_4
XANTENNA__12440__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1163 net1171 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__buf_4
Xfanout1174 net1179 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__buf_4
XFILLER_0_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1185 net1188 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_2
Xfanout1196 net1197 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__clkbuf_4
X_14987_ net1222 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16726_ net1450 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_135_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13938_ net1218 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XANTENNA__10113__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16657_ clknet_leaf_101_wb_clk_i _02776_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13869_ net1231 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15608_ clknet_leaf_19_wb_clk_i _01748_ _00416_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09806__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16588_ clknet_leaf_96_wb_clk_i _02707_ _01381_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16524__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08592__C net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09050__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11613__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15539_ clknet_leaf_86_wb_clk_i _01679_ _00347_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\] net775 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08011_ _03681_ _03713_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__xor2_2
XFILLER_0_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12615__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold602 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold613 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold624 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09585__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold635 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold646 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold657 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\] net752 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09337__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08913_ net1488 _04438_ net930 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__mux2_1
X_09893_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\] net821 net817 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\]
+ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout296_A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1302 team_02_WB.instance_to_wrap.ramaddr\[26\] vssd1 vssd1 vccd1 vccd1 net2760
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12350__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ net151 net1037 net1033 net1554 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16054__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08775_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\] net682 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\]
+ _04401_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout463_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _03406_ _03438_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07657_ _03345_ _03347_ _03351_ _03361_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout728_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07588_ team_02_WB.instance_to_wrap.top.a1.state\[1\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_81_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09327_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\] net818 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08076__A2 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09258_ net970 _04774_ net544 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08209_ _03897_ _03922_ _03923_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a21o_2
XANTENNA__12525__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09189_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\] net734 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\]
+ _04705_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10834__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11220_ _05974_ net665 _06723_ net668 _06724_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__o221a_1
XANTENNA__09576__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08784__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ _04997_ _05946_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09119__B net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__B team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10102_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\] net788 net685 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__a22o_1
XANTENNA__09328__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ net1000 _06590_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_21_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14910_ net1192 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
X_10033_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\] net823 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__a22o_1
XANTENNA__12260__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15890_ clknet_leaf_3_wb_clk_i _02030_ _00698_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10343__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ net1133 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10894__A1 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13880__A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14772_ net1090 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XANTENNA__15421__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08974__A team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ net270 net2037 net479 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
XANTENNA__16547__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16511_ clknet_leaf_37_wb_clk_i _02645_ _01318_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13723_ _03300_ _03016_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__nand2_1
X_10935_ net408 _06448_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16442_ clknet_leaf_64_wb_clk_i net1480 _01250_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ net1464 _04161_ net852 vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__mux2_1
X_10866_ _06380_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ net346 net2181 net438 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16373_ clknet_leaf_41_wb_clk_i _02513_ _01181_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13585_ net1548 net962 _03139_ net1066 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_45_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10797_ _06296_ _06312_ net414 vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_45_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15324_ clknet_leaf_63_wb_clk_i _01467_ _00137_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12536_ net354 net2363 net448 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08913__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12943__B _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15255_ clknet_leaf_66_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[14\]
+ _00068_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_10_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12435__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ net338 net2490 net453 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__mux2_1
XANTENNA__13024__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14206_ net1189 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XANTENNA__09567__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11418_ _06010_ _06011_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__xnor2_2
X_15186_ net1255 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12398_ net326 net2438 net460 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08775__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14137_ net1140 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
X_11349_ _06745_ _06848_ net397 vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__mux2_1
XANTENNA__09319__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14068_ net1091 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
XANTENNA__16077__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16821__1365 vssd1 vssd1 vccd1 vccd1 _16821__1365/HI net1365 sky130_fd_sc_hd__conb_1
XANTENNA__15047__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ team_02_WB.instance_to_wrap.top.pc\[31\] _06130_ vssd1 vssd1 vccd1 vccd1
+ _07539_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12170__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10334__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08560_ team_02_WB.instance_to_wrap.top.a1.hexop\[3\] _04228_ _04226_ vssd1 vssd1
+ vccd1 vccd1 _04229_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_102_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16709_ net1268 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
X_08491_ team_02_WB.instance_to_wrap.top.a1.data\[11\] net959 _04187_ vssd1 vssd1
+ vccd1 vccd1 _04188_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13036__C1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09112_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\] net738 _04625_ _04627_
+ _04628_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_21_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12853__B _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09043_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\] net885 _04559_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12345__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout309_A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09558__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold421 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold432 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12968__A_N _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08766__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold454 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13965__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1120_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold476 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold487 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold498 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 _04526_ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09945_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\] net920 net799 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\]
+ _05446_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__a221o_1
Xfanout912 _04523_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout580_A _07214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 _04513_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11117__A2 _06618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout678_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net946 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_4
Xfanout956 _04261_ vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12080__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout967 _02957_ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_4
X_09876_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\] net762 net698 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__a22o_1
XANTENNA__15444__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout978 _04281_ vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_4
Xhold1110 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 _04431_ vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_2
Xhold1121 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ net1611 net1042 net993 team_02_WB.instance_to_wrap.ramaddr\[4\] vssd1 vssd1
+ vccd1 vccd1 _02598_ sky130_fd_sc_hd__a22o_1
XANTENNA__09730__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1143 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1165 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1176 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ net848 _04360_ _04364_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__and3_4
Xhold1198 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _03302_ net425 vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08689_ net1057 _04278_ _04315_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__or3_2
XFILLER_0_71_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13290__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ _06144_ _06236_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10548__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10651_ net790 net552 _06166_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12250__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13370_ net1055 team_02_WB.instance_to_wrap.top.ru.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _03014_ sky130_fd_sc_hd__and2b_1
X_10582_ _06097_ _06098_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ net291 net1866 net567 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__mux2_1
XANTENNA__12255__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10564__A _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11457__A1_N net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09549__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ net1203 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
X_12252_ net268 net1951 net574 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11203_ net999 _06707_ _06708_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__o21bai_1
X_12183_ net256 net2458 net578 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ net667 _06641_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_53_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11108__A2 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15942_ clknet_leaf_42_wb_clk_i _02082_ _00750_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11065_ net398 _06448_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09182__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\] net684 _05528_ _05529_
+ _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__a2111oi_4
XANTENNA__09721__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ clknet_leaf_121_wb_clk_i _02013_ _00681_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15937__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14824_ net1175 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ net1131 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11967_ net337 net2456 net588 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10095__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ net1240 _03225_ _03226_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_47_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10918_ _06429_ _06431_ net396 vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__mux2_2
XFILLER_0_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14686_ net1191 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11898_ net330 net2084 net487 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16425_ clknet_leaf_104_wb_clk_i _02560_ _01233_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13637_ net2702 net963 _03186_ net1067 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__o211a_1
X_10849_ _04609_ net662 _06364_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__a21o_2
XFILLER_0_73_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16356_ clknet_leaf_0_wb_clk_i _02496_ _01164_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09788__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13568_ net1047 net1049 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] _03103_
+ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_97_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15307_ clknet_leaf_58_wb_clk_i team_02_WB.EN_VAL_REG _00120_ vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.testpc.en_latched sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_93_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12519_ net288 net2506 net448 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12165__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16287_ clknet_leaf_111_wb_clk_i _02427_ _01095_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13499_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\] _03063_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.lcd_en sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15238_ clknet_leaf_70_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[29\]
+ _00051_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ net1241 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XANTENNA__15467__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09960__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07991_ _03693_ net255 _03683_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09730_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\] net925 net913 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10307__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09712__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09661_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\] net727 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\]
+ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a221o_1
XANTENNA__08920__B1 _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ net84 net1578 net957 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__mux2_1
X_09592_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\] net916 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\]
+ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12848__B _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08543_ net1607 net793 net653 _04188_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
XANTENNA__13272__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout259_A _06530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08474_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__nor2_2
XFILLER_0_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12864__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1168_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12075__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09026_ net943 _04505_ _04509_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_76_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout795_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold240 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 team_02_WB.instance_to_wrap.ramstore\[2\] vssd1 vssd1 vccd1 vccd1 net1720
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold273 team_02_WB.instance_to_wrap.ramload\[0\] vssd1 vssd1 vccd1 vccd1 net1731
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout962_A _03027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 _04384_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_8
Xfanout731 net733 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09928_ _05444_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__inv_2
Xfanout742 net745 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_8
Xfanout753 _04376_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_4
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09164__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout775 net777 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
XANTENNA__09703__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout786 net789 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_8
X_09859_ net970 _05375_ net543 vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__o21a_1
Xfanout797 _04542_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12870_ _04423_ _07328_ _05877_ _05836_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_119_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11821_ net300 net2707 net590 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
XANTENNA__10559__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540_ net1072 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
X_11752_ net285 net1914 net599 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10703_ _06219_ _06218_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__and2b_1
XANTENNA__09015__A_N net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14471_ net1112 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
XANTENNA__10993__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _05970_ _07160_ _07168_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ clknet_leaf_5_wb_clk_i _02350_ _01018_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16820__1364 vssd1 vssd1 vccd1 vccd1 _16820__1364/HI net1364 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_23_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _03030_ _02765_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input91_A wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10634_ team_02_WB.instance_to_wrap.top.pc\[25\] _06150_ vssd1 vssd1 vccd1 vccd1
+ _06151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16141_ clknet_leaf_33_wb_clk_i _02281_ _00949_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13353_ net1580 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[15\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_52_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10565_ net546 net386 _06081_ net390 vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12304_ net358 net1901 net569 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16072_ clknet_leaf_15_wb_clk_i _02212_ _00880_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13284_ net1500 net983 net964 _02991_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__a22o_1
X_10496_ _05380_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15023_ net1223 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12235_ net2072 net331 net618 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10001__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ net323 net1935 net464 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ _04456_ _06618_ _06625_ net608 vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__o211a_4
X_12097_ net2254 net318 net581 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15925_ clknet_leaf_43_wb_clk_i _02065_ _00733_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11048_ team_02_WB.instance_to_wrap.top.pc\[24\] _06267_ team_02_WB.instance_to_wrap.top.pc\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__a21oi_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ clknet_leaf_41_wb_clk_i _01996_ _00664_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14807_ net1174 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
XANTENNA__10469__A _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15787_ clknet_leaf_14_wb_clk_i _01927_ _00595_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12999_ team_02_WB.instance_to_wrap.top.pc\[17\] _06192_ _07518_ vssd1 vssd1 vccd1
+ vccd1 _07519_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_52_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10068__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14738_ net1122 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13006__A2 _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14669_ net1154 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16408_ clknet_leaf_65_wb_clk_i _02543_ _01216_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11017__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15060__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08190_ _03906_ _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08969__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16339_ clknet_leaf_54_wb_clk_i _02479_ _01147_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10240__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12623__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09394__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13190__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09217__B _04733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ _03601_ _03645_ _03696_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__or3b_1
XFILLER_0_103_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09146__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ _05216_ _05217_ _05223_ _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__nor4_2
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12859__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09644_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\] net896 net893 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\] net776 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\]
+ _05091_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout543_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10059__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08526_ _04213_ net1614 net850 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11195__A2_N net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08457_ _04158_ _04160_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout710_A _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11702__S net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15632__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _04084_ _04085_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11559__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10350_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\] net741 _05865_ _05866_
+ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a211o_1
XANTENNA__10231__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09009_ _04295_ net944 _04505_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__and3_4
XFILLER_0_130_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15782__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10281_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\] net912 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12533__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10842__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12020_ net277 net1937 net476 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__mux2_1
XANTENNA__09385__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09137__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout561 _07219_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout572 _07217_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_4
Xfanout583 net584 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_8
X_13971_ net1254 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
Xfanout594 net596 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15710_ clknet_leaf_114_wb_clk_i _01850_ _00518_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12922_ _04489_ _06244_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11495__A1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12692__A0 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16690_ clknet_leaf_74_wb_clk_i _02807_ _01414_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11495__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08685__C team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ clknet_leaf_18_wb_clk_i _01781_ _00449_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12853_ _05231_ _06194_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14984__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] _04333_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_17_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15572_ clknet_leaf_13_wb_clk_i _01712_ _00380_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12784_ _06918_ _06946_ _07307_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__nand3_1
XFILLER_0_51_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14523_ net1185 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
X_11735_ net351 net1817 net604 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14454_ net1138 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
X_11666_ net513 _05511_ _06011_ _07151_ _05469_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13405_ _03300_ _03016_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__nor2_1
X_10617_ net552 _06133_ _06126_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_52_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14385_ net1107 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11597_ team_02_WB.instance_to_wrap.top.pc\[3\] net973 _04347_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\]
+ _07085_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16124_ clknet_leaf_44_wb_clk_i _02264_ _00932_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13336_ team_02_WB.instance_to_wrap.Wen _03297_ team_02_WB.instance_to_wrap.wb.curr_state\[0\]
+ _03301_ net2715 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10548_ _05231_ net406 vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16055_ clknet_leaf_14_wb_clk_i _02195_ _00863_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13267_ net1706 net985 net966 _02982_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a22o_1
XANTENNA__12443__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ _05878_ _05880_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__or2_2
X_15006_ net1229 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
XANTENNA__09376__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ net2545 net261 net617 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__mux2_1
XANTENNA__09915__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ _02953_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_write_i
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11059__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ net248 net2711 net462 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09128__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15505__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ clknet_leaf_0_wb_clk_i _02048_ _00716_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_07690_ _03385_ _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__xnor2_2
X_16888_ net1432 vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__buf_2
XFILLER_0_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15839_ clknet_leaf_109_wb_clk_i _01979_ _00647_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14894__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09360_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\] net843 _04871_ _04873_
+ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a2111o_1
XANTENNA__15655__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ _03997_ _03999_ _04018_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09291_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\] net826 net822 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12618__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_126_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_13 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ net224 _03957_ _03941_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__a21o_1
XANTENNA_24 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13222__A2_N net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_59_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08173_ _03849_ _03858_ _03891_ _03846_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_127_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10213__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__A1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12861__B _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12353__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1033_A _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_105_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XANTENNA__13163__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XANTENNA__09906__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_A _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput186 net186 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
Xoutput197 net197 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XANTENNA__12910__A1 _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1200_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _03661_ _03673_ _03679_ _03659_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__o22a_1
XANTENNA__13466__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A _04374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07888_ _03609_ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\] net698 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout925_A _04513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09558_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\] net886 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08509_ net1046 _04199_ _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12528__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\] net764 net748 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11520_ net945 _07007_ _07012_ net605 vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__o211a_2
XFILLER_0_0_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10556__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire236 _07326_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11451_ net656 _06942_ _06946_ net666 _06945_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10402_ net508 _05603_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10204__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14170_ net1184 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
X_11382_ _05378_ _05931_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__or2_1
XANTENNA__09070__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ net1026 _02891_ net1024 team_02_WB.instance_to_wrap.top.pc\[15\] vssd1 vssd1
+ vccd1 vccd1 _01496_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_103_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10333_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\] net909 net901 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10572__A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12263__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09358__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input54_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _07358_ _07359_ _07434_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__and3_1
X_10264_ _05770_ _05776_ _05780_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__nor3_2
XANTENNA__11165__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14979__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ net356 net2692 net478 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XANTENNA__12901__A1 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08030__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10195_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\] net890 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\]
+ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16811_ net1355 vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__buf_2
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout380 _06085_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_2
Xfanout391 _05856_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16742_ net1287 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_92_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13954_ net1213 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12905_ _07366_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__or2_1
X_16673_ clknet_leaf_73_wb_clk_i _02790_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13885_ net1251 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12417__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12836_ _04714_ _06143_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15624_ clknet_leaf_20_wb_clk_i _01764_ _00432_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12946__B _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08097__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15555_ clknet_leaf_125_wb_clk_i _01695_ _00363_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12767_ _05558_ _05921_ _07282_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12438__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14506_ net1156 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11718_ net284 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\] net601 vssd1
+ vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15486_ clknet_leaf_112_wb_clk_i _01626_ _00294_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12698_ net338 net2354 net433 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14437_ net1126 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11649_ net373 _06980_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__or2_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09597__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput44 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16303__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput55 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_1
X_14368_ net1148 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09061__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput66 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_1
Xinput77 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap514 net516 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold806 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ clknet_leaf_14_wb_clk_i _02247_ _00915_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput88 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
X_13319_ _07183_ _02959_ team_02_WB.instance_to_wrap.top.pc\[0\] net1051 vssd1 vssd1
+ vccd1 vccd1 _03009_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold828 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold839 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xinput99 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12173__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14299_ net1157 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
X_16038_ clknet_leaf_43_wb_clk_i _02178_ _00846_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11297__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08860_ net165 net1038 net1033 net1692 vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a22o_1
X_07811_ _03532_ _03533_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08791_ _04419_ _04417_ net551 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07742_ _03431_ _03464_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07673_ _03393_ _03394_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1
+ vccd1 vccd1 _03396_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_133_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09412_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\] net887 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13605__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _04853_ _04856_ _04858_ _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__nor4_2
XANTENNA_fanout241_A _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12348__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09274_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\] net755 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08225_ _03905_ _03914_ _03927_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1150_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09588__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ _03873_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10198__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12083__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ _03778_ _03780_ _03802_ _03806_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nand4_2
XANTENNA__10392__A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14799__A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout875_A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09760__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net944 _04503_ _04505_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09512__B1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ _06461_ _06462_ _06464_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__or3_1
XFILLER_0_98_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08866__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13670_ _03201_ _03202_ _03203_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__or3_1
X_10882_ net417 _06388_ _06396_ net373 vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12621_ net1738 net293 net553 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12258__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15340_ clknet_leaf_79_wb_clk_i _00008_ _00153_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12552_ net291 net2118 net443 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16326__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09291__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11503_ _05918_ _05923_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13878__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15271_ clknet_leaf_59_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[30\]
+ _00084_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12483_ net268 net2113 net557 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14222_ net1096 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
X_11434_ net669 _06915_ _06927_ _06930_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_80_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09043__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14153_ net1111 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
X_11365_ net606 _06858_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__and3_4
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_4_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13104_ _07466_ _07517_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__xnor2_1
X_10316_ _05829_ _05831_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__and2_1
XANTENNA__13127__B2 _07337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14084_ net1126 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11296_ net657 _06355_ _06797_ net418 vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13035_ _07439_ _02819_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10247_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\] net768 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1120 net1125 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09751__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1131 net1134 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1142 net1143 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__buf_4
XFILLER_0_94_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10178_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] net792 net652 _05694_
+ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a22oi_4
Xfanout1153 net1162 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_2
Xfanout1164 net1171 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_2
Xfanout1175 net1179 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1186 net1188 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_4
Xfanout1197 net1198 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14986_ net1245 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
XANTENNA__09503__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16725_ net1280 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
X_13937_ net1219 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13868_ net1233 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16656_ clknet_leaf_101_wb_clk_i _02775_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12819_ _07340_ _07341_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__nor2_1
X_15607_ clknet_leaf_116_wb_clk_i _01747_ _00415_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12168__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13799_ net1552 _03284_ net960 vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_100_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10477__A _05440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16587_ clknet_leaf_95_wb_clk_i _02706_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.lcd_rs
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09050__B _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15538_ clknet_leaf_11_wb_clk_i _01678_ _00346_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09282__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15469_ clknet_leaf_23_wb_clk_i _01609_ _00277_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08010_ _03726_ _03727_ _03731_ _03719_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__o31ai_2
XANTENNA__11800__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09034__A2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold603 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold614 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold625 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold658 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15843__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09961_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\] net704 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__a22o_1
XANTENNA__09990__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold669 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08912_ net1045 _04200_ _04211_ net1008 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__a32o_1
XFILLER_0_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09892_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\] net910 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a22o_1
XANTENNA__12631__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13207__A1_N _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08843_ net152 net1039 net1035 net1523 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1303 team_02_WB.instance_to_wrap.ramload\[23\] vssd1 vssd1 vccd1 vccd1 net2761
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15993__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08774_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] _04296_ _04302_ net931
+ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__and4_1
XFILLER_0_135_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ _03413_ _03446_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12867__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout456_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1198_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ _03345_ _03361_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16349__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_74_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12078__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07587_ _03311_ _03312_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_81_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09326_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\] net895 net939 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09273__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16499__CLK clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ _04764_ _04773_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nor2_4
XANTENNA__12806__S _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08208_ _03897_ _03922_ _03923_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_1390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\] net746 net843 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10834__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08139_ _03849_ _03855_ _03857_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13109__B2 _07337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11150_ net1899 net281 net641 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
XANTENNA__09981__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10101_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\] net753 net693 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__a22o_1
XANTENNA__08023__C team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12541__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ _06172_ net655 net495 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] net497
+ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14322__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _05542_ _05544_ _05546_ _05548_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__or4_1
X_14840_ net1196 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771_ net1169 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11983_ net261 net2482 net479 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13722_ _03016_ net950 _03235_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__and3_1
X_16510_ clknet_leaf_7_wb_clk_i _02644_ _01317_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10934_ _06345_ _06447_ net372 vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16441_ clknet_leaf_64_wb_clk_i net1640 _01249_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dfrtp_1
X_13653_ net1476 _04163_ net851 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__mux2_1
X_10865_ net368 _06041_ _06379_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15716__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12604_ net351 net1854 net440 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16372_ clknet_leaf_15_wb_clk_i _02512_ _01180_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13584_ team_02_WB.instance_to_wrap.top.a1.row2\[16\] _03124_ _03129_ _03131_ _03138_
+ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_67_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10796_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15323_ clknet_leaf_63_wb_clk_i _01466_ _00136_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12535_ net357 net2256 net446 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11071__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11620__S net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13401__A team_02_WB.instance_to_wrap.ramload\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15254_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[13\]
+ _00067_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12466_ net331 net2019 net452 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__mux2_1
X_14205_ net1085 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11417_ net2541 net315 net642 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15185_ net1255 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
X_12397_ net323 net2145 net460 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10031__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14136_ net1193 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11348_ _06793_ _06847_ net371 vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__mux2_1
X_14067_ net1165 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
XANTENNA__12451__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14232__A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ net670 _06768_ _06781_ net838 _06780_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__o221a_2
XFILLER_0_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09724__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ _07446_ _07537_ _07444_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13193__A1_N net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13284__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14969_ net1249 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16708_ net1267 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_72_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08490_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[11\] _04177_ vssd1 vssd1 vccd1
+ vccd1 _04187_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16639_ clknet_leaf_102_wb_clk_i _02758_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09255__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\] net782 net742 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12626__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09042_ net943 _04528_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__nor2_4
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold400 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\] vssd1
+ vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold422 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10022__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold455 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10573__A1 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold466 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold477 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16021__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout902 _04525_ vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_6
XFILLER_0_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold488 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\] net811 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\]
+ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout913 _04523_ vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12361__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold499 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1113_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout924 _04513_ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09715__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout935 _02960_ vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout946 _04456_ vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_2
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 _04261_ vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_2
X_09875_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\] net750 net734 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__a22o_1
Xfanout968 _04496_ vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_4
Xhold1100 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout573_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout979 _04281_ vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_2
Xhold1111 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ net1732 net1042 net990 net1694 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1133 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16171__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1166 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ _04359_ _04360_ _04361_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_87_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1177 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1188 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08794__B _04422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15739__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10089__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11705__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _03400_ _03428_ _03429_ _03430_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_68_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ net1058 _04315_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__or3b_1
XFILLER_0_75_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09494__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07639_ team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] _03335_ _03336_ _03361_ vssd1
+ vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11006__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ _04494_ _06166_ _06126_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_14_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15889__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09246__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11589__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\] net723 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11053__A2 _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12536__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10581_ _04886_ net405 vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_131_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11440__S net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10261__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ net276 net2252 net565 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12251_ net261 net2665 net574 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11202_ _06184_ net654 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] net496
+ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__a221o_1
XANTENNA__10013__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09954__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12182_ net250 net2009 net577 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11133_ net374 _06311_ _06342_ net378 _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__o221a_1
XANTENNA__11676__A _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12271__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__A _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15941_ clknet_leaf_34_wb_clk_i _02081_ _00749_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11064_ net668 _06573_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07592__C team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13891__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10015_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\] net741 _05530_ _05531_
+ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_30_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ clknet_leaf_107_wb_clk_i _02012_ _00680_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08985__A team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14823_ net1101 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13266__B1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14754_ net1207 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
X_11966_ _07013_ net2140 net587 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09485__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\]
+ _03222_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__and3_1
X_10917_ net389 _06286_ _06430_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_47_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14685_ net1083 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11897_ net334 net1917 net487 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16424_ clknet_leaf_67_wb_clk_i _02559_ _01232_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13636_ _03023_ _03183_ _03185_ _03164_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__or4b_1
X_10848_ net673 _06283_ _06284_ net672 _06363_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__a221o_1
XANTENNA__09237__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16355_ clknet_leaf_127_wb_clk_i _02495_ _01163_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13567_ net1047 _03103_ _03104_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__and3_1
XANTENNA__12446__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10779_ _06294_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15306_ clknet_leaf_71_wb_clk_i _01450_ _00119_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10252__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12518_ net278 net2401 net446 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__mux2_1
X_16286_ clknet_leaf_113_wb_clk_i _02426_ _01094_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13498_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\] _03019_ _03062_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] vssd1 vssd1 vccd1 vccd1 _03063_
+ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_93_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15237_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[28\]
+ _00050_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[28\]
+ sky130_fd_sc_hd__dfrtp_2
X_12449_ net262 net1760 net451 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap636_A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10004__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09945__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15168_ net1242 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ net1112 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
XANTENNA__12181__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07990_ _03683_ _03693_ _03703_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__nand3_2
X_15099_ net1098 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16194__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09660_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\] net779 net747 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08611_ net85 team_02_WB.START_ADDR_VAL_REG\[21\] net954 vssd1 vssd1 vccd1 vccd1
+ _02649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13257__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09591_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\] net880 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08542_ team_02_WB.instance_to_wrap.top.a1.state\[2\] net794 vssd1 vssd1 vccd1 vccd1
+ _04224_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13025__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08473_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ team_02_WB.instance_to_wrap.top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_63_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09228__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12864__B _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12356__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09025_ _04504_ _04516_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__nor2_4
XFILLER_0_5_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13976__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1230_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08739__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15411__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold230 team_02_WB.instance_to_wrap.ramload\[11\] vssd1 vssd1 vccd1 vccd1 net1688
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13085__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold241 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09400__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold252 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold263 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 net133 vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12091__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 team_02_WB.instance_to_wrap.top.a1.row2\[11\] vssd1 vssd1 vccd1 vccd1 net1743
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold296 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 _04386_ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_8
Xfanout721 _04384_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_4
Xfanout732 net733 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09927_ _04326_ _05441_ _05443_ net652 vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a22oi_4
Xfanout743 net745 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout754 _04375_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__buf_6
XANTENNA_fanout955_A _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 _04373_ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_4
Xfanout776 net777 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_6
Xfanout787 net789 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_4
XFILLER_0_99_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09858_ _05370_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__nor2_2
XANTENNA__10849__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout798 _04542_ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_4
X_08809_ net1788 net1042 net992 team_02_WB.instance_to_wrap.ramaddr\[22\] vssd1 vssd1
+ vccd1 vccd1 _02616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09789_ _05298_ _05299_ _05301_ _05305_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11259__C1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11820_ net292 net2186 net589 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09467__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10559__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11751_ net275 net1955 net597 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11274__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13650__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10702_ team_02_WB.instance_to_wrap.top.pc\[18\] _06188_ vssd1 vssd1 vccd1 vccd1
+ _06219_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14470_ net1089 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _04842_ _04861_ _05971_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__o211a_1
XANTENNA__09219__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13421_ net1065 _03031_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10633_ _06128_ _06149_ _04490_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__a21oi_4
XANTENNA__16067__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12266__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16140_ clknet_leaf_21_wb_clk_i _02280_ _00948_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10234__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13352_ net2098 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[14\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_106_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input84_A wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10564_ _04589_ net386 vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12303_ net341 net2073 net572 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__mux2_1
X_16071_ clknet_leaf_29_wb_clk_i _02211_ _00879_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13283_ team_02_WB.instance_to_wrap.top.pc\[18\] net1052 _06759_ net934 vssd1 vssd1
+ vccd1 vccd1 _02991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10495_ _05993_ _06010_ _05992_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__a21o_1
X_15022_ net1218 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
XANTENNA__07884__A team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12234_ net2717 net335 net618 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12165_ net319 net2121 net462 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net1000 _06623_ _06624_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_9_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12096_ net2104 net313 net581 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XANTENNA__13487__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13240__A_N _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11047_ _06150_ net655 net495 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] net497
+ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15924_ clknet_leaf_11_wb_clk_i _02064_ _00732_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08919__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12949__B _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15855_ clknet_leaf_38_wb_clk_i _01995_ _00663_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14806_ net1090 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
XANTENNA__09458__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15786_ clknet_leaf_0_wb_clk_i _01926_ _00594_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12998_ _07466_ _07517_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14737_ net1106 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11949_ net261 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\] net586 vssd1
+ vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14668_ net1071 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16407_ clknet_leaf_66_wb_clk_i _02542_ _01215_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12176__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08418__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ team_02_WB.instance_to_wrap.top.a1.row1\[11\] _03110_ _03121_ team_02_WB.instance_to_wrap.top.a1.row1\[115\]
+ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__a22o_1
X_14599_ net1112 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16338_ clknet_leaf_3_wb_clk_i _02478_ _01146_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09091__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16269_ clknet_leaf_24_wb_clk_i _02409_ _01077_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09918__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13190__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07973_ _03647_ _03674_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13478__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09712_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\] net676 _05213_ _05226_
+ _05228_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_103_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09697__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\] net916 _05157_ _05159_
+ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout271_A _06626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout369_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09574_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\] net752 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09449__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08525_ net1046 _04211_ _04212_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1180_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08456_ _04149_ _04150_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11008__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12086__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08387_ _04094_ _04096_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout703_A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire429 _05623_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09082__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09621__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15927__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09008_ _04295_ _04501_ _04507_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__and3_4
XFILLER_0_131_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\] net896 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10842__B net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13469__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
Xfanout562 _07219_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_4
Xfanout573 net576 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_6
X_13970_ net1251 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
Xfanout584 _07209_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_8
XFILLER_0_57_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _07352_ _07440_ _07350_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08685__D team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15640_ clknet_leaf_19_wb_clk_i _01780_ _00448_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12852_ _05231_ _06194_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_17_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ net345 net2455 net593 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__mux2_1
X_12783_ _06536_ _06569_ net416 vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__a21o_1
X_15571_ clknet_leaf_55_wb_clk_i _01711_ _00379_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15457__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11734_ net362 net1999 net602 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__mux2_1
X_14522_ net1180 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14453_ net1214 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
X_11665_ net513 _05511_ net512 _05556_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10207__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10616_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] net995 _06127_ vssd1
+ vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__a21oi_1
X_13404_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _03016_
+ sky130_fd_sc_hd__nand3_1
XANTENNA__09073__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14384_ net1100 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
X_11596_ net998 _07084_ net946 vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09612__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13335_ _03296_ team_02_WB.instance_to_wrap.Ren team_02_WB.instance_to_wrap.wb.curr_state\[0\]
+ _03301_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _00014_
+ sky130_fd_sc_hd__a32o_1
X_16123_ clknet_leaf_127_wb_clk_i _02263_ _00931_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10547_ _05271_ net384 vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__nor2_1
XANTENNA__08820__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16054_ clknet_leaf_45_wb_clk_i _02194_ _00862_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13266_ net935 _02962_ _02981_ net1054 team_02_WB.instance_to_wrap.top.pc\[26\] vssd1
+ vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a32o_1
X_10478_ net548 net403 vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15005_ net1234 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
X_12217_ net1925 net264 net617 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__mux2_1
X_13197_ team_02_WB.instance_to_wrap.top.d_ready _03308_ _04286_ _04289_ vssd1 vssd1
+ vccd1 vccd1 _02953_ sky130_fd_sc_hd__or4_2
XFILLER_0_27_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12148_ net253 net2572 net464 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net1733 net240 net581 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XANTENNA__14240__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ clknet_leaf_125_wb_clk_i _02047_ _00715_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16887_ net1431 vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__buf_2
XFILLER_0_56_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15838_ clknet_leaf_118_wb_clk_i _01978_ _00646_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire504_A _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15769_ clknet_leaf_16_wb_clk_i _01909_ _00577_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11803__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08310_ _04009_ _04023_ _04017_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_129_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15071__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09290_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\] net926 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09851__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08241_ _03949_ _03957_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_14 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_36 _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ _03806_ _03840_ _03847_ _03859_ _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a41o_1
XFILLER_0_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09603__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12634__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08811__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_28_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_11_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
Xoutput187 net187 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput198 net198 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout486_A _07198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _03678_ _03657_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__and2b_1
XANTENNA__08878__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] net316 _03597_ vssd1 vssd1
+ vccd1 vccd1 _03610_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\] net786 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09557_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\] net918 _05072_ _05073_
+ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout820_A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_A _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11713__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[7\] net980 vssd1 vssd1 vccd1
+ vccd1 _04200_ sky130_fd_sc_hd__or2_1
X_09488_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\] net845 _05002_ _05004_
+ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09842__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08439_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04125_ vssd1 vssd1 vccd1
+ vccd1 _04144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11450_ net416 _06504_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__or2_1
XANTENNA__09055__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10401_ _05648_ _05917_ _05647_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07605__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08802__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ net795 _06874_ _06876_ net656 _06879_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12544__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10853__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _06834_ net233 _02890_ net978 _02888_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__o221a_1
X_10332_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\] net816 net812 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\]
+ _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__a221o_1
XANTENNA__16105__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13051_ _07532_ _02832_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__xnor2_1
X_10263_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\] net772 _05764_ _05778_
+ _05779_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__a2111o_1
X_12002_ net342 net2731 net481 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
XANTENNA__12901__A2 _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08030__B2 _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\] net855 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__a22o_1
X_16810_ net1354 vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__buf_2
XFILLER_0_79_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 net371 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_2
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_4
X_16741_ net1286 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
Xfanout392 net401 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_4
X_13953_ net1236 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13159__A_N net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12904_ _05103_ _06188_ _07423_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__a21o_1
X_16672_ clknet_leaf_73_wb_clk_i _02789_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ net1238 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
XANTENNA__10140__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15623_ clknet_leaf_27_wb_clk_i _01763_ _00431_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12835_ net542 _06139_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15554_ clknet_leaf_123_wb_clk_i _01694_ _00362_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09294__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12766_ _05467_ _05514_ _05879_ _07289_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13090__A1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09833__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14505_ net1101 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
X_11717_ net275 net2139 net601 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
X_15485_ clknet_leaf_51_wb_clk_i _01625_ _00293_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12697_ net331 net2472 net432 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09046__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11648_ net409 _07053_ _07132_ _07133_ net378 vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__a221o_1
X_14436_ net1130 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12962__B _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput34 gpio_in[19] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
XFILLER_0_80_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput45 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
X_14367_ net1169 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12454__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11579_ net945 _07064_ _07068_ net605 vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__o211a_4
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput56 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
XFILLER_0_52_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold807 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
Xinput67 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
X_16106_ clknet_leaf_129_wb_clk_i _02246_ _00914_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput78 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__buf_1
X_13318_ net1633 net986 net967 _03008_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput89 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
Xhold818 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ net1180 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
X_16037_ clknet_leaf_33_wb_clk_i _02177_ _00845_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13249_ team_02_WB.instance_to_wrap.top.pc\[31\] net1054 _06124_ _02968_ _02969_
+ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a221o_1
XANTENNA__11156__A1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07810_ _03483_ _03529_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__xnor2_4
X_08790_ net1057 net650 _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__a21o_1
XANTENNA__15622__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire621_A _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ _03461_ _03462_ _03436_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_74_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11459__A2 _06950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07672_ _03393_ _03394_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09411_ net614 vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_94_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12629__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__A _05715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09342_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\] net826 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\]
+ _04844_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09824__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09273_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\] net743 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16699__1266 vssd1 vssd1 vccd1 vccd1 _16699__1266/HI net1266 sky130_fd_sc_hd__conb_1
XFILLER_0_69_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout234_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ net225 _03937_ _03939_ _03931_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09037__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08155_ _03827_ net226 _03820_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12364__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_A _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10198__A2 _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1143_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08086_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10392__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13984__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11147__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout770_A _04371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__B2 _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout868_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ team_02_WB.instance_to_wrap.top.a1.instruction\[21\] net951 team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__and3b_2
XFILLER_0_138_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10370__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07939_ _03601_ _03639_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10950_ _06238_ _06463_ net975 vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__and3b_1
XFILLER_0_39_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10122__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ net531 _05122_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__nand2_1
X_10881_ _06394_ _06395_ net393 vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__mux2_1
XANTENNA__12539__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input101_A wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12620_ net2442 net286 net555 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13072__B2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10567__B net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ net276 net2424 net442 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11502_ _05923_ _06005_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09028__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12482_ net260 net1988 net558 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__mux2_1
X_15270_ clknet_leaf_70_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[29\]
+ _00083_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11433_ net673 _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__nand2_1
X_14221_ net1141 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
XANTENNA__12274__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14152_ net1177 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11364_ _06197_ net654 _06837_ _06863_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10315_ _05829_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__nand2_2
XANTENNA__13894__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13103_ net1027 _02876_ net1024 team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1
+ vccd1 vccd1 _01499_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13127__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14083_ net1131 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11295_ _06579_ _06796_ net413 vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11138__A1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15645__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ _07353_ _07354_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__nand2_1
XANTENNA__08003__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10246_ net969 _05742_ _05761_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__o21a_1
XANTENNA__09200__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1110 net1116 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_2
Xfanout1121 net1122 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_4
XANTENNA__08554__A2 _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1132 net1133 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_4
X_10177_ _05668_ _05693_ net551 vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__mux2_1
Xfanout1143 net1144 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1154 net1162 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__buf_4
XANTENNA__08500__B net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1165 net1171 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__buf_4
Xfanout1176 net1179 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13221__A2_N net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1187 net1188 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_4
X_14985_ net1245 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
Xfanout1198 net1199 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__buf_4
X_16724_ net1279 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
X_13936_ net1200 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
XANTENNA__10113__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16655_ clknet_leaf_101_wb_clk_i _02774_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13867_ net1233 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
XANTENNA__12449__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15606_ clknet_leaf_48_wb_clk_i _01746_ _00414_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12818_ _04172_ _04180_ _03317_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09267__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16586_ clknet_leaf_93_wb_clk_i _02705_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ _03284_ _03285_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09806__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15537_ clknet_leaf_22_wb_clk_i _01677_ _00345_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12749_ _04906_ _04993_ _05038_ _05081_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15468_ clknet_leaf_20_wb_clk_i _01608_ _00276_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14419_ net1163 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16420__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12184__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15399_ clknet_leaf_29_wb_clk_i _01539_ _00207_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold604 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold615 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold626 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold637 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\] net764 net716 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\]
+ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a221o_1
Xhold659 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ net1542 _04437_ net930 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__mux2_1
X_09891_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\] net833 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\]
+ _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12877__A1 _07388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08842_ net153 net1040 net1036 net1585 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a22o_1
Xhold1304 team_02_WB.instance_to_wrap.ramaddr\[9\] vssd1 vssd1 vccd1 vccd1 net2762
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10352__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08773_ _04359_ _04364_ _04370_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07724_ _03413_ _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10104__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11301__B2 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09522__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ _03363_ _03368_ _03376_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12359__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_A _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11263__S net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A _07224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07586_ team_02_WB.instance_to_wrap.top.pad.count\[0\] _03310_ vssd1 vssd1 vccd1
+ vccd1 _03312_ sky130_fd_sc_hd__or2_1
XANTENNA__13054__A1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09258__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09325_ net532 vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1260_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ _04766_ _04768_ _04770_ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__or4_2
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08207_ _03911_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__and2_2
Xclkbuf_leaf_43_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12094__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09187_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\] net762 net698 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08138_ _03849_ _03855_ _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09430__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout985_A _02956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13109__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ _03788_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__or2_2
XFILLER_0_102_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10100_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\] net773 net757 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__a22o_1
XANTENNA__08023__D team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11080_ team_02_WB.instance_to_wrap.top.pc\[24\] _06267_ vssd1 vssd1 vccd1 vccd1
+ _06590_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10031_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\] net835 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\]
+ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10343__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ net1123 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ net266 net2749 net479 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__mux2_1
XANTENNA__09497__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13293__B2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13721_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _03235_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09432__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10933_ net542 _05901_ _06316_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12269__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ clknet_leaf_104_wb_clk_i _02575_ _01248_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09249__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ net368 _06047_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__nand2_1
X_13652_ net1469 _04165_ net851 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13889__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ net362 net2105 net440 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16371_ clknet_leaf_56_wb_clk_i _02511_ _01179_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16443__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10795_ _06303_ _06310_ net392 vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__mux2_1
X_13583_ _03132_ _03134_ _03137_ _03136_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__or4b_1
XANTENNA__08990__B team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11901__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15322_ clknet_leaf_64_wb_clk_i _01465_ _00135_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07887__A team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12534_ net341 net2149 net449 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15253_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[12\]
+ _00066_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12465_ net333 net1761 net452 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14204_ net1152 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11416_ net945 _06908_ _06913_ net605 vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__o211a_2
XANTENNA__09421__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12396_ net319 net1876 net458 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15184_ net1239 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ net1173 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11347_ _06308_ _06330_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__or2_1
XANTENNA__08775__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09607__A _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14066_ net1117 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
X_11278_ _05942_ _05980_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13017_ _07448_ _07536_ vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__or2_1
X_10229_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\] net857 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10334__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1 team_02_WB.instance_to_wrap.busy_o vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14968_ net1193 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16707_ net1445 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
X_13919_ net1200 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
XANTENNA__12179__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14899_ net1165 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16638_ clknet_leaf_102_wb_clk_i _02757_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13036__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16569_ clknet_leaf_94_wb_clk_i _02693_ _01376_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11811__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09110_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\] net774 net762 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\]
+ _04626_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_119_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09660__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09041_ _04554_ _04555_ _04556_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__or4_1
XFILLER_0_128_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09412__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold401 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold412 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold434 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12642__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15960__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold456 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold467 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold478 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09943_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\] net916 net896 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__a22o_1
Xhold489 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout903 _04525_ vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout914 _04518_ vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_6
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10670__B _05625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout925 _04513_ vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_4
Xfanout936 _02955_ vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout399_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout947 _04456_ vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
X_09874_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\] net686 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__a22o_1
XANTENNA__10325__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout958 net959 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_2
XANTENNA__16316__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1106_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout969 _04496_ vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_4
Xhold1101 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09191__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08825_ net1628 net1042 net990 team_02_WB.instance_to_wrap.ramaddr\[6\] vssd1 vssd1
+ vccd1 vccd1 _02600_ sky130_fd_sc_hd__a22o_1
Xhold1123 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1145 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _04359_ _04360_ _04364_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_87_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1178 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
X_07707_ _03364_ _03399_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12089__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ net1057 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _04316_ sky130_fd_sc_hd__nor2_1
XANTENNA__10398__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07638_ _03356_ _03359_ team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] _03329_ vssd1
+ vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07569_ net1069 vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout900_A _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11721__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09308_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\] net691 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10941__A1_N _04694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10580_ _04928_ net386 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09239_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\] net886 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12250_ net264 net1756 net574 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__mux2_1
XANTENNA__09403__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11201_ _06265_ _06706_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12181_ net253 net1824 net579 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__mux2_1
XANTENNA__12552__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ _06296_ _06638_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold990 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ net416 _06569_ _06572_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__a21o_1
X_15940_ clknet_leaf_4_wb_clk_i _02080_ _00748_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11513__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\] net772 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__a22o_1
XANTENNA__09182__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15871_ clknet_leaf_110_wb_clk_i _02011_ _00679_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14822_ net1072 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
XANTENNA__15164__A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13266__A1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14753_ net1209 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11965_ net333 net2637 net587 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\] _03222_ net1553 vssd1
+ vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10916_ net389 _06291_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_47_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14684_ net1146 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09890__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ net326 net2291 net486 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__mux2_1
XANTENNA__15833__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16423_ clknet_leaf_67_wb_clk_i _02558_ _01231_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13635_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] team_02_WB.instance_to_wrap.top.a1.row1\[101\]
+ _03184_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__and3_1
X_10847_ net668 _06344_ _06360_ net657 _06362_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_15_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16354_ clknet_leaf_122_wb_clk_i _02494_ _01162_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13206__A1_N _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13566_ _03290_ _03115_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__and3_1
X_10778_ _06291_ _06293_ net368 vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09642__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15305_ clknet_leaf_75_wb_clk_i _01449_ _00118_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12517_ net281 net2190 net447 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16285_ clknet_leaf_52_wb_clk_i _02425_ _01093_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15983__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13497_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15236_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[27\]
+ _00049_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[27\]
+ sky130_fd_sc_hd__dfrtp_2
X_12448_ net264 net1604 net451 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12970__B _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12462__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10771__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ net1244 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
X_12379_ net251 net1836 net461 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16339__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ net1082 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098_ net1098 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14049_ net1159 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10307__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11806__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ net86 net1509 net957 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
X_09590_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\] net827 net892 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\]
+ _05106_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09072__A _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08541_ _03291_ net794 _03319_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08472_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ team_02_WB.instance_to_wrap.top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__nor3b_2
XTAP_TAPCELL_ROW_63_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12637__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14418__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09633__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout314_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1056_A team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ _04519_ _04527_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 team_02_WB.instance_to_wrap.ramstore\[26\] vssd1 vssd1 vccd1 vccd1 net1678
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08739__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12372__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 net128 vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 team_02_WB.instance_to_wrap.top.a1.row2\[19\] vssd1 vssd1 vccd1 vccd1 net1700
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 team_02_WB.instance_to_wrap.ramaddr\[4\] vssd1 vssd1 vccd1 vccd1 net1722
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold275 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 team_02_WB.instance_to_wrap.ramstore\[14\] vssd1 vssd1 vccd1 vccd1 net1744
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout683_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout700 net701 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_6
Xhold297 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 _04386_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__buf_4
Xfanout722 _04383_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_6
XFILLER_0_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09926_ _04417_ _05442_ net552 vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__mux2_1
Xfanout733 _04381_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_8
Xfanout744 net745 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_8
Xfanout755 _04375_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09164__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout766 _04372_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_8
Xfanout777 _04369_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_4
X_09857_ _05359_ _05361_ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__or3_1
Xfanout788 net789 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_6
XFILLER_0_77_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout799 _04542_ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__buf_6
XFILLER_0_119_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11716__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ net1546 net1041 net990 team_02_WB.instance_to_wrap.ramaddr\[23\] vssd1 vssd1
+ vccd1 vccd1 _02617_ sky130_fd_sc_hd__a22o_1
X_09788_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\] net726 _05302_ _05304_
+ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15856__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08739_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_55_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ net288 net2338 net599 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__mux2_1
XANTENNA__09872__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10701_ team_02_WB.instance_to_wrap.top.pc\[17\] _06190_ _06217_ vssd1 vssd1 vccd1
+ vccd1 _06218_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12547__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11681_ _05982_ _07165_ _07166_ _06019_ _04862_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_42_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ team_02_WB.instance_to_wrap.top.lcd.currentState\[2\] team_02_WB.instance_to_wrap.top.lcd.nextState\[2\]
+ net962 vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__mux2_1
X_10632_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] net995 vssd1 vssd1 vccd1
+ vccd1 _06149_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13351_ net1713 net1016 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[13\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_91_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10563_ _04631_ net404 vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12302_ net337 net2550 net572 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__mux2_1
X_16070_ clknet_leaf_44_wb_clk_i _02210_ _00878_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input77_A wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13282_ net1496 net985 net966 _02990_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10494_ _05992_ _05993_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and2b_2
XFILLER_0_122_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15021_ net1204 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
XANTENNA__12282__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ net2155 net327 net618 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12164_ net315 net2394 net462 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15386__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ net975 _06620_ _06621_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16631__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12095_ net1949 net307 net581 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11046_ _06151_ _06152_ _06233_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__o21ai_1
X_15923_ clknet_leaf_85_wb_clk_i _02063_ _00731_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15854_ clknet_leaf_8_wb_clk_i _01994_ _00662_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10170__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14805_ net1187 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15785_ clknet_leaf_118_wb_clk_i _01925_ _00593_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12997_ _07467_ _07516_ _07469_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__a21oi_1
X_14736_ net1077 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11948_ net265 net2385 net586 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ net1151 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XANTENNA__12457__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11879_ net256 net1845 net488 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16406_ clknet_leaf_66_wb_clk_i _02541_ _01214_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13618_ team_02_WB.instance_to_wrap.top.a1.row2\[11\] _03122_ _03124_ team_02_WB.instance_to_wrap.top.a1.row2\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__a22o_1
XANTENNA__09615__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14598_ net1073 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
XANTENNA__10225__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08969__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16337_ clknet_leaf_22_wb_clk_i _02477_ _01145_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13549_ net1049 _03290_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__nor2_1
XANTENNA__09091__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16161__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16268_ clknet_leaf_25_wb_clk_i _02408_ _01076_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13175__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15219_ clknet_leaf_63_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[10\]
+ _00032_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15729__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12192__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16199_ clknet_leaf_29_wb_clk_i _02339_ _01007_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09394__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07972_ _03684_ _03693_ _03680_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__a21o_1
XANTENNA__13478__A1 team_02_WB.START_ADDR_VAL_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\] net725 net681 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\]
+ _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a221o_1
XANTENNA__09146__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09642_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\] net870 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\]
+ _05158_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a221o_1
XANTENNA__10161__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09573_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\] net788 net845 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout264_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08524_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[3\] net980 vssd1 vssd1 vccd1
+ vccd1 _04212_ sky130_fd_sc_hd__or2_2
XANTENNA__09854__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13650__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08455_ _04149_ _04152_ _04150_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12367__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_A _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1173_A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11271__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15259__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08386_ _04087_ _04089_ _04093_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o31a_1
XFILLER_0_50_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout898_A _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ _04313_ net943 _04507_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16654__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09385__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09137__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout552 _04356_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_4
X_09909_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\] net788 _05423_ _05425_
+ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__a211o_1
Xfanout563 _07219_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_6
Xfanout574 net576 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_8
Xfanout585 _07202_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_8
X_12920_ _07353_ _07439_ _07354_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__a21bo_1
Xfanout596 _07192_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12851_ net522 _06192_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__16034__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11802_ net348 net2663 net595 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ clknet_leaf_6_wb_clk_i _01710_ _00378_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09845__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12782_ _07295_ _07302_ _07303_ _07305_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14521_ net1140 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11733_ net354 net2635 net602 vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__mux2_1
XANTENNA__12277__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10586__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14058__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16184__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14452_ net1075 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
X_11664_ _05919_ _07146_ _07147_ _07149_ _07140_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__a41o_1
XFILLER_0_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ net2675 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\] vssd1 vssd1 vccd1
+ vccd1 _03015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10615_ _03293_ _06130_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14383_ net1111 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11595_ team_02_WB.instance_to_wrap.top.pc\[3\] team_02_WB.instance_to_wrap.top.pc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16122_ clknet_leaf_120_wb_clk_i _02262_ _00930_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13334_ _04243_ _04247_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10546_ _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08820__B2 team_02_WB.instance_to_wrap.ramaddr\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16053_ clknet_leaf_41_wb_clk_i _02193_ _00861_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13265_ _06523_ _02961_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10477_ _05440_ _05464_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__nand2_1
X_15004_ net1229 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12216_ net1887 net258 net617 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09376__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13196_ net1055 team_02_WB.instance_to_wrap.top.ru.state\[6\] team_02_WB.instance_to_wrap.Wen
+ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a21o_4
X_16789__1333 vssd1 vssd1 vccd1 vccd1 _16789__1333/HI net1333 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12147_ net238 net2405 net462 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09128__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ net2677 net246 net583 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11029_ net419 _06536_ _06539_ net376 vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__a22o_1
X_15906_ clknet_leaf_123_wb_clk_i _02046_ _00714_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16886_ net1430 vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__buf_2
XFILLER_0_56_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15837_ clknet_leaf_50_wb_clk_i _01977_ _00645_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15768_ clknet_leaf_19_wb_clk_i _01908_ _00576_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09836__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16527__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09300__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14719_ net1189 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
XANTENNA__12187__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15699_ clknet_leaf_55_wb_clk_i _01839_ _00507_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08240_ _03910_ _03942_ _03954_ _03955_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__or4_2
XFILLER_0_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_15 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_26 _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08171_ _03778_ _03842_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08811__A1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_112_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09367__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput188 net188 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XANTENNA__12650__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14431__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput199 net199 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1019_A _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07955_ _03652_ _03655_ _03670_ _03672_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_103_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout381_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10134__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ net316 _03597_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1
+ vccd1 vccd1 _03609_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09625_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\] net780 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09556_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\] net914 net817 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\]
+ _05062_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09827__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08507_ team_02_WB.instance_to_wrap.top.a1.data\[7\] net958 vssd1 vssd1 vccd1 vccd1
+ _04199_ sky130_fd_sc_hd__or2_1
XANTENNA__12097__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout813_A _04521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09487_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\] net744 net708 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\]
+ _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08438_ net1850 net1005 net981 _04143_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08369_ _04073_ _04079_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ _05912_ _05915_ _05691_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_104_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11380_ _06877_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10331_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\] net835 net905 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13050_ _07452_ _07453_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__and2b_1
X_10262_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\] net764 net712 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__a22o_1
XANTENNA__09358__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12001_ net339 net1878 net480 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08030__A2 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\] net809 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\]
+ _05697_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__a221o_1
XANTENNA__12560__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10373__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout360 net363 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13311__B1 _07064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16740_ net1285 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
Xfanout382 _06084_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_2
Xfanout393 net395 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_4
X_13952_ net1236 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
XANTENNA__10125__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _07370_ _07422_ _07368_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__a21oi_1
X_16671_ clknet_leaf_73_wb_clk_i _02788_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09530__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13883_ net1259 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
XANTENNA__11904__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15622_ clknet_leaf_42_wb_clk_i _01762_ _00430_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12834_ _04631_ _06134_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15553_ clknet_leaf_124_wb_clk_i _01693_ _00361_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15574__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08097__A2 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12765_ _04567_ _06116_ _07283_ _07288_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__or4_1
XFILLER_0_70_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14504_ net1177 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11716_ net290 net2245 net601 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
X_15484_ clknet_leaf_49_wb_clk_i _01624_ _00292_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12696_ net334 net2327 net432 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14435_ net1131 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11647_ net389 _06285_ _07128_ net396 vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__o31a_1
XFILLER_0_68_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09597__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput35 gpio_in[20] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
X_14366_ net1190 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput46 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11578_ team_02_WB.instance_to_wrap.top.pc\[4\] net973 _04347_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\]
+ _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput57 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput68 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16105_ clknet_leaf_119_wb_clk_i _02245_ _00913_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap505 net506 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_2
X_13317_ team_02_WB.instance_to_wrap.top.pc\[1\] net1051 _07122_ net933 vssd1 vssd1
+ vccd1 vccd1 _03008_ sky130_fd_sc_hd__a22o_2
Xhold808 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10529_ net505 net385 vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__and2_1
Xinput79 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_1
Xmax_cap527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold819 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14297_ net1138 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
X_16036_ clknet_leaf_1_wb_clk_i _02176_ _00844_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13248_ _06124_ _02959_ _02966_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__nor3_1
XFILLER_0_122_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12470__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ _07048_ net235 _02937_ _04281_ _02939_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__o221a_1
XANTENNA__10364__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09345__A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11086__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07740_ _03461_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10116__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11313__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire614_A _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07671_ _03356_ _03359_ _03388_ _03358_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__o22ai_4
X_16869_ net1413 vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__buf_2
XANTENNA__15082__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ _04915_ _04921_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__nor3_2
XANTENNA__11814__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09809__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\] net907 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\]
+ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09272_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\] net787 net707 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\]
+ _04788_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_115_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08223_ _03931_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12645__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08154_ _03820_ _03827_ net226 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__and3_1
XANTENNA__09588__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08424__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08085_ _03777_ _03804_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_70_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout596_A _07192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1244_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15447__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout763_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\] _04502_ vssd1 vssd1
+ vccd1 vccd1 _04504_ sky130_fd_sc_hd__or2_1
X_07938_ _03652_ _03655_ _03657_ _03659_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__o211ai_2
XANTENNA__10602__A1_N net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09512__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07869_ _03523_ _03562_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11724__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ _05103_ _05122_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10880_ _06092_ _06096_ net371 vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09539_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\] net726 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__a22o_1
XANTENNA__12766__D _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13072__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16788__1332 vssd1 vssd1 vccd1 vccd1 _16788__1332/HI net1332 sky130_fd_sc_hd__conb_1
XFILLER_0_94_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12550_ net282 net1860 net444 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ net2353 net335 net643 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ net266 net2579 net558 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__mux2_1
XANTENNA__12555__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14220_ net1071 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09579__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ _06011_ _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14151_ net1105 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
XANTENNA__16222__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11363_ net973 _06209_ _06859_ _06862_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13102_ net978 _07423_ _02874_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__o31a_1
X_10314_ net396 net498 vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__nand2_1
X_14082_ net1207 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
X_11294_ net407 _06690_ _06795_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13033_ _07448_ _07536_ _02817_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a21o_1
X_10245_ net969 _05742_ _05761_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12290__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10346__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1100 net1103 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__buf_2
Xfanout1111 net1112 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_4
XFILLER_0_24_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10176_ team_02_WB.instance_to_wrap.top.a1.instruction\[16\] net650 _05692_ vssd1
+ vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__a21o_1
Xfanout1122 net1124 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_4
XANTENNA__09751__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10897__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1133 net1134 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__buf_4
XANTENNA__10897__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1144 net1198 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_2
Xfanout1155 net1162 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1166 net1171 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__buf_2
Xfanout1177 net1179 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_4
X_14984_ net1238 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1188 net1198 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_2
Xfanout1199 net1265 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_4
X_13935_ net1219 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
X_16723_ net1278 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XANTENNA__09503__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16654_ clknet_leaf_100_wb_clk_i _02773_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13866_ net1233 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08509__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15605_ clknet_leaf_43_wb_clk_i _01745_ _00413_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12817_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[1\]
+ team_02_WB.instance_to_wrap.top.a1.state\[0\] _03317_ vssd1 vssd1 vccd1 vccd1 _07340_
+ sky130_fd_sc_hd__and4b_1
X_16585_ clknet_leaf_93_wb_clk_i _02704_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dfxtp_1
X_13797_ net1651 _03282_ net960 vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_100_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15536_ clknet_leaf_39_wb_clk_i _01676_ _00344_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12748_ _04568_ _04609_ _04948_ _06113_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__or4_1
XFILLER_0_85_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15467_ clknet_leaf_116_wb_clk_i _01607_ _00275_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12465__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ net265 net2124 net430 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14418_ net1122 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15398_ clknet_leaf_42_wb_clk_i _01538_ _00206_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14349_ net1154 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
Xhold605 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold638 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09990__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11809__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08910_ net1045 _04196_ _04208_ net1008 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__a32o_1
X_16019_ clknet_leaf_55_wb_clk_i _02159_ _00827_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_09890_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\] net898 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ net1631 net1039 net1035 team_02_WB.instance_to_wrap.ramstore\[23\] vssd1
+ vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a22o_1
XANTENNA__09742__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1305 team_02_WB.instance_to_wrap.ramload\[14\] vssd1 vssd1 vccd1 vccd1 net2763
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08772_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\] net686 net843 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07723_ _03416_ _03445_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07654_ _03369_ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10668__B _05580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09258__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07585_ net2321 _03311_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1086_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09324_ _04834_ _04836_ _04838_ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__nor4_1
XFILLER_0_118_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16245__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09255_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\] net925 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\]
+ _04771_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold1194_A team_02_WB.instance_to_wrap.top.a1.row2\[33\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1253_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08206_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] _03858_ vssd1 vssd1 vccd1
+ vccd1 _03924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09186_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\] net750 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\]
+ _04697_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a221o_1
XANTENNA__08769__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08137_ _03812_ _03850_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__xor2_2
XFILLER_0_82_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09430__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08068_ _03770_ _03787_ _03775_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__o21a_1
XANTENNA__09981__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout880_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11719__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09194__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\] net900 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08941__B1 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ net258 net2324 net479 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13720_ _03015_ net949 _03234_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10932_ net416 _06438_ _06441_ net376 _06445_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ net1467 _04167_ net851 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__mux2_1
X_10863_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12602_ net353 net2732 net440 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16370_ clknet_leaf_5_wb_clk_i _02510_ _01178_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13582_ team_02_WB.instance_to_wrap.top.a1.row1\[16\] _03111_ _03118_ team_02_WB.instance_to_wrap.top.a1.row2\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10794_ _06306_ _06309_ net367 vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15321_ clknet_leaf_120_wb_clk_i _01464_ _00134_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12533_ net339 net2625 net448 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12285__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15252_ clknet_leaf_63_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[11\]
+ _00065_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_10_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12464_ net328 net2522 net452 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14203_ net1159 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11415_ net994 _06910_ _06912_ _06837_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__a211o_1
X_15183_ net1239 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
X_12395_ net312 net2308 net458 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__mux2_1
XANTENNA__08999__A team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14134_ net1136 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
XANTENNA__10031__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ _05292_ net661 net658 _05293_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_91_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14065_ net1118 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
X_11277_ _06037_ _06770_ _06778_ _06779_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08511__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13016_ _07449_ _07535_ _07450_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__o21a_1
XANTENNA__09724__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\] net892 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2 team_02_WB.instance_to_wrap.top.pad.button_control.debounce vssd1 vssd1 vccd1
+ vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\] net913 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14967_ net1122 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10769__A _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13284__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10098__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16706_ net1444 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_102_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13918_ net1203 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
X_14898_ net1124 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13849_ net1224 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
X_16637_ clknet_leaf_101_wb_clk_i _02756_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13036__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16568_ clknet_leaf_97_wb_clk_i _02692_ _01375_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11598__A2 _07083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12195__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15519_ clknet_leaf_109_wb_clk_i _01659_ _00327_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16499_ clknet_leaf_35_wb_clk_i _02633_ _01306_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09040_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\] net836 net823 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\]
+ _04552_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold402 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold413 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10022__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold424 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold435 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09963__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold446 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11539__S net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold468 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09942_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\] net892 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\]
+ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold479 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout904 _04525_ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_70_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout915 _04518_ vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__buf_4
Xfanout926 _04511_ vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__buf_6
XANTENNA__09715__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16787__1331 vssd1 vssd1 vccd1 vccd1 _16787__1331/HI net1331 sky130_fd_sc_hd__conb_1
X_09873_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\] net843 _05386_ _05387_
+ _05389_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__a2111o_1
Xfanout937 _02955_ vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_2
XANTENNA_fanout294_A _06791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 _04178_ vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_2
Xhold1102 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ net135 net1044 net991 net1518 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a22o_1
Xhold1113 team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] vssd1 vssd1 vccd1 vccd1
+ net2571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1135 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ net848 _04363_ _04368_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__and3_4
Xhold1157 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout461_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1168 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1179 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ _03399_ _03400_ net425 vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a21boi_2
XANTENNA__10089__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__A1 _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ _04312_ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10398__B _05690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07637_ team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] _03329_ _03356_ _03359_ vssd1
+ vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA_fanout726_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07568_ team_02_WB.instance_to_wrap.top.ru.state\[0\] vssd1 vssd1 vccd1 vccd1 _03308_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09100__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09307_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\] net755 net703 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11589__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09238_ net539 vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__inv_2
XANTENNA__10261__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13220__A2_N net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\] _04559_ _04676_
+ _04685_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ team_02_WB.instance_to_wrap.top.pc\[20\] _06264_ vssd1 vssd1 vccd1 vccd1
+ _06706_ sky130_fd_sc_hd__nor2_1
XANTENNA__10013__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ net237 net1982 net577 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ net416 net413 vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold991 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09706__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ net381 _06570_ _06571_ net376 vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10013_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\] net728 net676 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ clknet_leaf_112_wb_clk_i _02010_ _00678_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ net1128 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10589__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14752_ net1152 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
XANTENNA__11277__A1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11964_ net325 net1591 net587 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13703_ net1718 _03222_ _03224_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__o21a_1
X_10915_ net368 _06287_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__nand2_1
X_14683_ net1156 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11895_ net321 net2724 net487 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11029__A1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15180__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16422_ clknet_leaf_67_wb_clk_i _02557_ _01230_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13634_ net1048 _03108_ _03135_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__o21ai_1
X_10846_ net379 net796 _06347_ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__o31a_1
XFILLER_0_41_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16560__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16353_ clknet_leaf_121_wb_clk_i _02493_ _01161_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ net1049 _03107_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ _05624_ net403 _06292_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15304_ clknet_leaf_71_wb_clk_i _01448_ _00117_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12516_ net271 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\] net447 vssd1
+ vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__mux2_1
X_16284_ clknet_leaf_45_wb_clk_i _02424_ _01092_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10252__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13496_ net191 net71 net104 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__and3b_1
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15235_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[26\]
+ _00048_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_87_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12447_ net259 net2400 net450 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10004__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09945__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15166_ net1249 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
X_12378_ net237 net2561 net458 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__mux2_1
XANTENNA__10771__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14117_ net1093 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11329_ net671 _06817_ _06829_ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15097_ net1078 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09158__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14048_ net1147 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13257__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16090__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15999_ clknet_leaf_110_wb_clk_i _02139_ _00807_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11268__A1 _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ _03313_ _04184_ net1673 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_82_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09330__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08471_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] _04169_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_63_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11822__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15090__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09023_ _04297_ _04500_ _04509_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12653__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout307_A _06891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09397__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 team_02_WB.instance_to_wrap.top.d_ready vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13193__B2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold232 _02596_ vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold243 team_02_WB.instance_to_wrap.ramstore\[8\] vssd1 vssd1 vccd1 vccd1 net1701
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10173__S _04496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold265 team_02_WB.START_ADDR_VAL_REG\[11\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold276 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 team_02_WB.instance_to_wrap.top.a1.row2\[32\] vssd1 vssd1 vccd1 vccd1 net1745
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1216_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout701 _04391_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_4
Xhold298 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 _04386_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__clkbuf_8
X_09925_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] _04330_ net651 team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a22o_2
Xfanout723 _04383_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout734 _04380_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_8
Xfanout745 _04378_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_4
XANTENNA_fanout676_A _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16433__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 _04375_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_8
Xfanout767 _04372_ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_4
X_09856_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\] net866 _05357_ _05372_
+ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__a211o_1
Xfanout778 _04367_ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout789 _04362_ vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__buf_4
X_08807_ net1609 net1043 net993 team_02_WB.instance_to_wrap.ramaddr\[24\] vssd1 vssd1
+ vccd1 vccd1 _02618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09787_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\] net778 net843 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\]
+ _05303_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__a221o_1
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout843_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11259__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08738_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] _04363_ _04365_ vssd1
+ vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__and3_4
XANTENNA__11259__B2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09321__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08669_ _04295_ _04296_ _04297_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11732__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ _06216_ _06215_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11680_ _04928_ _04947_ _04994_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_42_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10631_ team_02_WB.instance_to_wrap.top.pc\[26\] _06147_ vssd1 vssd1 vccd1 vccd1
+ _06148_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_27_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13350_ net1683 net1016 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[12\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10234__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10562_ net542 net405 vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13708__B1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12301_ net330 net2460 net571 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__mux2_1
XANTENNA__12563__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ _06731_ _02959_ team_02_WB.instance_to_wrap.top.pc\[19\] net1053 vssd1 vssd1
+ vccd1 vccd1 _02990_ sky130_fd_sc_hd__a2bb2o_1
X_10493_ _05468_ _06009_ _05994_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_134_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15020_ net1229 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
XANTENNA__09388__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13184__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ net2481 net321 net618 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__mux2_1
XANTENNA__09927__A2 _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11195__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12163_ net304 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\] net462 vssd1
+ vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11114_ _06267_ _06622_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12094_ net2080 net299 net584 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13487__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15175__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15922_ clknet_leaf_3_wb_clk_i _02062_ _00730_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11045_ net673 _06533_ _06555_ net672 _06554_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__a221o_2
XANTENNA__11498__B2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15800__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15853_ clknet_leaf_24_wb_clk_i _01993_ _00661_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14804_ net1074 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
X_15784_ clknet_leaf_15_wb_clk_i _01924_ _00592_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12996_ team_02_WB.instance_to_wrap.top.pc\[15\] _06197_ _07515_ vssd1 vssd1 vccd1
+ vccd1 _07516_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09312__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14735_ net1121 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
X_11947_ net257 net2584 net587 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13423__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14666_ net1139 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ _06498_ net2358 net486 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08517__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16405_ clknet_leaf_66_wb_clk_i _02540_ _01213_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13617_ _03164_ _03168_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__nor2_1
X_16786__1330 vssd1 vssd1 vccd1 vccd1 _16786__1330/HI net1330 sky130_fd_sc_hd__conb_1
XFILLER_0_131_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10829_ net547 net405 _06317_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__a21o_1
X_14597_ net1087 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11422__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16336_ clknet_leaf_39_wb_clk_i _02476_ _01144_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13548_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ _03289_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__and3_2
XFILLER_0_54_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09091__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16267_ clknet_leaf_115_wb_clk_i _02407_ _01075_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10782__A _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12473__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13479_ team_02_WB.START_ADDR_VAL_REG\[19\] net1070 _04259_ vssd1 vssd1 vccd1 vccd1
+ net202 sky130_fd_sc_hd__a21o_1
XFILLER_0_124_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15218_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[9\]
+ _00031_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09379__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09918__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16198_ clknet_leaf_44_wb_clk_i _02338_ _01006_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07929__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15330__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15149_ net1246 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ _03684_ _03693_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__nand2_1
XANTENNA__13478__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\] net769 net761 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__a22o_1
XANTENNA__11817__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11489__A1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09551__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\] net906 net939 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\] net740 _05086_ _05088_
+ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_65_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08523_ team_02_WB.instance_to_wrap.top.a1.data\[3\] net958 vssd1 vssd1 vccd1 vccd1
+ _04211_ sky130_fd_sc_hd__or2_1
XANTENNA__12648__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10957__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout257_A _06530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ _03307_ _04154_ _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10676__B _05740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08385_ _04072_ _04077_ _04083_ _04078_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__o31a_1
XFILLER_0_129_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout424_A _05715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1166_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10216__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09082__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12383__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09006_ _04295_ net943 _04505_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__and3_4
XANTENNA__09909__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12913__A1 _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09790__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15823__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13469__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\] net724 net716 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\]
+ _05424_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__a221o_1
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout564 _07219_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_4
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_6
XANTENNA__13205__A1_N net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout586 _07202_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout597 _07191_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_6
X_09839_ _05355_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__inv_2
XANTENNA__10152__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12919__A2_N _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15973__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ net526 _06190_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ net361 net1957 net595 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12558__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _06637_ _06696_ _06751_ _07304_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__and4_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14520_ net1195 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
XANTENNA__13243__A _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11732_ net359 net2485 net601 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10586__B _06102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14451_ net1166 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11663_ _07141_ _07148_ _05913_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__or3b_1
XFILLER_0_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13402_ team_02_WB.instance_to_wrap.ramload\[31\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[31\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07608__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10614_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__inv_2
XANTENNA__10207__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14382_ net1114 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
XANTENNA__09073__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11594_ net795 _07074_ _07082_ net656 _07081_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_49_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16121_ clknet_leaf_17_wb_clk_i _02261_ _00929_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13333_ net1055 team_02_WB.instance_to_wrap.top.ru.state\[2\] net1484 vssd1 vssd1
+ vccd1 vccd1 _00010_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11698__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15353__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12293__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10545_ _05314_ net402 vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08820__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ clknet_leaf_12_wb_clk_i _02192_ _00860_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13157__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13264_ net1520 net985 net966 _02980_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__a22o_1
X_10476_ _05419_ net518 vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15003_ net1228 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
XANTENNA__12904__A1 _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ net1858 net249 net616 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__mux2_1
XANTENNA__10107__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13195_ net1026 _02952_ net1023 team_02_WB.instance_to_wrap.top.pc\[2\] vssd1 vssd1
+ vccd1 vccd1 _01483_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_104_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12146_ net247 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\] net462 vssd1
+ vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09781__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12077_ net1697 net241 net584 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09533__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15905_ clknet_leaf_124_wb_clk_i _02045_ _00713_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11028_ _06385_ _06394_ net393 vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__mux2_1
X_16885_ net1429 vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__buf_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15836_ clknet_leaf_45_wb_clk_i _01976_ _00644_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12468__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15767_ clknet_leaf_116_wb_clk_i _01907_ _00575_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12979_ _07495_ _07498_ _07493_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14718_ net1192 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13066__A2_N net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15698_ clknet_leaf_8_wb_clk_i _01838_ _00506_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14649_ net1137 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_16 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _06914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ _03854_ _03860_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__xnor2_2
XANTENNA_38 _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09064__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16319_ clknet_leaf_109_wb_clk_i _02459_ _01127_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08811__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15846__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XANTENNA__14712__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10017__A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08575__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput189 net189 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__15996__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12659__A0 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07954_ _03660_ _03664_ _03673_ _03676_ _03643_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__o32a_2
XFILLER_0_103_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13320__B2 _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ _03576_ _03577_ _03598_ _03606_ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a32o_2
XFILLER_0_39_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09624_ _05129_ _05133_ _05137_ _05140_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15226__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\] net898 net805 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_37_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12378__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08506_ net1998 net850 _03319_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09486_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\] net784 net676 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15376__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ _04135_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout806_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08368_ _04060_ _04070_ _04063_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09055__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08802__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08299_ _03983_ _04011_ _04013_ _03987_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_46_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10070__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10330_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\] _04529_ _04530_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\]
+ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13139__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10261_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\] net788 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\]
+ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12000_ net331 net2042 net480 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XANTENNA__09763__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10192_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\] net878 _05696_ _05708_
+ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__a211o_1
XANTENNA__16001__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout350 net351 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_2
Xfanout361 net363 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_121_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09515__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 _05857_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13311__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout383 _06084_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_4
X_13951_ net1213 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12902_ _07369_ _07421_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__nand2_1
X_16670_ clknet_leaf_72_wb_clk_i _02787_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13882_ net1259 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16151__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15621_ clknet_leaf_34_wb_clk_i _01761_ _00429_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12833_ _04631_ _06134_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12288__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10597__A _04464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15552_ clknet_leaf_108_wb_clk_i _01692_ _00360_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12764_ _07284_ _07285_ _07286_ _07287_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09294__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14503_ net1102 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
X_11715_ net277 net2537 net603 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15483_ clknet_leaf_126_wb_clk_i _01623_ _00291_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12695_ net325 net2705 net432 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__mux2_1
XANTENNA__11920__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11646_ net388 _07089_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14434_ net1205 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
XANTENNA__09046__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15869__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_14365_ net1086 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
Xinput36 gpio_in[21] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
XANTENNA__10536__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ net998 _07066_ net945 vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__o21ai_1
Xinput47 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13316_ net2100 net986 net967 _03007_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__a22o_1
X_16104_ clknet_leaf_16_wb_clk_i _02244_ _00912_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput58 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
Xinput69 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
X_10528_ net500 net403 vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14296_ net1220 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
Xhold809 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap517 net518 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_2
Xmax_cap539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_21_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13247_ _02967_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16035_ clknet_leaf_2_wb_clk_i _02175_ _00843_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10459_ _04996_ _05041_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13178_ net228 _07501_ _02938_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__nand3_1
XFILLER_0_62_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12129_ net304 net2095 net466 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
XANTENNA__15249__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13302__B2 _03000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07670_ _03378_ _03387_ _03390_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__a211o_4
X_16868_ net1412 vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15399__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15819_ clknet_leaf_14_wb_clk_i _01959_ _00627_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13066__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12198__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13605__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16799_ net1343 vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_133_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16644__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09340_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\] net919 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\] net783 net734 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11830__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ _03921_ _03927_ _03901_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09037__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08153_ _03828_ _03858_ _03869_ _03870_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10052__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08084_ _03804_ _03777_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16024__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12661__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1129_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09745__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout491_A _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08986_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\] _04502_ vssd1 vssd1
+ vccd1 vccd1 _04503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07937_ _03652_ _03655_ _03657_ _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__o211a_1
X_16765__1309 vssd1 vssd1 vccd1 vccd1 _16765__1309/HI net1309 sky130_fd_sc_hd__conb_1
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout756_A _04375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07868_ _03558_ _03565_ _03567_ _03590_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09607_ _05103_ _05122_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__and2_1
X_07799_ _03490_ _03491_ _03496_ _03492_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout923_A _04513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09538_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\] net738 _05043_ _05047_
+ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09276__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09469_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\] net810 net903 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\]
+ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11740__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ net945 _06989_ _06993_ net605 vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12480_ net257 net2443 net560 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__mux2_1
XANTENNA__09028__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13240__B _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11431_ _05465_ _05927_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_134_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10043__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14150_ net1074 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
XANTENNA__09984__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11362_ net999 _06861_ _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1
+ vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13101_ net229 _02873_ _06761_ net233 vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_81_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ net407 net498 vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__nand2_1
XANTENNA__12571__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14081_ net1209 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
X_11293_ net407 _06794_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09736__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ net230 _07537_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__nand2_1
XANTENNA__16517__CLK clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08988__C team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ net970 _05760_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__or2_1
XANTENNA_input52_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09200__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16744__1289 vssd1 vssd1 vccd1 vccd1 _16744__1289/HI net1289 sky130_fd_sc_hd__conb_1
Xfanout1101 net1103 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__buf_4
Xfanout1112 net1116 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_125_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] net997 _04329_ net1056
+ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__a22o_1
Xfanout1123 net1124 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_4
Xfanout1134 net1135 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__clkbuf_2
Xfanout1145 net1153 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1156 net1157 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__buf_4
Xfanout1167 net1168 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_4
XANTENNA__13296__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14983_ net1243 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
XANTENNA__15541__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1178 net1179 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11915__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1189 net1197 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__buf_4
X_16722_ net1277 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XANTENNA__15183__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13934_ net1201 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16653_ clknet_leaf_100_wb_clk_i _02772_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13865_ net1231 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15604_ clknet_leaf_15_wb_clk_i _01744_ _00412_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12816_ team_02_WB.instance_to_wrap.top.edg2.flip1 _03299_ _04305_ vssd1 vssd1 vccd1
+ vccd1 _07339_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16584_ clknet_leaf_95_wb_clk_i _02703_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dfxtp_2
XANTENNA__09267__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13796_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\]
+ _03280_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15535_ clknet_leaf_38_wb_clk_i _01675_ _00343_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _07093_ _07094_ _07270_ _07074_ _07059_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10282__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12678_ net259 net2154 net433 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__mux2_1
X_15466_ clknet_leaf_127_wb_clk_i _01606_ _00274_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10821__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10774__B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08525__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16047__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14417_ net1106 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11629_ net838 _07113_ _07115_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13220__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15397_ clknet_leaf_34_wb_clk_i _01537_ _00205_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10034__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09975__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14348_ net1071 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold606 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold617 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12481__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14279_ net1107 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold639 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16197__CLK clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07575__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16018_ clknet_leaf_3_wb_clk_i _02158_ _00826_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08840_ net1625 net1039 net1035 team_02_WB.instance_to_wrap.ramstore\[24\] vssd1
+ vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1306 team_02_WB.instance_to_wrap.ramload\[23\] vssd1 vssd1 vccd1 vccd1 net2764
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08771_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] _04296_ _04302_ net931
+ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__and4b_1
XFILLER_0_97_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13287__B1 _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11825__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07722_ _03410_ _03415_ net425 vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07653_ _03370_ _03371_ _03373_ _03374_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07584_ team_02_WB.instance_to_wrap.top.pad.count\[0\] _03310_ vssd1 vssd1 vccd1
+ vccd1 _03311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09258__A2 _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09323_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\] net787 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\]
+ _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12656__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10273__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\] net877 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1079_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08205_ _03862_ _03896_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09185_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\] net710 _04699_ _04700_
+ _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1246_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__B1 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ _03849_ _03855_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__and2_1
XANTENNA__09966__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09430__A2 _04946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08067_ _03770_ _03775_ _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nor3_1
XFILLER_0_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12391__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09718__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13278__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\] net769 net681 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11735__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ net249 net2670 net478 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09497__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ _06442_ _06443_ _06444_ net399 net383 vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10862_ net389 _06043_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__or2_1
X_13650_ net1466 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] net852 vssd1 vssd1
+ vccd1 vccd1 _02733_ sky130_fd_sc_hd__mux2_1
XANTENNA__09249__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12601_ net358 net1921 net438 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13581_ _03135_ team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] _03105_ vssd1
+ vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__or3b_1
XANTENNA__12566__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10793_ _06307_ _06308_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13251__A _06365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15320_ clknet_leaf_104_wb_clk_i _01463_ _00133_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ net332 net1927 net448 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15251_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[10\]
+ _00064_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10086__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ net321 net2746 net452 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ net998 _06911_ _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1
+ vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14202_ net1180 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
X_15182_ net1250 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
X_12394_ net306 net2740 net458 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__mux2_1
XANTENNA__09421__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08999__B team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ net1214 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11345_ net421 _06313_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15907__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14064_ net1091 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
X_11276_ net422 _06776_ _06358_ _06123_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_120_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13015_ team_02_WB.instance_to_wrap.top.pc\[27\] _06147_ _07534_ vssd1 vssd1 vccd1
+ vccd1 _07535_ sky130_fd_sc_hd__a21oi_1
X_10227_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\] net912 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a22o_1
XANTENNA__08932__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10158_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\] net820 _04529_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\]
+ _05674_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13269__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 team_02_WB.instance_to_wrap.top.ru.state\[1\] vssd1 vssd1 vccd1 vccd1 net1461
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\] net776 net689 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14966_ net1138 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09488__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16705_ net1443 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_37_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13917_ net1149 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
XANTENNA__16737__A team_02_WB.instance_to_wrap.top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14897_ net1105 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16636_ clknet_leaf_101_wb_clk_i _02755_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13848_ net1221 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11047__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12476__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__A _05440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16567_ clknet_leaf_96_wb_clk_i _02691_ _01374_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_13779_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] _03271_
+ net961 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_80_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10255__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15518_ clknet_leaf_113_wb_clk_i _01658_ _00326_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16498_ clknet_leaf_37_wb_clk_i _02632_ _01305_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09660__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15449_ clknet_leaf_17_wb_clk_i _01589_ _00257_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07713__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764__1308 vssd1 vssd1 vccd1 vccd1 _16764__1308/HI net1308 sky130_fd_sc_hd__conb_1
XFILLER_0_5_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09412__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15587__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 team_02_WB.instance_to_wrap.top.a1.row1\[108\] vssd1 vssd1 vccd1 vccd1 net1861
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold425 team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] vssd1 vssd1 vccd1 vccd1
+ net1883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold436 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold447 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09941_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\] net831 _05447_ _05457_
+ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__a211o_1
Xhold469 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout905 _04525_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout916 _04518_ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__buf_6
Xfanout927 _04511_ vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_4
X_09872_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\] net786 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\]
+ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__a221o_1
Xfanout938 _02954_ vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_8
XANTENNA__14720__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout949 _03233_ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08823_ net136 net1041 net992 net1549 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a22o_1
Xhold1103 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1125 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout287_A _06766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1136 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net847 _04363_ _04365_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__and3_4
Xhold1147 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1169 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10679__B _05785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07705_ net425 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08685_ net1056 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] team_02_WB.instance_to_wrap.top.a1.instruction\[26\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 _04314_
+ sky130_fd_sc_hd__or4_1
XANTENNA__11286__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16212__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07636_ _03357_ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07567_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__inv_2
XANTENNA__12235__A1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12386__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout719_A _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13071__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16743__1288 vssd1 vssd1 vccd1 vccd1 _16743__1288/HI net1288 sky130_fd_sc_hd__conb_1
X_09306_ net535 _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_135_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09237_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\] net721 _04747_ _04752_
+ _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09168_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\] net824 net811 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout990_A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09403__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08119_ _03829_ _03836_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\] net786 net714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ net424 net412 vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold970 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold981 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11061_ _06435_ _06439_ net392 vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__mux2_1
Xhold992 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\] net712 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__a22o_1
XANTENNA__08914__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08914__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13246__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ net1127 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ net1182 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
XANTENNA__11277__A2 _06770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11963_ net323 net2526 net587 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__mux2_1
X_13702_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\] _03222_ net1240 vssd1
+ vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10914_ net672 _06427_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__nand2_1
X_14682_ net1180 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
X_11894_ net318 net2514 net486 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09890__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16421_ clknet_leaf_67_wb_clk_i _02556_ _01229_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13633_ team_02_WB.instance_to_wrap.top.a1.row1\[109\] _03160_ _03168_ _03181_ _03182_
+ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__a2111o_1
X_10845_ _04610_ net659 net665 _04611_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_32_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12296__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16352_ clknet_leaf_118_wb_clk_i _02492_ _01160_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08075__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10776_ net505 net403 vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__nand2_1
X_13564_ _03104_ _03109_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09642__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15303_ clknet_leaf_73_wb_clk_i _01447_ _00116_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12515_ net260 net2389 net447 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13495_ team_02_WB.instance_to_wrap.top.ru.state\[4\] team_02_WB.instance_to_wrap.top.ru.state\[6\]
+ net1055 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_dready sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_114_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16283_ clknet_leaf_125_wb_clk_i _02423_ _01091_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[25\]
+ _00047_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_12446_ net249 net1803 net450 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12377_ net246 net2341 net459 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__mux2_1
X_15165_ net1247 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
X_14116_ net1126 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
X_11328_ net837 _06828_ _06827_ _06826_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15096_ net1098 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14047_ net1175 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
X_11259_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] net494 _06762_ _04263_ net496
+ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_max_cap517_A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16235__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15998_ clknet_leaf_113_wb_clk_i _02138_ _00806_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14949_ net1126 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08470_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\] team_02_WB.instance_to_wrap.top.a1.halfData\[1\]
+ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 _04169_
+ sky130_fd_sc_hd__nand3b_1
XFILLER_0_106_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09881__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12217__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16619_ clknet_leaf_96_wb_clk_i _02738_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10228__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09633__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09022_ _04313_ net943 _04505_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__and3_4
XFILLER_0_2_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold200 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1
+ net1658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold211 net143 vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 team_02_WB.instance_to_wrap.ramaddr\[12\] vssd1 vssd1 vccd1 vccd1 net1680
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold233 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1
+ net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _02570_ vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold255 team_02_WB.instance_to_wrap.ramload\[13\] vssd1 vssd1 vccd1 vccd1 net1713
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold288 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net705 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_6
Xhold299 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] _04330_ net650 team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__a22o_2
XFILLER_0_121_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14450__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout713 _04386_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__buf_2
Xfanout724 _04383_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout735 _04380_ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1209_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout746 net749 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 _04375_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_4
X_09855_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\] net813 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\]
+ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout571_A _07217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 _04372_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__buf_8
Xfanout779 _04367_ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout669_A _05965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ net1656 net1043 net993 team_02_WB.instance_to_wrap.ramaddr\[25\] vssd1 vssd1
+ vccd1 vccd1 _02619_ sky130_fd_sc_hd__a22o_1
X_09786_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\] net742 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08737_ net848 _04360_ _04365_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__and3_4
XANTENNA__11259__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08668_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__and2_2
X_16879__1423 vssd1 vssd1 vccd1 vccd1 _16879__1423/HI net1423 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_137_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09872__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07619_ _03332_ _03335_ _03341_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__a21oi_1
X_08599_ _03309_ net1003 vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_46_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10630_ _06128_ _06146_ _04490_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_27_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09085__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11967__A0 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ _06074_ _06077_ net369 vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14625__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ net333 net2713 net571 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13280_ net1598 net983 net964 _02989_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10492_ net513 _05511_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a21o_1
XANTENNA__11719__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12231_ net2237 net318 net616 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09388__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16835__1379 vssd1 vssd1 vccd1 vccd1 _16835__1379/HI net1379 sky130_fd_sc_hd__conb_1
XFILLER_0_32_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12162_ net297 net1928 net463 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11113_ team_02_WB.instance_to_wrap.top.pc\[23\] _06266_ vssd1 vssd1 vccd1 vccd1
+ _06622_ sky130_fd_sc_hd__nor2_1
XANTENNA__16258__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12093_ net2520 net308 net583 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
XANTENNA__14360__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15921_ clknet_leaf_21_wb_clk_i _02061_ _00729_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11044_ _06027_ _06531_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09454__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08899__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11498__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15852_ clknet_leaf_20_wb_clk_i _01992_ _00660_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10170__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16763__1307 vssd1 vssd1 vccd1 vccd1 _16763__1307/HI net1307 sky130_fd_sc_hd__conb_1
X_14803_ net1169 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15783_ clknet_leaf_27_wb_clk_i _01923_ _00591_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12995_ _07470_ _07514_ vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__nor2_1
XANTENNA__11923__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14734_ net1163 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11946_ net248 net2277 net585 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14665_ net1100 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ net252 net2091 net488 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16404_ clknet_leaf_66_wb_clk_i _02539_ _01212_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13616_ _03103_ _03165_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__a21o_1
XANTENNA__09076__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10828_ net375 _06342_ _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11958__A0 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14596_ net1127 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
XANTENNA__09615__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16335_ clknet_leaf_34_wb_clk_i _02475_ _01143_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08823__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11422__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13547_ _03038_ _03057_ _03058_ _03040_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__o211a_1
XANTENNA__14535__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759_ net975 _06275_ _06274_ _06253_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16266_ clknet_leaf_128_wb_clk_i _02406_ _01074_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13478_ team_02_WB.START_ADDR_VAL_REG\[18\] net1068 net1002 vssd1 vssd1 vccd1 vccd1
+ net201 sky130_fd_sc_hd__a21o_1
XANTENNA__08533__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10782__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13281__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15217_ clknet_leaf_63_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[8\]
+ _00030_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] sky130_fd_sc_hd__dfrtp_4
X_12429_ net317 net2339 net454 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16197_ clknet_leaf_35_wb_clk_i _02337_ _01005_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15148_ net1245 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10933__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07970_ _03690_ _03691_ _03686_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__a21bo_1
X_15079_ net1252 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
X_16742__1287 vssd1 vssd1 vccd1 vccd1 _16742__1287/HI net1287 sky130_fd_sc_hd__conb_1
XANTENNA_wire637_A _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\] net884 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10161__A2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09571_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\] net764 net708 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\]
+ _05087_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11833__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ _04210_ net1581 net850 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09854__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07612__A team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11134__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09067__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08384_ _04077_ _04086_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08814__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12664__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout417_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1159_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09005_ net944 _04503_ _04507_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11177__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout786_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09907_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\] net684 net676 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout543 net545 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_2
Xfanout554 net556 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_6
Xfanout565 net568 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_6
XFILLER_0_96_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout576 _07216_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_8
X_09838_ _05348_ _05354_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__nor2_4
Xfanout587 _07202_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_6
Xfanout598 _07191_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09769_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\] net826 net911 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\]
+ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11743__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11800_ net354 net2003 net595 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12780_ _06965_ _06982_ _07002_ _07056_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_29_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11731_ net343 net2733 net603 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__mux2_1
X_14450_ net1122 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XANTENNA__09058__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11662_ net420 net502 _05914_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13401_ team_02_WB.instance_to_wrap.ramload\[30\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[30\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ net552 _06128_ _06129_ _06126_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__a31o_2
XANTENNA__08805__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12574__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11593_ net417 _06719_ _06921_ net375 _07073_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__a221o_2
X_14381_ net1141 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16120_ clknet_leaf_18_wb_clk_i _02260_ _00928_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13332_ _00008_ team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] vssd1 vssd1 vccd1
+ vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[4\] sky130_fd_sc_hd__or2_1
X_10544_ _05356_ net384 vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__nor2_1
XANTENNA_input82_A wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16051_ clknet_leaf_55_wb_clk_i _02191_ _00859_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13157__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13263_ _02963_ _02979_ team_02_WB.instance_to_wrap.top.pc\[27\] net1054 vssd1 vssd1
+ vccd1 vccd1 _02980_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10475_ net518 _05419_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11168__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15002_ net1222 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12214_ net2069 net253 net619 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__mux2_1
XANTENNA__12904__A2 _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13194_ net977 _02950_ _02951_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ net243 net2415 net465 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
XANTENNA__11918__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12117__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12076_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] _04452_ _06277_ _06279_
+ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__and4_4
XFILLER_0_100_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15904_ clknet_leaf_108_wb_clk_i _02044_ _00712_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11027_ net399 _06390_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16884_ net1428 vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__buf_2
XANTENNA__10143__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15835_ clknet_leaf_128_wb_clk_i _01975_ _00643_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15766_ clknet_leaf_48_wb_clk_i _01906_ _00574_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12978_ team_02_WB.instance_to_wrap.top.pc\[2\] _05836_ _07497_ vssd1 vssd1 vccd1
+ vccd1 _07498_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09836__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717_ net1084 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11929_ net323 net2681 net484 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__mux2_1
X_15697_ clknet_leaf_50_wb_clk_i _01837_ _00505_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14648_ net1194 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_17 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_28 _06914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12484__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_39 _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16423__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ net1174 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16318_ clknet_leaf_112_wb_clk_i _02458_ _01126_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10603__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16249_ clknet_leaf_17_wb_clk_i _02389_ _01057_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16573__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16878__1422 vssd1 vssd1 vccd1 vccd1 _16878__1422/HI net1422 sky130_fd_sc_hd__conb_1
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11828__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15096__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput179 net179 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07953_ _03601_ _03663_ _03674_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__and3b_1
XFILLER_0_128_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13320__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07884_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] _03543_ _03575_ vssd1 vssd1
+ vccd1 vccd1 _03607_ sky130_fd_sc_hd__or3_1
XANTENNA__10134__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\] net777 _05138_ _05139_
+ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12659__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09554_ _05064_ _05066_ _05068_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__or4_1
XANTENNA__09288__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09827__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08505_ net1046 _04185_ _04197_ _04198_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a31o_1
X_16834__1378 vssd1 vssd1 vccd1 vccd1 _16834__1378/HI net1378 sky130_fd_sc_hd__conb_1
X_09485_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\] net736 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a22o_1
XANTENNA__08990__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08436_ _04137_ _04140_ _04139_ _04130_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_77_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12394__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08367_ _04053_ _04074_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13188__A2_N net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ _03978_ _03985_ _04012_ _03962_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09460__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13139__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16762__1306 vssd1 vssd1 vccd1 vccd1 _16762__1306/HI net1306 sky130_fd_sc_hd__conb_1
XFILLER_0_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14903__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\] net784 net736 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a22o_1
XANTENNA__09212__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12898__A1 _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10191_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\] net833 net829 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\]
+ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10373__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout340 _07030_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout351 _07126_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11039__A _06549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13311__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout373 net374 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_2
X_13950_ net1213 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
Xfanout384 net385 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_2
XANTENNA__10125__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__dlymetal6s2s_1
X_12901_ _05187_ _06192_ _07420_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12569__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13881_ net1239 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
XANTENNA__13254__A _06415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15620_ clknet_leaf_2_wb_clk_i _01760_ _00428_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12832_ _07350_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__nor2_1
XANTENNA__09279__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08348__A team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10597__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15551_ clknet_leaf_86_wb_clk_i _01691_ _00359_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12822__A1 _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12763_ _04782_ _04864_ _04995_ _05040_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__or4_1
X_14502_ net1072 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11714_ net282 net2223 net603 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15482_ clknet_leaf_120_wb_clk_i _01622_ _00290_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12694_ net322 net2723 net432 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14433_ net1210 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
X_11645_ _05902_ net663 _06116_ _07128_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__o2bb2a_1
X_16741__1286 vssd1 vssd1 vccd1 vccd1 _16741__1286/HI net1286 sky130_fd_sc_hd__conb_1
XFILLER_0_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ net1152 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ _06254_ _07065_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__or2_1
XANTENNA__09451__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 gpio_in[22] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
Xinput48 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_16103_ clknet_leaf_29_wb_clk_i _02243_ _00911_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10061__A1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13315_ team_02_WB.instance_to_wrap.top.pc\[2\] net1051 _07104_ net933 vssd1 vssd1
+ vccd1 vccd1 _03007_ sky130_fd_sc_hd__a22o_2
Xinput59 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_10527_ _06041_ _06043_ net389 vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14295_ net1173 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap529 net530 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_126_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16034_ clknet_leaf_124_wb_clk_i _02174_ _00842_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13246_ net935 _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__nand2_1
X_10458_ _05127_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nand2_1
XANTENNA__09203__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13177_ _07489_ _07490_ _07500_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__nand3b_1
X_10389_ _05832_ _05905_ _05829_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10364__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12128_ net297 net2111 net469 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13302__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ net302 net1895 net471 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__mux2_1
XANTENNA__10116__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16867_ net1411 vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__buf_2
XANTENNA__12479__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10788__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15818_ clknet_leaf_128_wb_clk_i _01958_ _00626_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16798_ net1342 vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_87_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09809__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15749_ clknet_leaf_34_wb_clk_i _01889_ _00557_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09270_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\] net711 _04785_ _04786_
+ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08221_ _03936_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _03828_ _03858_ _03869_ _03870_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__o31a_1
XFILLER_0_83_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13204__A1_N _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09442__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08083_ _03771_ _03776_ _03787_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21o_1
XANTENNA__15963__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08548__A2 _04200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13219__A1_N net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10355__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1024_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] net951 vssd1 vssd1 vccd1
+ vccd1 _04502_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout484_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ _03646_ _03658_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11304__B2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07867_ _03558_ net329 _03565_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15343__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12389__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09606_ net531 _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07798_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09537_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\] net843 _05048_ _05050_
+ _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_6_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout916_A _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15493__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09468_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\] net923 net899 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10291__A1 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08419_ _04114_ _04121_ _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__or3_1
XANTENNA__08736__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09399_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\] net718 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ net666 _06918_ _06925_ net656 _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _06261_ _06860_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10312_ net396 net498 vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__or2_2
XFILLER_0_21_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13100_ _07368_ _07370_ _07422_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11292_ _06744_ _06793_ net371 vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__mux2_1
X_14080_ net1154 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13031_ net1027 _02816_ net1025 team_02_WB.instance_to_wrap.top.pc\[30\] vssd1 vssd1
+ vccd1 vccd1 _01511_ sky130_fd_sc_hd__a2bb2o_1
X_10243_ _05754_ _05757_ _05758_ _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__or4_2
XFILLER_0_63_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10346__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1102 net1103 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__buf_2
X_10174_ net505 _05690_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__nor2_1
Xfanout1113 net1116 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_4
Xfanout1124 net1125 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_4
Xfanout1135 net1144 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1146 net1153 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_4
Xfanout1157 net1162 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__buf_4
X_14982_ net1245 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
XANTENNA__13296__B2 _02997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1168 net1170 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__buf_4
Xfanout1179 net1198 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16721_ net1449 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
X_13933_ net1219 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12299__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08711__A2 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16652_ clknet_leaf_100_wb_clk_i _02771_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13864_ net1231 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
XANTENNA__13048__B2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15836__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15603_ clknet_leaf_56_wb_clk_i _01743_ _00411_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12815_ team_02_WB.instance_to_wrap.top.pc\[1\] team_02_WB.instance_to_wrap.top.testpc.en_latched
+ _07327_ _07336_ net1028 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__a32o_1
XANTENNA__08509__C _04200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16583_ clknet_leaf_95_wb_clk_i _02702_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__dfxtp_1
X_13795_ _03282_ _03283_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__nor2_1
X_16877__1421 vssd1 vssd1 vccd1 vccd1 _16877__1421/HI net1421 sky130_fd_sc_hd__conb_1
XFILLER_0_9_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11931__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ clknet_leaf_25_wb_clk_i _01674_ _00342_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12746_ _07269_ _07040_ _07023_ _07265_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__and4b_1
XANTENNA__09672__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07710__A team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15465_ clknet_leaf_105_wb_clk_i _01605_ _00273_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12677_ net249 net2672 net430 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_1
XANTENNA__15986__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14416_ net1077 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
X_11628_ _05996_ net664 _06116_ _05878_ _07114_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15396_ clknet_leaf_0_wb_clk_i _01536_ _00204_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14347_ net1200 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11559_ team_02_WB.instance_to_wrap.top.pc\[5\] net973 _04347_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\]
+ _07049_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold607 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold618 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold629 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14278_ net1089 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
X_16017_ clknet_leaf_22_wb_clk_i _02157_ _00825_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13229_ net1618 net1019 net938 _05760_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__a22o_1
X_16833__1377 vssd1 vssd1 vccd1 vccd1 _16833__1377/HI net1377 sky130_fd_sc_hd__conb_1
XFILLER_0_110_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11534__A1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11534__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_08770_ _04302_ net848 _04364_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__and3_4
XFILLER_0_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13287__B2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07721_ _03410_ net425 vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__nand2_1
XANTENNA__11298__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12002__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _03373_ _03374_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16761__1305 vssd1 vssd1 vccd1 vccd1 _16761__1305/HI net1305 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07583_ net1864 net1064 net34 vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11841__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\] net727 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13341__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09253_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\] net810 net883 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\]
+ _04769_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout232_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ _03917_ _03920_ _03903_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__a21o_2
XFILLER_0_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09184_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\] net778 net722 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\]
+ _04696_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a221o_1
XANTENNA__09415__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08135_ _03852_ _03854_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__and2b_1
XANTENNA__08769__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1141_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1239_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16141__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _03787_ _03321_ net1007 net1780 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13158__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout699_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15709__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16291__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\] net716 _04471_ _04484_
+ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__a211o_1
X_16740__1285 vssd1 vssd1 vccd1 vccd1 _16740__1285/HI net1285 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_51_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07919_ _03601_ _03639_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_51_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08899_ net27 net1031 net989 net2393 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10930_ _06323_ _06340_ net391 vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_92_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10861_ _06375_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11751__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ net341 net2446 net440 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13580_ net1049 _03115_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__nand2_1
XANTENNA__09654__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10792_ _05271_ net402 vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12531_ net335 net2216 net448 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15250_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[9\]
+ _00063_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09406__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12462_ net320 net2386 net450 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14201_ net1140 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11413_ team_02_WB.instance_to_wrap.top.pc\[12\] _06259_ vssd1 vssd1 vccd1 vccd1
+ _06911_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15181_ net1238 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XANTENNA__12582__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12393_ net296 net2167 net459 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14132_ net1091 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11344_ _05935_ _06843_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15389__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14063_ net1165 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
XANTENNA__09176__B _04692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11275_ _05980_ _06110_ _06775_ _06104_ _06777_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13014_ _07451_ _07533_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__nor2_1
XANTENNA__09185__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\] net896 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a22o_1
XANTENNA__11926__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\] net929 net925 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4 _00011_ vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10088_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\] net761 net732 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__a22o_1
X_14965_ net1217 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11227__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13916_ net1204 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
X_16704_ net1442 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XANTENNA__10131__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09893__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14896_ net1077 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16635_ clknet_leaf_101_wb_clk_i _02754_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_13847_ net1224 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14538__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16566_ clknet_leaf_92_wb_clk_i _02690_ _01373_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13778_ _03271_ _03272_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09645__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10785__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15517_ clknet_leaf_51_wb_clk_i _01657_ _00325_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12729_ _06585_ _06792_ _06817_ _07252_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__or4b_1
XFILLER_0_127_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16497_ clknet_leaf_30_wb_clk_i _02631_ _01304_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15448_ clknet_leaf_54_wb_clk_i _01588_ _00256_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16164__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12492__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15379_ clknet_leaf_78_wb_clk_i _01519_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold404 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold415 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold426 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold448 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09940_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\] net876 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold459 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11507__B2 _06084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout906 net909 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout917 _04518_ vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_2
X_09871_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\] net742 net722 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__a22o_1
Xfanout928 _04511_ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_8
Xfanout939 net940 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_4
XFILLER_0_123_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11836__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ net1531 net1041 net990 net2762 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10191__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1104 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net848 _04368_ _04370_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__and3_1
Xhold1148 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07704_ _03420_ _03425_ _03426_ _03393_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a22o_1
XANTENNA__10041__A _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08684_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09884__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07635_ team_02_WB.instance_to_wrap.top.a1.dataIn\[30\] _03324_ _03328_ vssd1 vssd1
+ vccd1 vccd1 _03358_ sky130_fd_sc_hd__and3_1
XANTENNA__12667__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1091_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1189_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07566_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 _03306_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09636__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10246__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ net971 _04821_ net543 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__o21a_1
XANTENNA__09100__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09236_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\] net767 net689 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09167_ _04678_ _04680_ _04682_ _04683_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15531__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13097__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14183__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08118_ _03793_ _03830_ _03831_ _03790_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__a22o_1
XANTENNA__08611__A1 team_02_WB.START_ADDR_VAL_REG\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\] net778 net730 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\]
+ _04612_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout983_A _02956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ _03763_ _03764_ _03769_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_129_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14911__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold960 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold971 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold982 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
X_16876__1420 vssd1 vssd1 vccd1 vccd1 _16876__1420/HI net1420 sky130_fd_sc_hd__conb_1
X_11060_ _06440_ _06444_ net393 vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__mux2_1
XANTENNA__15681__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold993 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11746__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _05516_ _05520_ _05524_ _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__or4_2
XANTENNA__08914__A2 _04203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10182__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16037__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ net1193 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
X_11962_ net319 net1762 net585 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09875__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13701_ _03222_ _03223_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10913_ _04695_ _06031_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12577__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14681_ net1136 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11893_ net315 net2203 net486 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11481__S net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16420_ clknet_leaf_67_wb_clk_i _02555_ _01228_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13632_ team_02_WB.instance_to_wrap.top.a1.row1\[13\] _03109_ _03114_ _03117_ team_02_WB.instance_to_wrap.top.a1.row1\[61\]
+ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__a32o_1
XANTENNA__16187__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10844_ net423 _06354_ _06357_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09627__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16832__1376 vssd1 vssd1 vccd1 vccd1 _16832__1376/HI net1376 sky130_fd_sc_hd__conb_1
XFILLER_0_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16351_ clknet_leaf_109_wb_clk_i _02491_ _01159_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13563_ net1047 net1049 _03290_ _03103_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__and4_1
X_10775_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__nand2_1
XANTENNA__08075__B _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15302_ clknet_leaf_71_wb_clk_i _01446_ _00115_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12514_ net264 net2246 net447 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__mux2_1
X_16282_ clknet_leaf_119_wb_clk_i _02422_ _01090_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13494_ net1668 _04286_ _04289_ net2229 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_read_i
+ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_97_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[24\]
+ _00046_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15189__A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12445_ net253 net2143 net452 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15164_ net1246 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
X_12376_ net243 net1779 net461 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__mux2_1
X_16760__1304 vssd1 vssd1 vccd1 vccd1 _16760__1304/HI net1304 sky130_fd_sc_hd__conb_1
X_14115_ net1130 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11327_ _05939_ _05988_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__xnor2_1
X_15095_ net1104 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09158__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ net1194 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11258_ _06761_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10209_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\] net770 _05724_ _05725_
+ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_108_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11189_ net546 net397 _06692_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__or3_1
X_15997_ clknet_leaf_48_wb_clk_i _02137_ _00805_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14948_ net1127 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
XANTENNA__09866__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09330__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14879_ net1186 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12487__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16618_ clknet_leaf_98_wb_clk_i _02737_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09618__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16549_ clknet_leaf_96_wb_clk_i _02673_ _01356_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13900__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09021_ _04313_ net944 _04505_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and3_1
XANTENNA__15099__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09397__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 team_02_WB.instance_to_wrap.ramload\[25\] vssd1 vssd1 vccd1 vccd1 net1659
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold212 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1
+ net1670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 _02606_ vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold234 team_02_WB.instance_to_wrap.ramstore\[4\] vssd1 vssd1 vccd1 vccd1 net1692
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 team_02_WB.instance_to_wrap.ramaddr\[21\] vssd1 vssd1 vccd1 vccd1 net1703
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 team_02_WB.instance_to_wrap.top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1 net1725
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09149__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09923_ net515 vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__inv_2
Xfanout703 net705 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_4
Xhold289 net131 vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 net717 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_8
Xfanout725 _04383_ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout397_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout736 _04380_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_8
Xfanout747 net749 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_4
X_09854_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\] net910 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a22o_1
XANTENNA__10164__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout758 _04374_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1104_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 _04372_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
X_08805_ net1515 net1043 net993 net2760 vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a22o_1
X_09785_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\] net782 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout564_A _07219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08736_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__and3b_2
XANTENNA__09321__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08667_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout731_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout829_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13082__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] _03329_ _03338_ _03340_ vssd1
+ vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _04250_ _04251_ _04253_ _04258_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_46_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1
+ _03290_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10560_ _06075_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13169__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\] net703 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09719__B net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ net513 _05511_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_44_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12230_ net2430 net315 net616 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__mux2_1
XANTENNA__09388__A2 _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12161_ net309 net2120 net463 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11112_ _04494_ net654 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] net496
+ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__a221o_1
XANTENNA__09735__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ net2552 net303 net583 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
Xhold790 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15920_ clknet_leaf_40_wb_clk_i _02060_ _00728_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11043_ _06551_ _06552_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10155__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15427__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15851_ clknet_leaf_115_wb_clk_i _01991_ _00659_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14802_ net1119 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
X_15782_ clknet_leaf_50_wb_clk_i _01922_ _00590_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09848__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ _07471_ _07513_ _07472_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09312__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14733_ net1143 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11945_ net253 net1783 net588 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
XANTENNA__15577__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14664_ net1178 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12100__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ net238 net2335 net486 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ clknet_leaf_65_wb_clk_i _02538_ _01211_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13615_ team_02_WB.instance_to_wrap.top.lcd.nextState\[4\] _03105_ _03113_ _03165_
+ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__a32o_1
X_10827_ _05715_ _06313_ _06329_ net379 vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__o22a_1
X_14595_ net1131 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16334_ clknet_leaf_26_wb_clk_i _02474_ _01142_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13546_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _03061_ _03092_ net1067
+ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__o211a_1
X_10758_ _06242_ _06246_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16265_ clknet_leaf_105_wb_clk_i _02405_ _01073_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13477_ team_02_WB.START_ADDR_VAL_REG\[17\] _04260_ vssd1 vssd1 vccd1 vccd1 net200
+ sky130_fd_sc_hd__and2_1
X_10689_ _03294_ _06203_ _06205_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15216_ clknet_leaf_58_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[7\]
+ _00029_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12907__B1 _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ net312 net2194 net454 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09379__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16196_ clknet_leaf_1_wb_clk_i _02336_ _01004_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15147_ net1244 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12359_ net311 net2379 net563 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10933__A2 _05901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15078_ net1252 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14029_ net1133 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
XANTENNA__13167__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09000__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10146__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire532_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09551__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09570_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\] net780 net716 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08521_ net1046 _04208_ _04209_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12010__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ _04145_ _04153_ _04148_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_19_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08383_ _04082_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08814__B2 net1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09004_ _04297_ net944 _04503_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__and3_4
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12680__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14461__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09790__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout779_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16831__1375 vssd1 vssd1 vccd1 vccd1 _16831__1375/HI net1375 sky130_fd_sc_hd__conb_1
X_09906_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\] net764 net748 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10137__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_2
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_8
XFILLER_0_22_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout566 net568 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09542__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\] net742 _05350_ _05352_
+ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__a2111o_1
Xfanout577 net580 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_6
Xfanout588 _07202_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_4
Xfanout599 _07191_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout946_A _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09768_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\] net863 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__a22o_1
X_08719_ net1058 _04277_ _04323_ _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09699_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\] net721 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\]
+ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_29_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11730_ net338 net2491 net604 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _05624_ _05646_ _05920_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__or3b_1
XFILLER_0_77_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13400_ team_02_WB.instance_to_wrap.ramload\[29\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[29\] sky130_fd_sc_hd__and2_1
X_10612_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] net995 vssd1 vssd1 vccd1
+ vccd1 _06129_ sky130_fd_sc_hd__nand2_1
X_14380_ net1073 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ net666 _07076_ _07078_ _07080_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13331_ net1491 _03013_ _03010_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[3\]
+ sky130_fd_sc_hd__or3b_1
X_10543_ net388 _06055_ _06056_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__a31o_1
XANTENNA__16225__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16050_ clknet_leaf_3_wb_clk_i _02190_ _00858_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13262_ _06490_ _02962_ _02959_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a21o_1
XANTENNA_input75_A wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10474_ _05314_ _05334_ _05377_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15001_ net1228 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
XANTENNA__11168__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ net1765 net240 net616 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__mux2_1
XANTENNA__12590__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ net231 _02949_ team_02_WB.instance_to_wrap.top.pc\[2\] net232 vssd1 vssd1
+ vccd1 vccd1 _02951_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10376__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ net647 _07212_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__nand2_1
XANTENNA__09781__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13314__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ net346 net1832 net470 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10404__A _05579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09533__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ net397 _06395_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__or2_1
X_15903_ clknet_leaf_112_wb_clk_i _02043_ _00711_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_16883_ net1427 vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__buf_2
XFILLER_0_95_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11934__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15834_ clknet_leaf_117_wb_clk_i _01974_ _00642_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11628__B1 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15765_ clknet_leaf_41_wb_clk_i _01905_ _00573_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12977_ _07334_ _07496_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11235__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11928_ net317 net2605 net482 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__mux2_1
X_14716_ net1146 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
X_15696_ clknet_leaf_39_wb_clk_i _01836_ _00504_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14647_ net1172 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
X_11859_ net312 net2517 net490 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14546__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14578_ net1124 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_29 _06914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16317_ clknet_leaf_50_wb_clk_i _02457_ _01125_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13529_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] _03061_ _03080_ _03089_
+ net1067 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16248_ clknet_leaf_19_wb_clk_i _02388_ _01056_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_109_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16179_ clknet_leaf_54_wb_clk_i _02319_ _00987_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_112_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10367__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XANTENNA__13305__B1 _07007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ _03663_ _03674_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__nand2_1
XANTENNA__12005__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07883_ net316 _03597_ _03578_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11844__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\] net772 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13344__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\] net940 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\]
+ _05069_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08504_ team_02_WB.instance_to_wrap.top.a1.row1\[16\] net850 vssd1 vssd1 vccd1 vccd1
+ _04198_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09484_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\] net700 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08435_ _04139_ _04140_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__and2b_1
XANTENNA__16248__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12675__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14456__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1171_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13360__A team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_110_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08366_ _04075_ _04076_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08297_ _03306_ _03746_ _03964_ _03972_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10070__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout896_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09285__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09763__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\] net926 net898 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_2
Xfanout341 _07051_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout352 _07087_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09515__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 _07107_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_2
Xfanout374 _06088_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_2
Xfanout385 _05901_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_2
XANTENNA__11754__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 net401 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_4
X_12900_ _07371_ _07419_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__and2_1
X_13880_ net1256 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12831_ _04589_ _06131_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12283__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15550_ clknet_leaf_113_wb_clk_i _01690_ _00358_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12762_ _05126_ _05210_ _05293_ _05379_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14501_ net1087 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
XANTENNA__08067__C _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11713_ net270 net1794 net603 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
X_15481_ clknet_leaf_111_wb_clk_i _01621_ _00289_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12693_ net319 net2464 net430 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__mux2_1
XANTENNA__12585__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14432_ net1152 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
X_11644_ _07129_ _04462_ _06114_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__or3b_1
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14363_ net1156 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11575_ team_02_WB.instance_to_wrap.top.pc\[3\] team_02_WB.instance_to_wrap.top.pc\[2\]
+ team_02_WB.instance_to_wrap.top.pc\[4\] vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__a21oi_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
X_16102_ clknet_leaf_49_wb_clk_i _02242_ _00910_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ net1963 net983 net964 _03006_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__a22o_1
Xinput38 wb_rst_i vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
X_10526_ _05995_ _06042_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__or2_1
Xinput49 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10061__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14294_ net1093 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11929__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16033_ clknet_leaf_121_wb_clk_i _02173_ _00841_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13245_ _06365_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__nand2_1
XANTENNA__15765__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ _05972_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__nor2_2
XANTENNA__10349__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11010__A1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13176_ _07398_ _07400_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10388_ _05878_ _05903_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__or2_1
XANTENNA__08962__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ net308 net1821 net468 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09923__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12058_ net295 net1993 net472 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11313__A2 _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ _06122_ _06517_ _06520_ _06509_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__a211o_1
X_16866_ net1410 vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__buf_2
XANTENNA__10788__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15817_ clknet_leaf_104_wb_clk_i _01957_ _00625_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_16797_ net1341 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11077__A1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15748_ clknet_leaf_2_wb_clk_i _01888_ _00556_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12495__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15679_ clknet_leaf_111_wb_clk_i _01819_ _00487_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08493__A2 _04185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08220_ _03916_ _03926_ _03920_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__or3b_1
XFILLER_0_12_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16830__1374 vssd1 vssd1 vccd1 vccd1 _16830__1374/HI net1374 sky130_fd_sc_hd__conb_1
XFILLER_0_114_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08151_ _03849_ _03855_ _03857_ _03826_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10052__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08082_ _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13339__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09745__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08984_ net1056 net951 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__nand2_1
X_07935_ _03614_ _03637_ _03617_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout477_A _07206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13355__A team_02_WB.instance_to_wrap.ramload\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07866_ _03558_ _03563_ _03564_ net329 vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__nand4_1
XFILLER_0_97_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09605_ net970 net630 net543 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16070__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07797_ _03491_ _03514_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09536_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\] net774 _05051_ _05052_
+ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a211o_1
XANTENNA__15638__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09130__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10815__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\] net821 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\]
+ _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout811_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08418_ _04125_ _03321_ net1005 net1981 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__a2bb2o_1
X_09398_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\] net787 _04911_ _04912_
+ _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_65_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08349_ _04047_ _04049_ _04058_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14914__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10043__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09984__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11360_ team_02_WB.instance_to_wrap.top.pc\[14\] _06260_ vssd1 vssd1 vccd1 vccd1
+ _06860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10311_ _05811_ _05817_ _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__nor3_2
XANTENNA__11749__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11291_ _05187_ net404 _06332_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13030_ net978 _02815_ _07547_ _07544_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__o211a_1
XANTENNA__09736__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\] net827 net900 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\]
+ _05745_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10173_ _05671_ net622 _04496_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__mux2_4
Xfanout1103 net1125 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_2
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1114 net1116 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_4
Xfanout1125 net1199 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1136 net1137 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__buf_4
XANTENNA_input38_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1153 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__buf_4
Xfanout1158 net1161 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__buf_4
X_14981_ net1255 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13296__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16413__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1169 net1170 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__buf_4
XANTENNA__13265__A _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16720_ net1448 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
X_13932_ net1194 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13863_ net1228 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
X_16651_ clknet_leaf_100_wb_clk_i _02770_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13048__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12814_ team_02_WB.instance_to_wrap.top.testpc.en_latched team_02_WB.instance_to_wrap.top.i_ready
+ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15602_ clknet_leaf_9_wb_clk_i _01742_ _00410_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13794_ net1869 _03280_ net960 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_104_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16582_ clknet_leaf_94_wb_clk_i _02701_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09121__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16563__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15533_ clknet_leaf_22_wb_clk_i _01673_ _00341_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12745_ _06609_ _07267_ _07268_ _06643_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_100_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10282__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15464_ clknet_leaf_20_wb_clk_i _01604_ _00272_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12676_ net251 net2099 net433 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415_ net1121 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08525__C _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11627_ _05880_ net661 vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__nand2_1
X_15395_ clknet_leaf_127_wb_clk_i _01535_ _00203_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ net1142 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
Xwire550 _04415_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10034__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ net998 _07048_ net947 vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09975__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap316 _03596_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold608 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10509_ _06018_ _06019_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__or3_1
Xhold619 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ net1087 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11489_ net657 _06356_ _06981_ _06982_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__o31a_1
XFILLER_0_69_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16016_ clknet_leaf_39_wb_clk_i _02156_ _00824_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09188__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13228_ net621 net937 net1018 net1692 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13159_ net232 _06991_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16093__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13287__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ _03431_ _03436_ _03440_ _03441_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__a211o_1
XFILLER_0_100_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire612_A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07651_ _03336_ _03341_ _03361_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__and3_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16849_ net1393 vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13903__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07582_ net2518 net1064 net35 vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\] net711 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\]
+ _04837_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15930__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09252_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\] net898 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a22o_1
XANTENNA__10273__A2 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11470__B2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08203_ _03917_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09183_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\] net774 net718 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14734__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ _03780_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10025__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09966__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__A team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08065_ _03782_ _03786_ _03755_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_114_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1134_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09718__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout594_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10733__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\] net745 net704 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_A _04374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13278__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07918_ _03627_ _03640_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08898_ net28 net1029 net987 net1808 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_123_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15460__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09351__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07849_ _03546_ net329 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14909__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10860_ _06373_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09103__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09519_ net970 net633 net544 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10791_ _05314_ net384 vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12530_ net326 net1815 net448 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12461_ net312 net2211 net450 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14200_ net1193 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11412_ _06205_ _06909_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_10_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10016__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09957__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15180_ net1238 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12392_ net310 net2180 net461 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14131_ net1166 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
X_11343_ _05294_ _05934_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09709__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14062_ net1163 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11274_ _05167_ net662 net659 _05168_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13013_ _07452_ _07532_ _07453_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__o21a_1
X_10225_ team_02_WB.instance_to_wrap.top.a1.instruction\[24\] net792 net652 _05741_
+ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__a22o_4
XFILLER_0_101_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09590__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\] net921 net799 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\]
+ _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__a221o_1
XANTENNA__13269__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 team_02_WB.instance_to_wrap.top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 net1463
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12103__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ _05579_ _05603_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__nand2_1
X_14964_ net1074 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09342__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ net1441 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11227__B _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13915_ net1216 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14895_ net1122 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
XANTENNA__10131__B _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15953__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16634_ clknet_leaf_102_wb_clk_i _02753_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13846_ net1226 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
XANTENNA__13426__C1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13777_ net2680 _03269_ net961 vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__o21ai_1
X_16565_ clknet_leaf_92_wb_clk_i _02689_ _01372_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13218__A1_N net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ _04783_ _06028_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_80_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__B _04177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15516_ clknet_leaf_45_wb_clk_i _01656_ _00324_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10255__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16309__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12728_ _06841_ _06893_ _07251_ _06867_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__nor4b_1
XTAP_TAPCELL_ROW_61_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16496_ clknet_leaf_7_wb_clk_i _02630_ _01303_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12659_ net315 net2199 net434 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__mux2_1
X_15447_ clknet_leaf_14_wb_clk_i _01587_ _00255_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12401__A0 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15378_ clknet_leaf_78_wb_clk_i _01518_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold405 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14329_ net1139 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold416 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold427 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold438 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout907 net909 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_4
XFILLER_0_110_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09870_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\] net758 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a22o_1
Xfanout918 _04515_ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout929 _04511_ vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__buf_2
XANTENNA__15483__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09581__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ net1582 net1044 net990 team_02_WB.instance_to_wrap.ramaddr\[10\] vssd1 vssd1
+ vccd1 vccd1 _02604_ sky130_fd_sc_hd__a22o_1
Xhold1105 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1116 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _04358_ _04360_ _04368_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__and3_1
Xhold1127 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1138 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12013__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1149 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ _03392_ _03421_ _03390_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09333__B1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08683_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] team_02_WB.instance_to_wrap.top.a1.instruction\[29\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] team_02_WB.instance_to_wrap.top.a1.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__or4_1
XANTENNA__10041__B _05556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07634_ team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] _03353_ team_02_WB.instance_to_wrap.top.a1.dataIn\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07565_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 _03305_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_76_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13432__A2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09304_ _04814_ _04820_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout1084_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12640__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10246__A2 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09235_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\] net674 _04748_ _04751_
+ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_131_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12683__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout607_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14464__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1251_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09166_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\] net816 net873 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\]
+ _04674_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08117_ _03793_ _03830_ _03831_ _03790_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_47_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09097_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\] net754 net726 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08048_ _03765_ _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_1400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold950 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold961 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold972 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold983 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold994 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\] net760 _05525_ _05526_
+ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_34_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\] net768 net748 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\]
+ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__a221o_1
XANTENNA__15976__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13120__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ net313 net1990 net585 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11762__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13700_ net1627 _03221_ net1065 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__o21ai_1
X_10912_ _05956_ _06425_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__or2_1
XANTENNA__07886__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14680_ net1186 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
XANTENNA__11682__A1 _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11892_ net305 net2196 net486 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13631_ team_02_WB.instance_to_wrap.top.a1.row1\[101\] _03162_ vssd1 vssd1 vccd1
+ vccd1 _03181_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10843_ net414 net397 net546 vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11434__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16350_ clknet_leaf_114_wb_clk_i _02490_ _01158_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13562_ net1048 _03113_ _03115_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__and4b_4
XFILLER_0_82_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ net500 net385 vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15301_ clknet_leaf_67_wb_clk_i _01445_ _00114_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12513_ net256 net1975 net447 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16281_ clknet_leaf_111_wb_clk_i _02421_ _01089_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15356__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13493_ _03061_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.edg2.button_i
+ sky130_fd_sc_hd__inv_2
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12593__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15232_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[23\]
+ _00045_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_12444_ net240 net1900 net450 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15163_ net1246 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
X_12375_ net645 _07195_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__nand2_4
XFILLER_0_23_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14114_ net1208 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
X_11326_ net421 _06037_ _06070_ _06104_ _06823_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__a32oi_1
X_15094_ net1098 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11937__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14045_ net1084 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11257_ team_02_WB.instance_to_wrap.top.pc\[18\] _06263_ vssd1 vssd1 vccd1 vccd1
+ _06761_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10208_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\] net754 net698 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a22o_1
XANTENNA__09563__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10173__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ _06693_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10139_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\] net732 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15996_ clknet_leaf_45_wb_clk_i _02136_ _00804_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13647__C1 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14947_ net1131 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14878_ net1191 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12870__B1 _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16131__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16617_ clknet_leaf_99_wb_clk_i _02736_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13829_ net1232 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10228__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11425__B2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16548_ clknet_leaf_97_wb_clk_i _02672_ _01355_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16479_ clknet_leaf_89_wb_clk_i net1599 _01287_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_112_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09020_ net943 _04507_ _04509_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__and3_4
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold202 net111 vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 team_02_WB.instance_to_wrap.ramstore\[18\] vssd1 vssd1 vccd1 vccd1 net1671
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 team_02_WB.instance_to_wrap.ramaddr\[24\] vssd1 vssd1 vccd1 vccd1 net1682
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold235 _02566_ vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _02615_ vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold257 team_02_WB.instance_to_wrap.ramstore\[17\] vssd1 vssd1 vccd1 vccd1 net1715
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 team_02_WB.instance_to_wrap.ramload\[28\] vssd1 vssd1 vccd1 vccd1 net1726
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11847__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold279 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\] net784 _05434_ _05435_
+ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__a2111oi_2
Xfanout704 net705 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_8
Xfanout715 net717 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_8
Xfanout726 net729 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_8
Xfanout737 _04380_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_4
X_09853_ _05363_ _05365_ _05367_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or4_1
XANTENNA__13347__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_6
Xfanout759 _04374_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout292_A _06791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ net125 net1043 net993 net1520 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a22o_1
X_09784_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\] net746 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\]
+ _05300_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__a221o_1
XANTENNA__13638__C1 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13102__A1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07580__A2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08735_ team_02_WB.instance_to_wrap.top.a1.instruction\[18\] net932 team_02_WB.instance_to_wrap.top.a1.instruction\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__and3b_2
XFILLER_0_20_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12678__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__and2_2
XFILLER_0_94_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] team_02_WB.instance_to_wrap.top.a1.dataIn\[21\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1 vccd1 _03340_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15379__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08597_ _04254_ _04255_ _04256_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout724_A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07548_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1
+ _03289_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09085__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09218_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10490_ _05559_ _06006_ net512 _05556_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_92_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__A1 _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09149_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\] net753 _04664_ _04665_
+ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a211o_1
XANTENNA__14922__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12160_ net301 net2575 net463 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__mux2_1
XANTENNA__09793__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _06230_ _06619_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11757__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ net2152 net295 net583 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
Xhold780 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 team_02_WB.START_ADDR_VAL_REG\[7\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09545__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _06038_ _06541_ _06548_ _06123_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_9_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08899__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15850_ clknet_leaf_129_wb_clk_i _01990_ _00658_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ net1118 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
X_15781_ clknet_leaf_31_wb_clk_i _01921_ _00589_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12588__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12993_ _07475_ _07512_ _07473_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__o21a_1
X_14732_ net1071 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11944_ net237 net2264 net585 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11875_ net247 net2748 net488 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
X_14663_ net1120 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16402_ clknet_leaf_65_wb_clk_i _02537_ _01210_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10826_ _06335_ _06341_ net393 vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__mux2_1
X_13614_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] _03108_ vssd1 vssd1 vccd1
+ vccd1 _03166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11407__B2 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09076__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14594_ net1208 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16333_ clknet_leaf_23_wb_clk_i _02473_ _01141_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10757_ net999 _06273_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__nor2_1
X_13545_ _03080_ _03101_ _03102_ net1067 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08823__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13476_ team_02_WB.START_ADDR_VAL_REG\[16\] net1068 net1002 vssd1 vssd1 vccd1 vccd1
+ net199 sky130_fd_sc_hd__a21o_1
X_16264_ clknet_leaf_15_wb_clk_i _02404_ _01072_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10688_ net790 _04419_ _06204_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__o21a_2
XFILLER_0_42_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08533__C _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15215_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[6\]
+ _00028_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] sky130_fd_sc_hd__dfrtp_4
X_12427_ net306 net2581 net454 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__mux2_1
X_16195_ clknet_leaf_12_wb_clk_i _02335_ _01003_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09784__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15146_ net1243 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
X_12358_ net300 net2568 net562 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ _06262_ _06810_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__or2_1
X_15077_ net1235 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
XANTENNA_max_cap522_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12289_ net272 net1995 net569 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14028_ net1073 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XANTENNA__09000__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12498__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14279__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15979_ clknet_leaf_114_wb_clk_i _02119_ _00787_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15521__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08520_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[4\] net980 vssd1 vssd1 vccd1
+ vccd1 _04209_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_65_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10600__A _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08451_ _04145_ _04153_ _04148_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__or3b_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08382_ _04059_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09067__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15671__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08275__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08814__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_118_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10082__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09003_ _04510_ _04519_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__nor2_4
XANTENNA__16027__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10909__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout305_A _06891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13049__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1214_A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09527__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09905_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\] net728 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\]
+ _05421_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout545 _04498_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_2
XANTENNA_fanout674_A _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout556 _07227_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_4
X_09836_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\] net766 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__a22o_1
Xfanout567 net568 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_6
Xfanout578 net580 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_8
Xfanout589 net592 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_6
XFILLER_0_77_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09767_ _05277_ _05279_ _05281_ _05283_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout841_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout939_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ _04268_ _04346_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__nor2_4
XANTENNA__11637__A1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09698_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\] net726 net703 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08649_ net1059 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _04278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11660_ _05738_ _05916_ _07141_ _07145_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09058__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10611_ _04283_ _04493_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__nand2_8
XFILLER_0_14_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11591_ net671 _07075_ _07079_ net837 vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08805__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10073__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13330_ team_02_WB.instance_to_wrap.top.a1.hexop\[1\] team_02_WB.instance_to_wrap.top.a1.hexop\[2\]
+ team_02_WB.instance_to_wrap.top.a1.hexop\[3\] vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__or3_1
X_10542_ net388 _06058_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ net2653 net986 net967 _02978_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ net519 _05333_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__nand2_1
X_15000_ net1228 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
X_12212_ net2285 net246 net617 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09766__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ _07390_ _07392_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input68_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09230__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ _06278_ _07190_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__nor2_1
XANTENNA__13268__A _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_88_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13314__B2 _03006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ net348 net2441 net473 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11025_ _06534_ _06535_ net413 vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__mux2_1
X_15902_ clknet_leaf_113_wb_clk_i _02042_ _00710_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16882_ net1426 vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__buf_2
XFILLER_0_99_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15833_ clknet_leaf_18_wb_clk_i _01973_ _00641_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12111__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15764_ clknet_leaf_12_wb_clk_i _01904_ _00572_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12976_ team_02_WB.instance_to_wrap.top.pc\[2\] _05835_ vssd1 vssd1 vccd1 vccd1 _07496_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14715_ net1160 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ net313 net2271 net482 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__mux2_1
X_15695_ clknet_leaf_38_wb_clk_i _01835_ _00503_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11950__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14646_ net1094 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11858_ net306 net2636 net490 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_19 _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10809_ _04755_ net404 vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13250__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14577_ net1119 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
X_11789_ net296 net2528 net594 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10064__A0 _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ clknet_leaf_45_wb_clk_i _02456_ _01124_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ _03084_ _03085_ _03087_ _03088_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__or4_1
XANTENNA__10603__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16247_ clknet_leaf_116_wb_clk_i _02387_ _01055_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13459_ team_02_WB.START_ADDR_VAL_REG\[0\] _03309_ net1003 vssd1 vssd1 vccd1 vccd1
+ _03060_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09757__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16178_ clknet_leaf_3_wb_clk_i _02318_ _00986_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XANTENNA__09221__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_2_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__13178__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
X_15129_ net1248 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_11_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09509__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ _03670_ _03672_ _03660_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__a21oi_2
XANTENNA__13305__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ _03585_ _03604_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09391__A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09621_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\] net753 net715 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09552_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\] net906 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__a22o_1
XANTENNA__12021__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12816__B1 _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ team_02_WB.instance_to_wrap.top.a1.data\[8\] net958 _04196_ vssd1 vssd1 vccd1
+ vccd1 _04197_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09483_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\] net684 _04998_ _04999_
+ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a211o_1
XANTENNA__11860__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ _04127_ _04133_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13360__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08365_ _04041_ _04054_ _04074_ _04053_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_50_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout422_A _05715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1164_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15417__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08296_ _03962_ _03988_ _03985_ _03980_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09460__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12691__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09212__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15567__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout889_A _04536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_86_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout320 _06936_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_15_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_2
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_2
Xfanout353 _07087_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_1
Xfanout364 _03496_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_4
Xfanout375 net376 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_2
XANTENNA__09920__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09819_ _05335_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__inv_2
Xfanout397 net400 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12830_ _04588_ _06130_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__nor2_1
XANTENNA__09279__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12761_ _04823_ _04909_ _05083_ _05168_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11770__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14500_ net1126 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10294__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11712_ net262 net2191 net603 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
X_15480_ clknet_leaf_53_wb_clk_i _01620_ _00288_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12692_ net315 net2304 net430 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14431_ net1170 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
X_11643_ _05995_ _06287_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__nor2_2
XFILLER_0_65_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10046__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09987__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14362_ net1181 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
X_11574_ _06583_ _07059_ _07060_ _07063_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_52_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09451__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_16101_ clknet_leaf_34_wb_clk_i _02241_ _00909_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput39 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_1
X_10525_ _05877_ net403 vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__nor2_1
X_13313_ team_02_WB.instance_to_wrap.top.pc\[3\] net1051 _07083_ net933 vssd1 vssd1
+ vccd1 vccd1 _03006_ sky130_fd_sc_hd__a22o_2
X_14293_ net1214 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13244_ _06415_ _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nand2_1
XANTENNA__09739__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16032_ clknet_leaf_106_wb_clk_i _02172_ _00840_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09476__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456_ _05080_ _05061_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and2b_1
XANTENNA__09203__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ net1026 _02936_ net1025 team_02_WB.instance_to_wrap.top.pc\[6\] vssd1 vssd1
+ vccd1 vccd1 _01487_ sky130_fd_sc_hd__a2bb2o_1
X_10387_ _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__inv_2
XANTENNA__10415__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12106__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12126_ net300 net2642 net469 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
XANTENNA__13299__B1 _06950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12057_ net286 net2679 net472 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11008_ _04777_ net663 net660 _04782_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__a221o_1
XANTENNA__09911__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16865_ net1409 vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__buf_2
X_15816_ clknet_leaf_20_wb_clk_i _01956_ _00624_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_16796_ net1340 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15747_ clknet_leaf_2_wb_clk_i _01887_ _00555_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12959_ team_02_WB.instance_to_wrap.top.pc\[11\] _05444_ vssd1 vssd1 vccd1 vccd1
+ _07479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14557__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10285__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15678_ clknet_leaf_118_wb_clk_i _01818_ _00486_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14629_ net1086 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13223__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10037__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ _03796_ _03824_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__nor2_1
XANTENNA__09978__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09442__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08081_ _03774_ net227 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__xor2_2
XFILLER_0_125_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11537__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12016__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08983_ net1056 net951 vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11855__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13636__A _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07934_ _03608_ _03653_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__xor2_4
XANTENNA__09902__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ _03556_ _03586_ _03587_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__nor3_1
XANTENNA__13355__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _05107_ _05115_ _05118_ _05120_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__nor4_1
XFILLER_0_97_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07796_ _03490_ _03497_ _03518_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09535_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\] net758 net714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12686__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10276__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09466_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\] net829 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16365__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10815__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__A team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08417_ _04113_ _04122_ _04124_ _04109_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__o2bb2a_2
X_09397_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\] net755 net711 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\]
+ _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a221o_1
XANTENNA__13214__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10028__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04059_ vssd1 vssd1 vccd1
+ vccd1 _04060_ sky130_fd_sc_hd__or2_1
XANTENNA__10579__A1 _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10934__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ _03962_ _03988_ _03976_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1
+ vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10310_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\] net784 _05818_ _05819_
+ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11290_ _05212_ _06016_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10241_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\] net823 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\]
+ _05744_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10200__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _05673_ _05684_ _05686_ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_110_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1104 net1108 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__buf_4
XANTENNA__11765__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1115 net1116 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__buf_4
Xfanout1126 net1135 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1137 net1144 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_4
X_14980_ net1238 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
Xfanout1148 net1153 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1159 net1161 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13931_ net1219 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11700__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16650_ clknet_leaf_100_wb_clk_i _02769_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13862_ net1226 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
X_15601_ clknet_leaf_19_wb_clk_i _01741_ _00409_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12813_ team_02_WB.instance_to_wrap.top.testpc.en_latched team_02_WB.instance_to_wrap.top.i_ready
+ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16581_ clknet_leaf_100_wb_clk_i _02700_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dfxtp_1
XANTENNA__12596__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13793_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\]
+ _03278_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_104_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15532_ clknet_leaf_10_wb_clk_i _01672_ _00340_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12744_ _06667_ _06700_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09672__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15463_ clknet_leaf_26_wb_clk_i _01603_ _00271_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13205__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12675_ net237 net2299 net430 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ net1164 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
X_11626_ _05902_ _05996_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__xor2_1
X_15394_ clknet_leaf_125_wb_clk_i _01534_ _00202_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_2
X_14345_ net1099 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11557_ _06255_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold609 team_02_WB.instance_to_wrap.ramload\[1\] vssd1 vssd1 vccd1 vccd1 net2067
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ _06022_ _06024_ _05984_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14276_ net1129 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
X_11488_ _06977_ _06981_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16015_ clknet_leaf_38_wb_clk_i _02155_ _00823_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13227_ net623 net936 net1020 net1851 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__a2bb2o_1
X_10439_ _04695_ _05955_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14840__A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12192__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13158_ net1026 _02922_ net1023 team_02_WB.instance_to_wrap.top.pc\[9\] vssd1 vssd1
+ vccd1 vccd1 _01490_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_97_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12109_ _06278_ _07188_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13089_ _06707_ net233 net229 _02863_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11298__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13692__B1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07650_ _03336_ _03361_ _03341_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__a21oi_1
X_16848_ net1392 vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15262__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07581_ net2050 net1064 net36 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a21o_1
X_16779_ net1323 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
X_09320_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\] net767 net743 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10258__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09663__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09251_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\] net817 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\]
+ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08202_ _03884_ _03918_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nor3_1
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09182_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\] net754 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\]
+ _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09415__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11758__A0 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08133_ _03842_ _03843_ _03844_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08732__B team_02_WB.instance_to_wrap.top.a1.instruction\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _03706_ _03784_ _03785_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__nor3_2
XFILLER_0_86_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1127_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10733__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\] net696 net677 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15605__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07917_ _03571_ _03600_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_51_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08897_ net29 net1031 net989 team_02_WB.instance_to_wrap.ramload\[5\] vssd1 vssd1
+ vccd1 vccd1 _02533_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout754_A _04375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07848_ _03537_ _03569_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__xor2_2
XFILLER_0_19_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07779_ _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14197__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10249__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09518_ _05020_ _05021_ _05030_ _05034_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__nor4_1
X_10790_ _06304_ _06305_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09654__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\] net759 _04964_ _04965_
+ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a211o_1
XANTENNA__08862__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13232__A2_N net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ net307 net2306 net450 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09406__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08923__A team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11411_ _03294_ net849 vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12391_ net302 net1608 net459 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14130_ net1123 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
X_11342_ net671 _06841_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14061_ net1133 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
X_11273_ _06546_ _06773_ net415 vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__mux2_1
X_13012_ team_02_WB.instance_to_wrap.top.pc\[25\] _06172_ _07531_ vssd1 vssd1 vccd1
+ vccd1 _07532_ sky130_fd_sc_hd__a21oi_1
X_10224_ _05693_ _05740_ net551 vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__mux2_1
XANTENNA_input50_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09754__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10155_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\] net823 net909 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16530__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14963_ net1166 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
X_10086_ _05583_ _05602_ net969 vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__mux2_1
Xhold6 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[4\] vssd1 vssd1 vccd1 vccd1
+ net1464 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16702_ net1440 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_106_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ net1204 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
XANTENNA__10488__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14894_ net1163 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09893__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16633_ clknet_leaf_100_wb_clk_i _02752_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13845_ net1224 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11437__C1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16564_ clknet_leaf_94_wb_clk_i _02688_ _01371_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13776_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] _03269_
+ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10988_ _05954_ _06499_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__and2_1
XANTENNA__09645__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15515_ clknet_leaf_128_wb_clk_i _01655_ _00323_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12727_ _06957_ _07250_ _06915_ _06937_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__nand4b_1
XTAP_TAPCELL_ROW_119_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16495_ clknet_leaf_4_wb_clk_i _02629_ _01302_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15446_ clknet_leaf_64_wb_clk_i _01586_ _00254_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12658_ net304 net2483 net434 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ _05833_ _05998_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15377_ clknet_leaf_78_wb_clk_i _01517_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12589_ net302 net2503 net439 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14328_ net1187 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold406 team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] vssd1 vssd1 vccd1 vccd1
+ net1864 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold417 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16060__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold428 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold439 team_02_WB.instance_to_wrap.ramload\[8\] vssd1 vssd1 vccd1 vccd1 net1897
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14259_ net1165 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08908__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08908__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09030__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_8
Xfanout919 _04515_ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08820_ net1528 net1041 net990 team_02_WB.instance_to_wrap.ramaddr\[11\] vssd1 vssd1
+ vccd1 vccd1 _02605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10191__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ net847 _04368_ _04370_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__and3_4
XFILLER_0_20_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15778__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1139 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07702_ _03422_ _03424_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__nor2_1
X_08682_ net1060 _04308_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nand2_1
XANTENNA__11140__A1 _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09884__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07633_ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] _03339_ _03342_ _03344_ _03355_
+ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__o41a_2
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07564_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 _03304_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_49_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09097__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09636__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09303_ _04816_ _04818_ _04819_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__or3_1
XANTENNA__08844__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16707__1445 vssd1 vssd1 vccd1 vccd1 net1445 _16707__1445/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_135_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13028__B1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1077_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09234_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\] net743 _04749_ _04750_
+ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09839__A _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\] net831 net925 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\]
+ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1244_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08116_ _03832_ _03834_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09096_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\] net734 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ _03725_ _03752_ _03767_ _03768_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_124_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold940 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold951 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold962 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold973 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold984 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout871_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout969_A _04496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12204__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09998_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\] net752 net705 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a22o_1
X_08949_ _04270_ _04273_ _04457_ _04465_ _04309_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13120__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ net304 net2125 net585 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09875__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10911_ _04695_ _05955_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11891_ net298 net1964 net488 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ net1494 net963 _03180_ net1066 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09088__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ net547 net420 vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09627__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ _03289_ net1047 _03113_ _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__and4_2
XANTENNA__08835__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ net609 net403 vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__nand2_1
X_15300_ clknet_leaf_67_wb_clk_i _01444_ _00113_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12512_ net248 net2319 net446 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__mux2_1
X_16280_ clknet_leaf_54_wb_clk_i _02420_ _01088_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input98_A wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ team_02_WB.instance_to_wrap.top.pad.button_control.debounce_dly team_02_WB.instance_to_wrap.top.pad.button_control.debounce
+ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__and2b_2
XFILLER_0_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15231_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[22\]
+ _00044_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_114_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12443_ net244 net2344 net451 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15162_ net1244 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12374_ net346 net2212 net561 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14113_ net1208 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
X_11325_ _05988_ net664 net656 _06825_ _06824_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__o221a_1
XFILLER_0_120_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15093_ net1078 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14044_ net1149 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11256_ _06218_ _06219_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10207_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\] net742 net714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a22o_1
XANTENNA__11519__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15920__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12114__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ net410 _06449_ _06692_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_108_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10138_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\] net784 net701 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\]
+ _05654_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a221o_1
X_15995_ clknet_leaf_127_wb_clk_i _02135_ _00803_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11953__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14946_ net1152 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
X_10069_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\] net916 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09866__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14877_ net1086 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16616_ clknet_leaf_98_wb_clk_i _02735_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13828_ net1252 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
XANTENNA__09079__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09618__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16547_ clknet_leaf_94_wb_clk_i _02671_ _01354_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15300__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ team_02_WB.instance_to_wrap.top.pad.button_control.debounce team_02_WB.instance_to_wrap.top.pad.button_control.noisy
+ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or2_1
XANTENNA__08826__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16426__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16478_ clknet_leaf_74_wb_clk_i net1497 _01286_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15429_ clknet_leaf_33_wb_clk_i _01569_ _00237_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09251__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 _02608_ vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold214 _02580_ vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold225 team_02_WB.instance_to_wrap.ramload\[12\] vssd1 vssd1 vccd1 vccd1 net1683
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold236 team_02_WB.instance_to_wrap.ramaddr\[5\] vssd1 vssd1 vccd1 vccd1 net1694
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] vssd1 vssd1
+ vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold258 _02579_ vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\] net776 _05436_ _05437_
+ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__a211o_1
Xhold269 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout705 _04389_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__buf_4
Xfanout716 net717 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_8
Xfanout727 net729 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_4
X_09852_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\] net829 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\]
+ _05368_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a221o_1
XANTENNA__12024__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout738 _04379_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_6
XANTENNA__10164__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout749 _04377_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_4
X_08803_ net1565 net1042 net992 team_02_WB.instance_to_wrap.ramaddr\[28\] vssd1 vssd1
+ vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
X_09783_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\] net774 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__a22o_1
XANTENNA__11863__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__A _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ net932 vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__and3b_2
XFILLER_0_119_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08738__A team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _03298_ _04278_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout452_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1194_A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] _03338_ vssd1 vssd1 vccd1
+ vccd1 _03339_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_137_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ net56 net55 net58 net57 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__or4_1
XFILLER_0_117_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12613__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08817__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12694__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11416__A2 _06908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09490__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09217_ _04714_ _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13202__A1_N net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09148_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\] net776 net769 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09242__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09079_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\] net887 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11110_ _06174_ _06175_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ net2467 net286 net581 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
Xhold770 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold781 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13217__A1_N _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold792 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net383 _06104_ _06549_ _06531_ _06110_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_9_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10155__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11773__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14800_ net1110 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
X_15780_ clknet_leaf_0_wb_clk_i _01920_ _00588_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12992_ _07476_ _07511_ _07477_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09848__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14731_ net1201 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11943_ net246 net2334 net586 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
XANTENNA__15323__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16449__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11074__A _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14662_ net1072 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11874_ net243 net1650 net488 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
X_16401_ clknet_leaf_64_wb_clk_i _02536_ _01209_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13613_ net1048 _03114_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__or2_1
XANTENNA__08808__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825_ _06337_ _06340_ net366 vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__mux2_1
XANTENNA__11407__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14593_ net1209 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XANTENNA__14385__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16332_ clknet_leaf_24_wb_clk_i _02472_ _01140_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15473__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] _03061_ vssd1 vssd1 vccd1
+ vccd1 _03102_ sky130_fd_sc_hd__or2_1
X_10756_ team_02_WB.instance_to_wrap.top.pc\[31\] _06272_ vssd1 vssd1 vccd1 vccd1
+ _06273_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09481__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16263_ clknet_leaf_29_wb_clk_i _02403_ _01071_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13475_ team_02_WB.START_ADDR_VAL_REG\[15\] net1069 net1003 vssd1 vssd1 vccd1 vccd1
+ net198 sky130_fd_sc_hd__a21o_1
X_10687_ net995 net552 _04417_ _06127_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15214_ clknet_leaf_58_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[5\]
+ _00027_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] sky130_fd_sc_hd__dfrtp_4
X_12426_ net296 net1826 net456 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__mux2_1
XANTENNA__09233__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16194_ clknet_leaf_117_wb_clk_i _02334_ _01002_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11948__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11040__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15145_ net1247 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12357_ net294 net2226 net564 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11308_ team_02_WB.instance_to_wrap.top.pc\[15\] _06261_ team_02_WB.instance_to_wrap.top.pc\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__a21oi_1
X_15076_ net1259 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ net290 net1997 net571 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__mux2_1
X_14027_ net1205 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
X_11239_ net670 _06742_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__nor2_1
XANTENNA__10146__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16706__1444 vssd1 vssd1 vccd1 vccd1 net1444 _16706__1444/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_69_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15978_ clknet_leaf_128_wb_clk_i _02118_ _00786_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13096__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14929_ net1117 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
XANTENNA_wire518_A _05400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10854__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08450_ _04145_ _04153_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_19_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08381_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04070_ vssd1 vssd1 vccd1
+ vccd1 _04091_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09389__A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12359__A0 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12019__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15966__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09002_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ net1056 _04499_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o31a_1
XFILLER_0_2_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09224__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11858__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13358__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09904_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\] net744 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10137__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1207_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\] net778 net698 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\]
+ _05351_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a221o_1
Xfanout557 _07223_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12689__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 _07218_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_6
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_8
XANTENNA_fanout667_A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09766_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\] net927 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\]
+ _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08717_ _04288_ _04320_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__nand2_2
XFILLER_0_94_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09697_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\] net747 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout834_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10845__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ _03298_ team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _04277_ sky130_fd_sc_hd__or2_2
XANTENNA__15496__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08579_ net1719 _04241_ _04225_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__mux2_1
XANTENNA__12598__A0 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10610_ _04283_ _04493_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__and2_2
XFILLER_0_92_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ _05906_ _05910_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ net517 net384 _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_107_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13260_ team_02_WB.instance_to_wrap.top.pc\[28\] net1054 net935 _02977_ vssd1 vssd1
+ vccd1 vccd1 _02978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10472_ _05295_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12211_ net2437 net242 net619 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__mux2_1
XANTENNA__11768__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ _07334_ _07496_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10376__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11573__B2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16121__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ net345 net2300 net467 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13268__B _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13314__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ net360 net2559 net472 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
XANTENNA__12522__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15901_ clknet_leaf_51_wb_clk_i _02041_ _00709_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11024_ _06381_ _06384_ net392 vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16881_ net1425 vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__buf_2
XFILLER_0_102_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12599__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16271__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15832_ clknet_leaf_53_wb_clk_i _01972_ _00640_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13078__A1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15763_ clknet_leaf_53_wb_clk_i _01903_ _00571_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11628__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12975_ _07493_ _07494_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__nor2_1
XANTENNA__12825__A1 _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14714_ net1181 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
X_11926_ net304 net2611 net482 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ clknet_leaf_25_wb_clk_i _01834_ _00502_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10300__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14645_ net1214 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
X_11857_ net297 net2674 net491 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XANTENNA__15989__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10808_ _04802_ net386 vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14576_ net1095 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
X_11788_ net309 net2676 net596 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10064__A1 _05580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16315_ clknet_leaf_126_wb_clk_i _02455_ _01123_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13527_ _03081_ _03082_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__nor2_1
XANTENNA__11251__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10739_ team_02_WB.instance_to_wrap.top.pc\[7\] team_02_WB.instance_to_wrap.top.pc\[6\]
+ _06255_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15219__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16246_ clknet_leaf_47_wb_clk_i _02386_ _01054_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13458_ _02768_ _03047_ _03059_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09206__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12409_ net242 net1953 net457 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__mux2_1
X_16177_ clknet_leaf_21_wb_clk_i _02317_ _00985_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13389_ team_02_WB.instance_to_wrap.ramload\[18\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[18\] sky130_fd_sc_hd__and2_1
XFILLER_0_109_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XANTENNA__10367__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
X_15128_ net1248 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15369__CLK clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13305__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ _03670_ _03672_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__and2_1
X_15059_ net1259 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10119__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire635_A _04860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ net316 _03597_ _03581_ _03584_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__a211o_1
X_09620_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\] net732 _05134_ _05136_
+ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a211o_1
XANTENNA__12302__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09551_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\] net825 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\]
+ _05067_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a221o_1
XANTENNA__11619__A2 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08502_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[8\] net980 vssd1 vssd1 vccd1
+ vccd1 _04196_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09482_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\] net712 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08433_ _04128_ _04130_ _04133_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08735__B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ _04030_ _04053_ _04074_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__nand3_1
XANTENNA__10055__A1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08295_ _03962_ _03988_ _03980_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14753__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13529__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16144__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10358__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout784_A _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16294__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08971__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout310 net311 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_100_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout321 net324 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
Xfanout332 _07013_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_2
Xfanout343 _07051_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_2
Xfanout354 _07087_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout365 net367 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 _06087_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_2
X_09818_ _05314_ _05333_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__or2_2
Xfanout387 _05901_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_2
XANTENNA__12212__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout398 net400 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_55_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09749_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\] net771 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\]
+ _05265_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12760_ _04694_ _05252_ _05335_ _05420_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__or4_1
XFILLER_0_90_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11711_ net265 net2539 net603 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11491__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12691_ net304 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\] net430 vssd1
+ vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11352__A _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14430_ net1191 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
X_11642_ net548 net385 vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09436__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361_ net1136 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11573_ net837 _07057_ _07058_ net669 _07062_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__o221a_1
X_16705__1443 vssd1 vssd1 vccd1 vccd1 net1443 _16705__1443/LO sky130_fd_sc_hd__conb_1
XFILLER_0_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14663__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16100_ clknet_leaf_4_wb_clk_i _02240_ _00908_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13312_ net1722 net986 net967 _03005_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__a22o_1
XANTENNA_input80_A wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10524_ _06039_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14292_ net1077 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16031_ clknet_leaf_86_wb_clk_i _02171_ _00839_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13243_ _06458_ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10455_ _05061_ _05080_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__and2b_1
XANTENNA__10349__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13174_ _07027_ net235 _02933_ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10386_ _05880_ _05902_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08962__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12125_ net294 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\] net467 vssd1
+ vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13299__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15661__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ net274 net2380 net470 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _04783_ _06111_ _06410_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12122__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16864_ net1408 vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15815_ clknet_leaf_27_wb_clk_i _01955_ _00623_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16017__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16795_ net1339 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_137_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11961__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15746_ clknet_leaf_123_wb_clk_i _01886_ _00554_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12958_ _07477_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__inv_2
XANTENNA__09675__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11909_ net244 net2602 net483 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15677_ clknet_leaf_51_wb_clk_i _01817_ _00485_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12889_ _07407_ _07408_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14628_ net1129 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14559_ net1190 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08080_ _03795_ _03800_ _03790_ _03792_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_114_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16229_ clknet_leaf_30_wb_clk_i _02369_ _01037_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08938__C1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08982_ _04275_ _04310_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07933_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__inv_2
XANTENNA__09902__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ _03571_ _03574_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__nand2b_2
XANTENNA__12032__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09603_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\] net811 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\]
+ _05119_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a221o_1
X_07795_ _03465_ _03474_ net364 _03488_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11871__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09534_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\] net778 net734 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a22o_1
XANTENNA__13462__A1 team_02_WB.START_ADDR_VAL_REG\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09130__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09465_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\] _04529_ _04530_
+ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\] _04981_ vssd1 vssd1 vccd1
+ vccd1 _04982_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08416_ _04104_ _04115_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__and2b_1
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09418__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\] net771 net731 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08347_ _04047_ _04058_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_102_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08278_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] _03989_ vssd1 vssd1 vccd1
+ vccd1 _03993_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout999_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12207__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10240_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\] net908 _05743_ _05756_
+ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a211o_1
XANTENNA__15684__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10736__C1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\] net836 net917 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\]
+ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_110_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1105 net1107 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_4
Xfanout1116 net1125 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__clkbuf_4
Xfanout1127 net1135 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_4
Xfanout1138 net1144 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_4
Xfanout1149 net1153 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__buf_4
X_13930_ net1218 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11700__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13861_ net1226 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15600_ clknet_leaf_39_wb_clk_i _01740_ _00408_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11781__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ net231 _07334_ _07335_ _07329_ _04280_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a32o_1
XFILLER_0_134_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16580_ clknet_leaf_95_wb_clk_i _02699_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13792_ _03280_ _03281_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__nor2_1
XANTENNA__09657__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09121__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15531_ clknet_leaf_112_wb_clk_i _01671_ _00339_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10267__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ _06728_ _06754_ _07266_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__nand3_1
XFILLER_0_57_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ clknet_leaf_49_wb_clk_i _01602_ _00270_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12674_ net246 net2081 net430 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10019__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14413_ net1141 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
X_11625_ net422 _06776_ _07111_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15393_ clknet_leaf_121_wb_clk_i _01533_ _00201_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14344_ net1177 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire530 net531 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire541 _04754_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__dlymetal6s2s_1
X_11556_ team_02_WB.instance_to_wrap.top.pc\[5\] _06254_ vssd1 vssd1 vccd1 vccd1 _07047_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10507_ _05972_ _05976_ _06023_ _06020_ _05977_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__o32a_1
XANTENNA__12117__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14275_ net1133 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11487_ net376 _06796_ _06980_ net381 vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16014_ clknet_leaf_9_wb_clk_i _02154_ _00822_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13226_ net649 net936 net1020 net1596 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09188__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10438_ _04779_ _05954_ _04734_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_1674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11956__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13157_ _06972_ net232 _02921_ net977 _02919_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10369_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\] net876 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a22o_1
XANTENNA_max_cap428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ net1922 net347 net581 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux2_1
X_13088_ _07365_ _07426_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12039_ net363 net1884 net477 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__mux2_1
XANTENNA__15407__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09360__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16847_ net1391 vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07580_ net1883 net1063 net37 vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a21o_1
X_16778_ net1322 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XANTENNA__09648__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09112__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15557__CLK clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15729_ clknet_leaf_23_wb_clk_i _01869_ _00537_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_115_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09250_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\] net927 net912 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08201_ _03886_ _03898_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__xor2_4
XFILLER_0_51_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\] net782 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08132_ _03850_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_133_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09820__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ _03711_ _03753_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12027__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09179__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16799__1343 vssd1 vssd1 vccd1 vccd1 _16799__1343/HI net1343 sky130_fd_sc_hd__conb_1
XANTENNA__11866__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1022_A _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10194__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__C1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08965_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\] net748 _04473_ _04475_
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_122_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout482_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07916_ _03605_ _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08896_ net30 net1029 net987 net1771 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__o22a_1
X_16704__1442 vssd1 vssd1 vccd1 vccd1 net1442 _16704__1442/LO sky130_fd_sc_hd__conb_1
XANTENNA__09887__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09860__A _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ _03537_ _03551_ net329 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12697__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14478__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07778_ _03467_ _03500_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09517_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\] net868 _05031_ _05033_
+ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__a211o_1
XANTENNA__09103__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16755__1299 vssd1 vssd1 vccd1 vccd1 _16755__1299/HI net1299 sky130_fd_sc_hd__conb_1
XFILLER_0_52_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout914_A _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09448_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\] net787 net755 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a22o_1
X_09379_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\] net805 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\]
+ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08923__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15102__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ net671 _06893_ _06907_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08614__A1 team_02_WB.START_ADDR_VAL_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12390_ net294 net2014 net460 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11341_ _05294_ _06015_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_112_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14060_ net1080 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11272_ net420 _06774_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13011_ _07530_ _07454_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__and2b_1
XANTENNA__11776__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] net650 _05739_ vssd1
+ vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10185__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input43_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10154_ team_02_WB.instance_to_wrap.top.a1.instruction\[26\] net792 _05670_ vssd1
+ vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09590__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14962_ net1122 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
X_10085_ _05594_ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__or2_2
Xhold7 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[8\] vssd1 vssd1 vccd1 vccd1
+ net1465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09878__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ net1439 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
X_13913_ net1218 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10488__B2 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14893_ net1140 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
X_13844_ net1217 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
X_16632_ clknet_leaf_100_wb_clk_i _02751_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12400__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13775_ _03269_ _03270_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16563_ clknet_leaf_94_wb_clk_i _02687_ _01370_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10987_ _04783_ _05953_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12726_ _06976_ _07014_ _07249_ _06995_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__and4bb_1
X_15514_ clknet_leaf_120_wb_clk_i _01654_ _00322_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16494_ clknet_leaf_35_wb_clk_i _02628_ _01301_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15445_ clknet_leaf_40_wb_clk_i _01585_ _00253_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12657_ net298 net2201 net435 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ net795 _07094_ _06117_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ clknet_leaf_78_wb_clk_i _01516_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__09802__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ net293 net2352 net439 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14327_ net1172 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
XANTENNA__16205__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11539_ net2082 net337 net643 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold407 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold418 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14258_ net1123 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold429 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13209_ net2036 net1020 net938 _04904_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14189_ net1141 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
Xfanout909 _04524_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__buf_4
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16355__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire548_A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1107 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
X_08750_ net847 _04360_ _04365_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__and3_2
Xhold1118 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1129 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09869__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07701_ _03383_ _03423_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__xor2_1
XANTENNA__09333__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08681_ net1062 net1060 _04266_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08541__B1 _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ _03328_ _03346_ _03352_ team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] team_02_WB.instance_to_wrap.top.a1.dataIn\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_90_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12310__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07563_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 _03303_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09302_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\] net899 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\]
+ _04808_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10100__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\] net783 net747 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout230_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout328_A _06975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09164_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\] net908 net897 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08115_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09095_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\] net678 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1237_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ _03744_ _03750_ _03766_ _03725_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold930 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold941 team_02_WB.instance_to_wrap.top.a1.row1\[58\] vssd1 vssd1 vccd1 vccd1 net2399
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold952 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold963 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold974 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\] vssd1
+ vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold985 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12712__C _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold996 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09572__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09997_ _05489_ _05511_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout864_A _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ _04310_ _04316_ _04317_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ net17 net1030 net988 net2259 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10910_ net1923 net239 net642 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__mux2_1
XANTENNA__12220__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ net309 net2736 net489 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10841_ _06355_ _06356_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13840__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13560_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__nor2_2
X_10772_ _06286_ _06287_ net389 vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12511_ net251 net2444 net448 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13491_ team_02_WB.START_ADDR_VAL_REG\[31\] net1070 net1004 vssd1 vssd1 vccd1 vccd1
+ net216 sky130_fd_sc_hd__a21o_1
XFILLER_0_82_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15230_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[21\]
+ _00043_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12442_ net241 net1847 net452 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15161_ net1243 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12373_ net350 net2423 net564 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__mux2_1
XANTENNA__15252__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14112_ net1158 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11324_ _06358_ _06821_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__or2_1
X_15092_ net1104 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14043_ net1157 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
X_11255_ _06743_ _06756_ _06758_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__or3b_2
XANTENNA__10158__B1 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10206_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\] net782 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\]
+ _05722_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__a221o_1
XANTENNA__09563__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11186_ net411 _06691_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10137_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\] net748 net677 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__a22o_1
X_15994_ clknet_leaf_120_wb_clk_i _02134_ _00802_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09315__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\] net811 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__a22o_1
X_14945_ net1211 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12130__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10330__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14876_ net1150 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16615_ clknet_leaf_99_wb_clk_i _02734_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13827_ net1232 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16798__1342 vssd1 vssd1 vccd1 vccd1 _16798__1342/HI net1342 sky130_fd_sc_hd__conb_1
X_13758_ team_02_WB.instance_to_wrap.top.pad.button_control.debounce team_02_WB.instance_to_wrap.top.pad.button_control.noisy
+ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16546_ clknet_leaf_94_wb_clk_i _02670_ _01353_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ _04325_ _04355_ _06162_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__or3_1
XANTENNA__11830__A0 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13689_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\]
+ _03200_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_14_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16477_ clknet_leaf_89_wb_clk_i net1501 _01285_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_14_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08563__B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13293__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15428_ clknet_leaf_0_wb_clk_i _01568_ _00236_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire498_A _05828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16703__1441 vssd1 vssd1 vccd1 vccd1 net1441 _16703__1441/LO sky130_fd_sc_hd__conb_1
XFILLER_0_53_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15359_ clknet_leaf_90_wb_clk_i _01499_ _00172_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14581__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold204 team_02_WB.instance_to_wrap.top.a1.row1\[121\] vssd1 vssd1 vccd1 vccd1 net1662
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold215 team_02_WB.instance_to_wrap.top.a1.row1\[109\] vssd1 vssd1 vccd1 vccd1 net1673
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 team_02_WB.instance_to_wrap.ramstore\[29\] vssd1 vssd1 vccd1 vccd1 net1684
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold237 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1
+ net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold248 team_02_WB.instance_to_wrap.ramaddr\[26\] vssd1 vssd1 vccd1 vccd1 net1706
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\] net704 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a22o_1
Xhold259 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15745__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12305__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10614__A _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16754__1298 vssd1 vssd1 vccd1 vccd1 _16754__1298/HI net1298 sky130_fd_sc_hd__conb_1
XFILLER_0_46_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout706 _04387_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout717 _04385_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_4
X_09851_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\] net833 net821 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__a22o_1
Xfanout728 net729 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _04379_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__clkbuf_4
X_08802_ net1503 net1043 net993 team_02_WB.instance_to_wrap.ramaddr\[29\] vssd1 vssd1
+ vccd1 vccd1 _02623_ sky130_fd_sc_hd__a22o_1
X_09782_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\] net758 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\]
+ _05296_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15895__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ _04358_ _04360_ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08664_ _04291_ _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__nor2_1
XANTENNA__12040__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07615_ _03324_ _03328_ _03325_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_137_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ net63 net62 net59 net60 vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_137_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1187_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09216_ net971 net637 net544 vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_134_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09147_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\] net785 net761 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_92_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\] net833 net926 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\]
+ _04594_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09793__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout981_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _03744_ _03750_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12215__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold760 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 team_02_WB.instance_to_wrap.top.ru.state\[0\] vssd1 vssd1 vccd1 vccd1 net2229
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold782 team_02_WB.instance_to_wrap.top.a1.row2\[40\] vssd1 vssd1 vccd1 vccd1 net2240
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09545__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _05951_ net662 net659 _04823_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__a22o_1
Xhold793 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13835__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12991_ team_02_WB.instance_to_wrap.top.pc\[11\] _05445_ _07510_ vssd1 vssd1 vccd1
+ vccd1 _07511_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11942_ net241 net1974 net588 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__mux2_1
X_14730_ net1142 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14661_ net1085 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
X_11873_ net647 _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__nand2_4
XANTENNA__16050__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16400_ clknet_leaf_65_wb_clk_i _02535_ _01208_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13612_ _03160_ _03163_ _03108_ _03135_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_131_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824_ _06338_ _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__or2_1
XANTENNA__15618__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14592_ net1158 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
XANTENNA__08808__B2 team_02_WB.instance_to_wrap.ramaddr\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11812__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13543_ team_02_WB.instance_to_wrap.top.edg2.button_i _03090_ _03099_ _03100_ vssd1
+ vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__or4_1
X_16331_ clknet_leaf_112_wb_clk_i _02471_ _01139_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10755_ team_02_WB.instance_to_wrap.top.pc\[30\] _06271_ vssd1 vssd1 vccd1 vccd1
+ _06272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16262_ clknet_leaf_44_wb_clk_i _02402_ _01070_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10091__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13474_ team_02_WB.START_ADDR_VAL_REG\[14\] _04260_ vssd1 vssd1 vccd1 vccd1 net197
+ sky130_fd_sc_hd__and2_1
XFILLER_0_10_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10686_ _06201_ _06202_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15213_ clknet_leaf_58_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[4\]
+ _00026_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] sky130_fd_sc_hd__dfrtp_4
X_12425_ net308 net2445 net457 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15768__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16193_ clknet_leaf_117_wb_clk_i _02333_ _01001_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10379__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15144_ net1245 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12356_ net285 net2407 net563 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__mux2_1
XANTENNA__09784__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13317__B1 _07122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ _06214_ _06808_ net974 vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__and3b_1
XFILLER_0_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15075_ net1256 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10434__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12125__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ net276 net1972 net569 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14026_ net1168 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
XANTENNA__09536__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ _05127_ _06597_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__xor2_1
XANTENNA__11964__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11169_ _06355_ _06674_ _06123_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07743__A team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15977_ clknet_leaf_104_wb_clk_i _02117_ _00785_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13096__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14928_ net1109 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
XANTENNA__10303__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14859_ net1205 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ _04087_ _04089_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16529_ clknet_leaf_60_wb_clk_i _00006_ _01336_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08275__A2 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10082__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09001_ _04516_ _04517_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__nor2_4
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15200__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12035__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09527__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09903_ net517 _05419_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11874__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_127_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09834_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\] net754 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__a22o_1
Xfanout547 _04489_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_2
XFILLER_0_67_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout558 _07223_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1102_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout569 _07217_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_8
X_09765_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\] net923 net875 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout562_A _07219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08716_ net1059 _04286_ _04316_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__or3b_1
XFILLER_0_55_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09696_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\] net780 net733 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09160__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08647_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] net997 vssd1 vssd1 vccd1
+ vccd1 _04276_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_29_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13390__A team_02_WB.instance_to_wrap.ramload\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _02811_ _04230_ _04227_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__o21a_1
XANTENNA__08484__A _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10519__A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15910__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10540_ net515 net402 vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__nand2_1
XANTENNA__10073__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10953__S net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ _05252_ _05937_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__nand2_2
XFILLER_0_134_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12210_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04291_ _04292_ _04333_
+ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__nor4_1
XANTENNA__15110__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09766__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13190_ team_02_WB.instance_to_wrap.top.pc\[3\] net1023 _02948_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01484_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12141_ net348 net2346 net468 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16797__1341 vssd1 vssd1 vccd1 vccd1 _16797__1341/HI net1341 sky130_fd_sc_hd__conb_1
X_12072_ net352 net2719 net472 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
Xhold590 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11784__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15900_ clknet_leaf_45_wb_clk_i _02040_ _00708_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11023_ net407 _06377_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__or2_1
X_16880_ net1424 vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__buf_2
XFILLER_0_95_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07563__A team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15831_ clknet_leaf_13_wb_clk_i _01971_ _00639_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11085__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16702__1440 vssd1 vssd1 vccd1 vccd1 net1440 _16702__1440/LO sky130_fd_sc_hd__conb_1
XFILLER_0_73_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15762_ clknet_leaf_9_wb_clk_i _01902_ _00570_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12974_ team_02_WB.instance_to_wrap.top.pc\[3\] _05787_ vssd1 vssd1 vccd1 vccd1 _07494_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__15440__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1290 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09151__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14713_ net1137 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
X_11925_ net296 net2433 net483 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
X_15693_ clknet_leaf_24_wb_clk_i _01833_ _00501_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11856_ net310 net2478 net493 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
X_14644_ net1090 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
X_16753__1297 vssd1 vssd1 vccd1 vccd1 _16753__1297/HI net1297 sky130_fd_sc_hd__conb_1
XFILLER_0_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ _06322_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14575_ net1121 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
XANTENNA__15590__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11787_ net301 net2558 net594 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13250__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16314_ clknet_leaf_117_wb_clk_i _02454_ _01122_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11261__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13526_ _03075_ _03086_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__nor2_1
X_10738_ team_02_WB.instance_to_wrap.top.pc\[5\] _06254_ vssd1 vssd1 vccd1 vccd1 _06255_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_137_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11959__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16245_ clknet_leaf_43_wb_clk_i _02385_ _01053_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13457_ _03056_ _03059_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__nand2_1
X_10669_ _06128_ _06185_ _04490_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__a21oi_4
XANTENNA__13002__A2 _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12408_ net645 _07197_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09757__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16176_ clknet_leaf_39_wb_clk_i _02316_ _00984_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13388_ team_02_WB.instance_to_wrap.ramload\[17\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[17\] sky130_fd_sc_hd__and2_1
XFILLER_0_3_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12339_ net362 net2374 net567 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__mux2_1
X_15127_ net1248 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15058_ net1259 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
XANTENNA__09509__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14009_ net1128 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
X_07880_ _03581_ _03598_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire530_A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire628_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\] net866 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_95_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13201__A1_N _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09142__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ net1046 _04185_ _04194_ _04195_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__a31o_1
XANTENNA__10827__A1 _05715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\] net780 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15933__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08432_ _04119_ _04131_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08735__C team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ _04060_ _04063_ _04067_ _04070_ _04066_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__a41o_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08595__D_N net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10055__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__B2 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ _03980_ _03990_ _04003_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11869__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout310_A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1052_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09748__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13369__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15313__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout300 net303 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_2
Xfanout311 _06840_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_2
Xfanout322 net324 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout333 net336 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10515__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 _07087_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_1
XANTENNA__08479__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout366 net367 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09381__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout377 net380 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_2
XANTENNA__09920__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09817_ _05333_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__inv_2
Xfanout388 net391 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_2
XANTENNA__16696__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12268__A0 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\] net751 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09679_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\] net915 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11710_ net256 net1872 net604 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_95_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15105__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10294__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ net297 net2708 net431 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11641_ net377 _06567_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14944__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14360_ net1220 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10046__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ net666 net377 _06432_ _07061_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09987__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11779__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13311_ team_02_WB.instance_to_wrap.top.pc\[4\] net1052 _07064_ net933 vssd1 vssd1
+ vccd1 vccd1 _03005_ sky130_fd_sc_hd__a22o_2
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_1
X_10523_ _05782_ net403 vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14291_ net1172 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
XANTENNA__08178__A1_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13242_ _06490_ _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__nor2_1
X_16030_ clknet_leaf_112_wb_clk_i _02170_ _00838_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09739__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input73_A wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _04802_ _04822_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08947__B1 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13173_ net977 _07403_ _02934_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__or3_1
X_10385_ net548 net385 vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12124_ net285 net1841 net467 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13299__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12055_ net290 net2016 net472 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__mux2_1
XANTENNA__12403__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ net383 _06513_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__nand2_1
XANTENNA__09372__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16863_ net1407 vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__buf_2
XFILLER_0_99_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09911__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11019__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15814_ clknet_leaf_44_wb_clk_i _01954_ _00622_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_16794_ net1338 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XANTENNA__09124__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15745_ clknet_leaf_121_wb_clk_i _01885_ _00553_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12957_ _03294_ _07378_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11908_ net243 net1819 net484 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__mux2_1
XANTENNA__10285__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15676_ clknet_leaf_44_wb_clk_i _01816_ _00484_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12888_ _05533_ _05536_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09013__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14627_ net1145 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
X_11839_ net647 _07195_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__nand2_8
X_16709__1268 vssd1 vssd1 vccd1 vccd1 _16709__1268/HI net1268 sky130_fd_sc_hd__conb_1
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13223__A2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10037__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11234__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09948__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09978__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14558_ net1194 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15336__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13509_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\] _03066_
+ _03067_ _03070_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__or4_1
XFILLER_0_86_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14489_ net1129 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16228_ clknet_leaf_0_wb_clk_i _02368_ _01036_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11537__A2 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16159_ clknet_leaf_111_wb_clk_i _02299_ _00967_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15486__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08981_ _04494_ net972 vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__nand2_1
X_07932_ _03613_ _03636_ _03653_ _03654_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__a22o_1
XANTENNA__12313__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07863_ _03578_ _03580_ _03583_ _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__o211a_2
XANTENNA__09902__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09602_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\] net924 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a22o_1
X_07794_ _03515_ _03516_ _03513_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__o21a_1
XANTENNA__09115__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09533_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\] net702 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\]
+ _05049_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout260_A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10276__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\] net895 net939 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16111__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08415_ _04113_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__and2_1
X_09395_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\] net707 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__a22o_1
X_16796__1340 vssd1 vssd1 vccd1 vccd1 _16796__1340/HI net1340 sky130_fd_sc_hd__conb_1
XFILLER_0_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08346_ _04058_ _03321_ net1006 net1809 vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10028__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09969__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11599__S net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ _03988_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15829__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout894_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10736__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10200__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10170_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\] net897 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_110_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_4
XFILLER_0_101_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12489__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1117 net1120 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__buf_4
X_16752__1296 vssd1 vssd1 vccd1 vccd1 _16752__1296/HI net1296 sky130_fd_sc_hd__conb_1
XANTENNA__10532__A _05579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12223__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1135 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__buf_4
Xfanout1139 net1144 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09354__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13843__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__A2 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13860_ net1231 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12811_ team_02_WB.instance_to_wrap.top.pc\[1\] _04422_ vssd1 vssd1 vccd1 vccd1 _07335_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__11448__A2_N net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ net1888 _03278_ net960 vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ clknet_leaf_1_wb_clk_i _01670_ _00338_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12742_ _06776_ _06797_ net418 vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15461_ clknet_leaf_33_wb_clk_i _01601_ _00269_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12673_ net241 net1742 net433 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14412_ net1080 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
X_11624_ net378 _07108_ _07110_ net373 _06961_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__o32a_1
X_15392_ clknet_leaf_118_wb_clk_i _01532_ _00200_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14343_ net1117 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
X_11555_ net669 _07031_ _07045_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__o21ai_4
Xwire520 _05313_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire531 _05102_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10506_ _05124_ _05973_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__nor2_1
X_14274_ net1207 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11486_ _06897_ _06979_ net395 vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16013_ clknet_leaf_32_wb_clk_i _02153_ _00821_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13225_ net1602 net1018 net938 _05602_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10437_ _04783_ _05953_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12922__A _04489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09593__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ _07410_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08611__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10368_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\] _04529_ net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12107_ net2193 net348 net584 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12133__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ _07522_ _02862_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__xnor2_1
X_10299_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\] net788 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\]
+ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__a221o_1
XANTENNA__13141__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ net352 net2589 net475 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16846_ net1390 vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_2
XFILLER_0_79_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16134__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09648__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16777_ net1321 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
X_13989_ net1126 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15728_ clknet_leaf_33_wb_clk_i _01868_ _00536_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10258__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16284__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15659_ clknet_leaf_114_wb_clk_i _01799_ _00467_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14584__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08200_ _03865_ _03906_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09180_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\] net786 net738 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08131_ _03809_ _03817_ _03814_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12308__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08062_ _03758_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__xor2_4
XFILLER_0_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08964_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\] net725 _04477_ _04478_
+ _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_55_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13132__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07915_ _03615_ _03618_ _03635_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__a21oi_1
X_08895_ net31 net1029 net987 net1948 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11882__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A _07206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07846_ _03551_ net329 vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07777_ _03473_ net364 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout642_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15501__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09516_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\] net815 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\]
+ _05032_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09447_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\] net727 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout907_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09378_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\] net813 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a22o_1
XANTENNA__15651__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08329_ _04035_ _04040_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nand2_1
XANTENNA__12218__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11340_ net2039 net308 net641 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11271_ _06550_ _06773_ net414 vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13010_ _07455_ _07529_ _07456_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__o21ai_1
X_10222_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\] net997 _04329_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a22o_1
XANTENNA__09575__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11358__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _05625_ _05668_ net551 vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__mux2_1
XANTENNA__16157__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16708__1267 vssd1 vssd1 vccd1 vccd1 _16708__1267/HI net1267 sky130_fd_sc_hd__conb_1
XFILLER_0_41_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09327__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ net1105 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
XANTENNA_input36_A gpio_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ _05597_ _05598_ _05600_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__or3_1
XANTENNA__11792__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[0\] vssd1 vssd1 vccd1 vccd1
+ net1466 sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ net1438 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13912_ net1218 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11685__A1 _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08667__A team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14892_ net1082 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16631_ clknet_leaf_100_wb_clk_i _02750_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13843_ net1224 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13426__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16562_ clknet_leaf_96_wb_clk_i _02686_ _01369_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11437__B2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13774_ net2070 _03267_ net960 vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__o21ai_1
X_10986_ net2033 net248 net642 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15513_ clknet_leaf_112_wb_clk_i _01653_ _00321_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12725_ _07248_ _07058_ _07031_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__and3b_1
XFILLER_0_128_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16493_ clknet_leaf_83_wb_clk_i _02627_ _01300_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08853__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15444_ clknet_leaf_11_wb_clk_i _01584_ _00252_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ net309 net2411 net435 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ net422 _06750_ _07092_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08066__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12128__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15375_ clknet_leaf_78_wb_clk_i _01515_ _00188_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_12587_ net286 net2585 net440 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14326_ net1094 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11538_ net947 _07026_ _07029_ net607 vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11967__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold408 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14257_ net1106 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
XANTENNA__10871__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11469_ _06547_ _06853_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13208_ net635 net936 net1021 net1763 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07746__A team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09030__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14188_ net1071 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ team_02_WB.instance_to_wrap.top.pc\[12\] net1023 _02906_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01493_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13186__C _07394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09318__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13114__A1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14579__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07700_ _03351_ _03386_ _03411_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08680_ net1062 _04266_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__nand2_4
XFILLER_0_20_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire610_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] _03353_ vssd1 vssd1 vccd1
+ vccd1 _03354_ sky130_fd_sc_hd__xor2_1
X_16829_ net1373 vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__buf_2
XFILLER_0_71_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11207__S net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07562_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 _03302_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_88_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11428__A1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15674__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09097__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09301_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\] net834 net894 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\]
+ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08844__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09232_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\] net786 net738 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16751__1295 vssd1 vssd1 vccd1 vccd1 _16751__1295/HI net1295 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_44_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09163_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\] net808 net869 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\]
+ _04679_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12038__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08114_ _03795_ _03818_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_20_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09094_ _04609_ _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_86_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11877__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08045_ _03725_ _03766_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold920 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold931 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold942 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold953 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold964 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold975 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11364__B1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold986 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold997 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09996_ _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__inv_2
XANTENNA__09309__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08947_ _04318_ _04339_ _04309_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout857_A _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13393__A team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__A1 _05440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11667__B2 _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ net18 net1032 net989 net2599 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07829_ _03532_ _03533_ _03511_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_101_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10840_ net546 net415 vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__or2_2
XFILLER_0_67_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09088__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10771_ net548 net403 vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__nor2_1
XANTENNA__08835__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__B _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ net239 net1835 net446 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__mux2_1
XANTENNA__15113__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13490_ team_02_WB.START_ADDR_VAL_REG\[30\] net1069 net1004 vssd1 vssd1 vccd1 vccd1
+ net215 sky130_fd_sc_hd__a21o_1
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12441_ net645 _07199_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15160_ net1249 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
X_12372_ net360 net2596 net563 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14111_ net1182 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
XANTENNA__11787__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11323_ _05252_ net658 _06113_ _05937_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_133_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15091_ net1104 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09548__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07566__A team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14042_ net1182 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
X_11254_ net838 _06741_ _06751_ net657 _06757_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10205_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\] net843 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a22o_1
XANTENNA__15547__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11185_ _06578_ _06690_ net398 vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\] net756 net737 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16775__1319 vssd1 vssd1 vccd1 vccd1 _16775__1319/HI net1319 sky130_fd_sc_hd__conb_1
X_15993_ clknet_leaf_112_wb_clk_i _02133_ _00801_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10067_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\] net896 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__a22o_1
X_14944_ net1158 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
XANTENNA__12411__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15697__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09720__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14875_ net1159 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16614_ clknet_leaf_79_wb_clk_i _02733_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13826_ net1232 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09079__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16545_ clknet_leaf_94_wb_clk_i _02669_ _01352_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13757_ _03256_ _03257_ _03066_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13280__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ net417 _06481_ _06355_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_46_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10094__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12708_ _06124_ _07231_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__nor2_1
X_16476_ clknet_leaf_72_wb_clk_i net1773 _01284_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\] _03200_ net1686 vssd1 vssd1
+ vccd1 vccd1 _03215_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_14_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15427_ clknet_leaf_124_wb_clk_i _01567_ _00235_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12639_ net645 _07210_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09787__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15358_ clknet_leaf_90_wb_clk_i _01498_ _00171_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09251__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold205 team_02_WB.instance_to_wrap.ramstore\[13\] vssd1 vssd1 vccd1 vccd1 net1663
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14309_ net1086 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold216 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ clknet_leaf_78_wb_clk_i _01433_ _00102_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold227 team_02_WB.instance_to_wrap.top.pad.button_control.noisy vssd1 vssd1 vccd1
+ vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09539__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold238 _02762_ vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 team_02_WB.instance_to_wrap.ramaddr\[25\] vssd1 vssd1 vccd1 vccd1 net1707
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16472__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 _04387_ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_4
X_09850_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\] net817 net886 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\]
+ _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a221o_1
Xfanout718 _04384_ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 _04382_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ net1600 net1042 net992 team_02_WB.instance_to_wrap.ramaddr\[30\] vssd1 vssd1
+ vccd1 vccd1 _02624_ sky130_fd_sc_hd__a22o_1
XANTENNA__09691__A _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09781_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\] net754 net698 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\]
+ _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13417__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08732_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__and3_1
XANTENNA__12321__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09711__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08663_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__nand2_2
XFILLER_0_59_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07614_ _03326_ _03330_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__and2_1
X_08594_ net46 net49 net48 net47 vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_137_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13271__B1 _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout340_A _07030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08817__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1082_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout438_A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09490__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09215_ _04725_ _04728_ _04730_ _04731_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__nor4_2
XFILLER_0_118_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout605_A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09146_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\] net709 net685 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_92_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09242__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13388__A team_02_WB.instance_to_wrap.ramload\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09077_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\] net826 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10805__A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08028_ _03744_ _03750_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold750 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold761 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold794 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09979_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\] net815 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\]
+ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__a221o_1
XANTENNA__11636__A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10540__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ _07481_ _07509_ _07479_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__o21a_1
XANTENNA__08505__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09702__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11941_ _04292_ net645 _07201_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__or3_4
XFILLER_0_93_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13851__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14660_ net1130 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11872_ _07190_ _07193_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__nor2_1
XANTENNA__08945__A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13611_ _03117_ _03161_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10823_ _04928_ net405 vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13262__B1 _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14591_ net1193 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
XANTENNA__08808__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ clknet_leaf_128_wb_clk_i _02470_ _01138_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10076__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13542_ _03078_ _03081_ _03072_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a21oi_1
X_10754_ team_02_WB.instance_to_wrap.top.pc\[29\] _06270_ vssd1 vssd1 vccd1 vccd1
+ _06271_ sky130_fd_sc_hd__and2_1
XANTENNA__16345__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09481__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ clknet_leaf_31_wb_clk_i _02401_ _01069_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13473_ team_02_WB.START_ADDR_VAL_REG\[13\] net1068 net1002 vssd1 vssd1 vccd1 vccd1
+ net196 sky130_fd_sc_hd__a21o_1
X_10685_ team_02_WB.instance_to_wrap.top.pc\[13\] _06200_ vssd1 vssd1 vccd1 vccd1
+ _06202_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09769__B1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15212_ clknet_leaf_58_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[3\]
+ _00025_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12424_ net301 net2582 net456 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__mux2_1
XANTENNA__09776__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16192_ clknet_leaf_109_wb_clk_i _02332_ _01000_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09233__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15143_ net1245 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12406__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ net272 net2704 net561 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__mux2_1
XANTENNA__11040__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13317__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _06195_ _06212_ _06213_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__nand3_1
X_15074_ net1259 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
X_12286_ net280 net2413 net570 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14025_ net1101 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
X_11237_ _05127_ _05943_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10000__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ _04996_ net665 _06667_ net796 _06668_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__o221a_1
X_16750__1294 vssd1 vssd1 vccd1 vccd1 _16750__1294/HI net1294 sky130_fd_sc_hd__conb_1
XFILLER_0_93_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10119_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\] net816 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\]
+ _05630_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12141__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099_ net415 _06107_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__or2_1
XANTENNA__10450__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ clknet_leaf_19_wb_clk_i _02116_ _00784_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14927_ net1165 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11980__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10854__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14858_ net1142 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13809_ net1228 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13253__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14789_ net1094 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10067__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16528_ clknet_leaf_70_wb_clk_i _00005_ _01335_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_85_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16459_ clknet_leaf_74_wb_clk_i net1487 _01267_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14592__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09000_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ _04499_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09224__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12316__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10625__A team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13308__B2 _03003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ net970 net625 net543 vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_35_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12840__A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09932__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09833_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\] net786 net718 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\]
+ _05349_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__a221o_1
Xfanout559 _07223_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__buf_6
XANTENNA__08999__C_N net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\] net806 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\]
+ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__a221o_1
XANTENNA__10360__A _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08715_ _04338_ _04340_ _04341_ _04343_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__and4b_1
X_09695_ _05207_ _05209_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11890__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout555_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08646_ _04265_ net1062 net1060 vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_90_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16368__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout722_A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ net1774 _04240_ _04225_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09999__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16774__1318 vssd1 vssd1 vccd1 vccd1 _16774__1318/HI net1318 sky130_fd_sc_hd__conb_1
XFILLER_0_8_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10470_ _05231_ _05251_ _05291_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a21o_1
XANTENNA__11558__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09129_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\] net906 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\]
+ _04645_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12226__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10230__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ net362 net2029 net468 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
XANTENNA__08005__A team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12071_ net357 net2626 net470 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold580 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold591 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _06531_ _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__xnor2_1
X_15830_ clknet_leaf_62_wb_clk_i _01970_ _00638_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15761_ clknet_leaf_21_wb_clk_i _01901_ _00569_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12973_ team_02_WB.instance_to_wrap.top.pc\[3\] _05787_ vssd1 vssd1 vccd1 vccd1 _07493_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_77_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1280 team_02_WB.instance_to_wrap.top.pad.keyCode\[5\] vssd1 vssd1 vccd1 vccd1
+ net2738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ net1215 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10297__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11924_ net310 net2235 net485 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__mux2_1
X_15692_ clknet_leaf_25_wb_clk_i _01832_ _00500_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ net1164 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ net301 net2567 net491 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XANTENNA__15735__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10049__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10806_ _06320_ _06321_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nor2_1
X_14574_ net1164 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
XANTENNA__11797__A0 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11786_ net292 net2059 net593 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16313_ clknet_leaf_17_wb_clk_i _02453_ _01121_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13525_ team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__or4b_1
XFILLER_0_32_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10737_ team_02_WB.instance_to_wrap.top.pc\[4\] team_02_WB.instance_to_wrap.top.pc\[3\]
+ team_02_WB.instance_to_wrap.top.pc\[2\] vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16244_ clknet_leaf_11_wb_clk_i _02384_ _01052_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15885__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13456_ _03038_ _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_58_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10668_ net994 _05580_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__nand2_1
XANTENNA__08614__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09206__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ net345 net2241 net458 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__mux2_1
X_16175_ clknet_leaf_38_wb_clk_i _02315_ _00983_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12136__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13387_ net2759 net1011 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[16\]
+ sky130_fd_sc_hd__and2_1
X_10599_ _04462_ _06114_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__or2_4
XANTENNA__10445__A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
X_15126_ net1227 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_84_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12338_ net352 net2648 net567 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15057_ net1263 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12269_ net339 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\] net576 vssd1
+ vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14008_ net1187 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
XANTENNA__09914__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15265__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire523_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15959_ clknet_leaf_14_wb_clk_i _02099_ _00767_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08500_ net2745 net850 vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__and2_1
XANTENNA__10827__A2 _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09480_ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08431_ _04119_ _04131_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16660__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08362_ _04060_ _04063_ _04070_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09445__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08293_ _03948_ _03967_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12835__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13529__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12046__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout303_A _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10212__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11885__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16040__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1212_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 net303 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09905__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout312 net314 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_2
XANTENNA__15608__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout323 net324 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_2
Xfanout334 net336 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout345 net347 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10515__B2 _04692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout356 net359 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_2
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_2
X_09816_ net970 net626 net543 vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__o21ai_1
Xfanout378 net380 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_2
Xfanout389 net391 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_2
XFILLER_0_119_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09747_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\] net844 _05261_ _05262_
+ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout937_A _02955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14497__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10279__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09678_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\] net818 net903 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\]
+ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__a221o_1
XANTENNA__09684__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08629_ net97 net1677 net956 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__mux2_1
XANTENNA__08892__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11491__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13323__A1_N team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11640_ net1985 net349 net644 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XANTENNA__09436__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ _05738_ _06110_ net658 _05737_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_64_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13310_ net1694 net984 net965 _03004_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__a22o_1
X_10522_ net498 net403 vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and2_1
X_14290_ net1119 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13241_ _06523_ _02961_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__nand2_1
X_10453_ _04802_ _04822_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10265__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10384_ net402 vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__inv_2
XANTENNA_input66_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13172_ _07387_ _07401_ _07402_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11795__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ net272 net2543 net466 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15288__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16533__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12054_ net278 net2657 net470 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11005_ net418 _06516_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__nor2_1
X_16862_ net1406 vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout890 _04533_ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_6
X_15813_ clknet_leaf_31_wb_clk_i _01953_ _00621_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_16793_ net1337 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15744_ clknet_leaf_105_wb_clk_i _01884_ _00552_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_16889__1433 vssd1 vssd1 vccd1 vccd1 _16889__1433/HI net1433 sky130_fd_sc_hd__conb_1
X_12956_ _03294_ _07378_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__nand2_1
XANTENNA__08609__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11907_ net647 _07199_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__nand2_1
X_15675_ clknet_leaf_126_wb_clk_i _01815_ _00483_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12887_ _07404_ _07406_ _07386_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14626_ net1202 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11838_ _07188_ _07193_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__nor2_2
XANTENNA__09427__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14557_ net1084 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11769_ net350 net2103 net600 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\]
+ _03065_ _03069_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__or4_1
XFILLER_0_114_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14488_ net1194 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16227_ clknet_leaf_125_wb_clk_i _02367_ _01035_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13439_ _03043_ _03044_ _03040_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16845__1389 vssd1 vssd1 vccd1 vccd1 _16845__1389/HI net1389 sky130_fd_sc_hd__conb_1
XFILLER_0_109_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16158_ clknet_leaf_113_wb_clk_i _02298_ _00966_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09060__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15109_ net1108 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ _04491_ _04493_ net972 vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__and3_4
X_16089_ clknet_leaf_17_wb_clk_i _02229_ _00897_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire640_A _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07931_ _03575_ _03612_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15900__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ _03549_ _03572_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09601_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\] net807 _05104_ _05117_
+ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__a211o_1
X_16773__1317 vssd1 vssd1 vccd1 vccd1 _16773__1317/HI net1317 sky130_fd_sc_hd__conb_1
X_07793_ _03451_ _03478_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09532_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\] net754 net746 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09666__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09463_ _04973_ _04975_ _04979_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__or3_1
XFILLER_0_91_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08414_ _04119_ _04120_ _04115_ _04116_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09394_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\] net743 net723 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\]
+ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13137__A2_N net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09418__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08345_ _04050_ _04051_ _04057_ _04043_ _04037_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_30_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1162_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08276_ _03962_ _03987_ _03964_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10984__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08929__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15430__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_A _04536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12504__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1107 net1108 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1118 net1120 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_4
XANTENNA__10532__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1129 net1135 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15580__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15116__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ _04422_ team_02_WB.instance_to_wrap.top.pc\[1\] vssd1 vssd1 vccd1 vccd1 _07334_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__11644__A _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13790_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\] _03278_
+ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09657__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08656__C _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09114__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ net377 _06550_ _07001_ _07262_ _07264_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15460_ clknet_leaf_2_wb_clk_i _01600_ _00268_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12672_ net645 _07212_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__nand2_4
XANTENNA__09409__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14411_ net1200 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16086__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11623_ net389 _06039_ _06042_ _07109_ net392 vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__o311a_1
X_15391_ clknet_leaf_18_wb_clk_i _01531_ _00199_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14342_ net1089 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
X_11554_ net837 _07032_ _07039_ _06117_ _07044_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__o221a_1
Xwire521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09290__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire532 net533 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_4
XFILLER_0_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10975__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10505_ _04994_ _06021_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__nand2_1
X_14273_ net1159 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ _06938_ _06978_ net367 vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14690__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16012_ clknet_leaf_15_wb_clk_i _02152_ _00820_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13224_ net2754 _00012_ net938 _05555_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10436_ _05950_ _05952_ _04823_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12922__B _06244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ _07384_ _07385_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__or2_1
XANTENNA__12414__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\] net922 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__a22o_1
X_12106_ net1727 net361 net584 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__mux2_1
X_10298_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\] net760 net744 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__a22o_1
X_13086_ _07461_ _07462_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13141__A2 _07332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12037_ net357 net2461 net474 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09896__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16845_ net1389 vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16776_ net1320 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ net1128 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
XANTENNA__09648__A2 _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15727_ clknet_leaf_34_wb_clk_i _01867_ _00535_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08856__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ team_02_WB.instance_to_wrap.top.pc\[22\] _06180_ vssd1 vssd1 vccd1 vccd1
+ _07459_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15658_ clknet_leaf_129_wb_clk_i _01798_ _00466_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14609_ net1118 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15589_ clknet_leaf_34_wb_clk_i _01729_ _00397_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08130_ _03809_ _03814_ _03817_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15453__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09281__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09820__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08061_ _03709_ _03740_ _03710_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_133_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12324__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__A1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08963_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\] net785 net845 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\]
+ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07914_ _03632_ _03634_ _03621_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__a21o_1
XANTENNA__13944__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08894_ net32 net1031 net989 net1897 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09887__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07845_ _03558_ _03566_ _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout468_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ _03465_ _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09515_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\] net924 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08847__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14775__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09446_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\] net763 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout802_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\] net874 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\]
+ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a221o_1
XANTENNA__10808__A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08328_ _04030_ _04040_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__and2_1
XANTENNA__09272__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09811__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ _03925_ _03960_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11270_ _06664_ _06772_ net397 vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__mux2_1
X_16888__1432 vssd1 vssd1 vccd1 vccd1 _16888__1432/HI net1432 sky130_fd_sc_hd__conb_1
XFILLER_0_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10221_ _05736_ _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__and2b_2
XANTENNA__12234__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10185__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10152_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] net650 _05668_ vssd1
+ vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a21o_1
XANTENNA__11358__B _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10083_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\] net857 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\]
+ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__a221o_1
X_14960_ net1099 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
XANTENNA__09878__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[1\] vssd1 vssd1 vccd1 vccd1
+ net1467 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ net1204 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14891_ net1151 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
XANTENNA__11685__A2 _04692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08667__B team_02_WB.instance_to_wrap.top.a1.instruction\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16630_ clknet_leaf_100_wb_clk_i _02749_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13842_ net1222 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10893__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16561_ clknet_leaf_96_wb_clk_i _02685_ _01368_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_16844__1388 vssd1 vssd1 vccd1 vccd1 _16844__1388/HI net1388 sky130_fd_sc_hd__conb_1
XANTENNA__08838__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13773_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\]
+ _03265_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11437__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10985_ net606 _06491_ _06497_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_84_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15512_ clknet_leaf_54_wb_clk_i _01652_ _00320_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12724_ _05833_ net669 _07075_ _07175_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16492_ clknet_leaf_95_wb_clk_i _02626_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08683__A team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15443_ clknet_leaf_57_wb_clk_i _01583_ _00251_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ net301 net2616 net435 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__mux2_1
XANTENNA__12409__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ net421 _06749_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15374_ clknet_leaf_80_wb_clk_i _01514_ _00187_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12586_ net274 net2116 net438 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09802__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14325_ net1214 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
X_16772__1316 vssd1 vssd1 vccd1 vccd1 _16772__1316/HI net1316 sky130_fd_sc_hd__conb_1
X_11537_ team_02_WB.instance_to_wrap.top.pc\[6\] net976 _04347_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\]
+ _07028_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14256_ net1092 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
X_11468_ net376 _06773_ _06961_ net381 _06962_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08622__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13207_ _04821_ net936 net1020 net1474 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_81_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10419_ net612 _05251_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14187_ net1203 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10453__A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _06847_ _06896_ net366 vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16101__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13138_ _04280_ _02904_ _02905_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a21o_1
XANTENNA__11983__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13069_ _07430_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1109 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09869__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16251__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13169__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] _03349_ vssd1 vssd1 vccd1
+ vccd1 _03353_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16828_ net1372 vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__buf_2
XANTENNA__15819__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07561_ net1 vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__inv_2
XANTENNA__08829__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16759_ net1303 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_18_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09300_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\] net810 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08593__A net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10100__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09231_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\] net760 net731 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12319__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15969__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09162_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\] net905 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a22o_1
XANTENNA__09254__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08113_ _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13107__A1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ _04588_ _04608_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12843__A _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08044_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03722_ vssd1 vssd1 vccd1
+ vccd1 _03766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold910 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold921 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold932 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold943 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12054__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1125_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold998 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09995_ _05489_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout585_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _04318_ _04339_ _04309_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11116__A1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ net19 net1030 net988 net1659 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout752_A _04376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ _03546_ _03550_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__nand2_1
XANTENNA__15499__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07759_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10770_ net498 net385 _06285_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09493__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09429_ _04934_ _04941_ _04944_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__or4_4
XFILLER_0_17_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12229__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10538__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12440_ net344 net2349 net454 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09245__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13849__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ net355 net2262 net563 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14110_ net1191 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
XANTENNA__16124__CLK clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322_ _06821_ _06822_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__nor2_1
X_15090_ net1098 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14041_ net1136 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11253_ _05127_ net665 _06754_ net795 _06755_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10158__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10204_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\] net746 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11184_ _06629_ _06689_ net370 vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10135_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\] net693 _05650_ _05651_
+ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15992_ clknet_leaf_19_wb_clk_i _02132_ _00800_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08678__A _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11107__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14943_ net1182 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
X_10066_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__inv_2
XANTENNA_output135_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14874_ net1184 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10330__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13825_ net1232 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16613_ clknet_leaf_99_wb_clk_i _02732_ _01406_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12607__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16544_ clknet_leaf_93_wb_clk_i _02668_ _01351_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13756_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10968_ net410 _06480_ _06359_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__o21a_1
XANTENNA__09484__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12707_ _04355_ _06163_ _06249_ _07123_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__o22a_1
X_16475_ clknet_leaf_79_wb_clk_i net1545 _01283_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
X_13687_ net1691 _03200_ _03214_ net1240 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_2_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12139__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10899_ _06413_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15426_ clknet_leaf_124_wb_clk_i _01566_ _00234_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12638_ net2404 net346 net554 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09236__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11978__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15357_ clknet_leaf_88_wb_clk_i _01497_ _00170_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_12569_ net352 net2750 net443 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14308_ net1132 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
X_15288_ clknet_leaf_78_wb_clk_i _01432_ _00101_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold206 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 team_02_WB.instance_to_wrap.top.a1.hexop\[1\] vssd1 vssd1 vccd1 vccd1 net1675
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold228 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ net1686 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ net1189 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
Xhold239 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10149__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout708 _04387_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_6
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout719 _04384_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__clkbuf_4
X_08800_ net1510 net1043 net993 team_02_WB.instance_to_wrap.ramaddr\[31\] vssd1 vssd1
+ vccd1 vccd1 _02625_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12602__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\] net770 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15641__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ net932 vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_59_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08662_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10321__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ _03332_ _03335_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__nand2_1
XANTENNA__13031__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08593_ net52 net51 net54 net53 vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__or4_1
XANTENNA__15791__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16887__1431 vssd1 vssd1 vccd1 vccd1 _16887__1431/HI net1431 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_46_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09475__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13271__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12049__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1075_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\] net890 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\]
+ _04716_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__a221o_1
XANTENNA__09227__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13023__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11888__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\] net788 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1242_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09076_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\] net899 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\]
+ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16297__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08027_ _03712_ _03738_ _03749_ _03745_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__o31a_2
XANTENNA__11189__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold740 team_02_WB.instance_to_wrap.ramload\[20\] vssd1 vssd1 vccd1 vccd1 net2198
+ sky130_fd_sc_hd__dlygate4sd3_1
X_16843__1387 vssd1 vssd1 vccd1 vccd1 _16843__1387/HI net1387 sky130_fd_sc_hd__conb_1
Xhold751 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold762 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold773 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold795 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_A _02957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09978_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\] net868 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a22o_1
XANTENNA__12512__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] net1009 _04447_ _04448_ vssd1
+ vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__a22o_1
XANTENNA__10540__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08505__A2 _04185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\] _04333_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__or3b_2
XFILLER_0_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16771__1315 vssd1 vssd1 vccd1 vccd1 _16771__1315/HI net1315 sky130_fd_sc_hd__conb_1
XFILLER_0_73_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11871_ net344 net2231 net490 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11652__A _04482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ _03289_ net1048 _03127_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__nor3_1
X_10822_ _04971_ net386 vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__nor2_1
X_14590_ net1194 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
XANTENNA__13262__A1 _06490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09466__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10076__A1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ _03078_ _03086_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10753_ team_02_WB.instance_to_wrap.top.pc\[28\] team_02_WB.instance_to_wrap.top.pc\[27\]
+ _06269_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16260_ clknet_leaf_1_wb_clk_i _02400_ _01068_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input96_A wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13472_ team_02_WB.START_ADDR_VAL_REG\[12\] net1068 net1002 vssd1 vssd1 vccd1 vccd1
+ net195 sky130_fd_sc_hd__a21o_1
X_10684_ team_02_WB.instance_to_wrap.top.pc\[13\] _06200_ vssd1 vssd1 vccd1 vccd1
+ _06201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[2\]
+ _00024_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__11798__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12423_ net292 net2429 net455 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__mux2_1
X_16191_ clknet_leaf_111_wb_clk_i _02331_ _00999_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10379__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15142_ net1243 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12354_ net288 net2644 net563 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13317__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11099__A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ _06800_ _06803_ _06806_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_56_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15073_ net1238 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12285_ net271 net2375 net570 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14024_ net1177 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11236_ net1793 net273 net642 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12930__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12422__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ net421 _06673_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10118_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\] net819 net909 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\]
+ _05631_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ clknet_leaf_24_wb_clk_i _02115_ _00783_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11098_ net410 _06606_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14926_ net1113 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
X_10049_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\] net720 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10303__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14857_ net1099 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_118_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ net1226 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13253__A1 team_02_WB.instance_to_wrap.ramaddr\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09457__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14788_ net1132 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16527_ clknet_leaf_67_wb_clk_i _02660_ _01334_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.busy_o
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13739_ _03245_ _03246_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09209__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16458_ clknet_leaf_64_wb_clk_i net1562 _01266_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15409_ clknet_leaf_50_wb_clk_i _01549_ _00217_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16389_ clknet_leaf_97_wb_clk_i _02524_ _01197_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11501__S net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13308__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12516__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09901_ _05405_ _05412_ _05415_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nor4_1
XFILLER_0_22_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13428__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09832_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\] net710 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__a22o_1
XANTENNA__12332__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09763_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\] net830 net887 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout283_A _06657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ _04311_ _04276_ _04320_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__mux2_1
XANTENNA__13952__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09694_ _05207_ _05209_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__or2_1
XANTENNA__09696__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09160__A2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08645_ _04271_ _04273_ _04268_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout450_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1192_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09448__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08576_ _04180_ _04239_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15537__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout715_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10816__A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11558__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09128_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\] net890 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09059_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\] net734 net844 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\]
+ _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ net343 net2751 net473 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
Xhold570 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold592 team_02_WB.instance_to_wrap.top.pad.keyCode\[2\] vssd1 vssd1 vccd1 vccd1
+ net2050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13180__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ _04863_ _05950_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__nor2_1
XANTENNA__15119__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12242__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14958__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15760_ clknet_leaf_33_wb_clk_i _01900_ _00568_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12972_ _07490_ _07491_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__and2_1
XANTENNA__09687__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1270 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14711_ net1174 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
Xhold1281 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09151__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11923_ net300 net2576 net483 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__mux2_1
Xhold1292 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
X_15691_ clknet_leaf_114_wb_clk_i _01831_ _00499_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14642_ net1123 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ net294 net2119 net492 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XANTENNA__09439__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10805_ _04842_ net405 vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__nor2_1
X_14573_ net1154 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11785_ net287 net1806 net595 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__mux2_1
XANTENNA__16462__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13524_ _03073_ _03077_ _03061_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16312_ clknet_leaf_53_wb_clk_i _02452_ _01120_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10736_ _06245_ net655 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] net496
+ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12925__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16243_ clknet_leaf_56_wb_clk_i _02383_ _01051_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13455_ _03036_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__nand2_1
X_10667_ _06128_ _06183_ _04490_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__a21oi_4
XANTENNA__12417__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12406_ net351 net2008 net461 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__mux2_1
X_16174_ clknet_leaf_9_wb_clk_i _02314_ _00982_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13386_ net2757 net1011 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[15\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_10_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09611__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10598_ _04462_ _06114_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15125_ net1227 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
XANTENNA__08965__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
X_12337_ net358 net2647 net565 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15056_ net1258 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12268_ net332 net2627 net575 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__mux2_1
X_16886__1430 vssd1 vssd1 vccd1 vccd1 _16886__1430/HI net1430 sky130_fd_sc_hd__conb_1
XANTENNA__08630__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ net1123 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
X_11219_ _05081_ _06113_ _06116_ _05082_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__o22a_1
XANTENNA__12152__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ net322 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\] net579 vssd1
+ vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11991__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15958_ clknet_leaf_52_wb_clk_i _02098_ _00766_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09678__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09142__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire516_A _05439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14909_ net1084 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15889_ clknet_leaf_19_wb_clk_i _02029_ _00697_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08430_ _04135_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16842__1386 vssd1 vssd1 vccd1 vccd1 _16842__1386/HI net1386 sky130_fd_sc_hd__conb_1
X_08361_ _04042_ _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08292_ _03969_ _04002_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09850__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12835__B _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12327__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09602__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16770__1314 vssd1 vssd1 vccd1 vccd1 _16770__1314/HI net1314 sky130_fd_sc_hd__conb_1
XFILLER_0_63_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08956__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12851__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1038_A _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12062__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_2
Xfanout324 _06955_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_2
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16335__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout346 net347 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_2
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout357 net359 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_2
X_09815_ _05325_ _05328_ _05329_ _05331_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__nor4_1
XFILLER_0_96_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09381__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 net372 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_2
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_2
XANTENNA_fanout665_A _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\] net767 net703 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\]
+ _05253_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__a221o_1
X_09677_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\] net887 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08628_ net98 net1517 net957 vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold243_A team_02_WB.instance_to_wrap.ramstore\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08559_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04169_ vssd1 vssd1 vccd1
+ vccd1 _04228_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11570_ _05736_ net661 net656 _07056_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09841__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10521_ _04461_ _05963_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12237__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13240_ _06556_ _06588_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_17_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10452_ net615 _04733_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13171_ net228 _07502_ _02932_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10383_ _04422_ net969 _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12122_ net290 net1810 net467 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input59_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ net281 net1911 net471 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11004_ _06514_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__and2_1
XANTENNA__09372__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16861_ net1405 vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_2
XFILLER_0_79_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14688__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 net881 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__buf_6
Xfanout891 _04533_ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_4
X_15812_ clknet_leaf_3_wb_clk_i _01952_ _00620_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12700__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__A team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16792_ net1336 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09124__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15743_ clknet_leaf_110_wb_clk_i _01883_ _00551_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12955_ _07473_ _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11906_ _06280_ _07193_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15674_ clknet_leaf_119_wb_clk_i _01814_ _00482_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12886_ _07386_ _07405_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__nand2_1
XANTENNA__08883__B2 team_02_WB.instance_to_wrap.ramload\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_114_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11219__B1 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11837_ net346 net2175 net589 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
X_14625_ net1215 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14556_ net1149 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11768_ net362 net2109 net599 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__mux2_1
XANTENNA__09832__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16208__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13507_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ _03064_ _03068_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__or4_1
X_10719_ team_02_WB.instance_to_wrap.top.pc\[26\] _06147_ _06235_ vssd1 vssd1 vccd1
+ vccd1 _06236_ sky130_fd_sc_hd__a21oi_1
X_14487_ net1173 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
XANTENNA__12147__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ net1001 net994 _07123_ team_02_WB.instance_to_wrap.top.pc\[0\] vssd1 vssd1
+ vccd1 vccd1 _07185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16226_ clknet_leaf_122_wb_clk_i _02366_ _01034_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13438_ _03043_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11986__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16157_ clknet_leaf_51_wb_clk_i _02297_ _00965_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ team_02_WB.instance_to_wrap.ramload\[31\] net1016 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[31\] sky130_fd_sc_hd__and2_1
XFILLER_0_84_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15232__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16358__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ net1078 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
X_16088_ clknet_leaf_54_wb_clk_i _02228_ _00896_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07930_ _03612_ _03613_ _03636_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__a21oi_2
X_15039_ net1204 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09899__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire633_A _05035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15382__CLK clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\] net831 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\]
+ _05116_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a221o_1
XANTENNA__12610__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07792_ _03490_ _03491_ _03492_ net364 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08596__A net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09531_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\] net722 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__a22o_1
XANTENNA__09115__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11458__B1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09462_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\] net818 _04976_ _04978_
+ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08413_ _04119_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__nor2_1
X_09393_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\] net767 net759 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12846__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout246_A _06372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08344_ _04040_ _04052_ _04024_ _04035_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__and4b_1
XFILLER_0_47_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09823__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12057__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08275_ net1745 _03315_ net982 _03990_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout413_A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1155_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13291__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11896__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10736__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_A _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15725__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1125 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1119 net1120 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_2
XFILLER_0_100_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09354__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12520__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15875__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09729_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\] net830 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\]
+ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ net379 _06347_ _06407_ _06453_ _07263_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08656__D net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08865__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10121__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12671_ net344 net2484 net434 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__B _04463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14410_ net1168 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
X_11622_ net389 _07071_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15390_ clknet_leaf_112_wb_clk_i _01530_ _00198_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09814__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14341_ net1087 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ net795 _07040_ _07041_ net666 _07043_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire511 _05533_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_64_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire533 net534 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10975__A2 _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10504_ _04970_ _04992_ _05039_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14272_ net1151 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
X_11484_ _06298_ _06300_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__or2_1
X_16011_ clknet_leaf_115_wb_clk_i _02151_ _00819_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13223_ net1472 net1018 net938 _05510_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10435_ _04863_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__or2_1
XANTENNA__10188__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09593__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13154_ net228 _07507_ _02918_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__nand3_1
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10366_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\] net926 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12105_ net2607 net352 net582 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
X_16841__1385 vssd1 vssd1 vccd1 vccd1 _16841__1385/HI net1385 sky130_fd_sc_hd__conb_1
XANTENNA__16650__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13085_ net1026 _02861_ net1024 team_02_WB.instance_to_wrap.top.pc\[21\] vssd1 vssd1
+ vccd1 vccd1 _01502_ sky130_fd_sc_hd__a2bb2o_1
X_10297_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\] net692 net846 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a22o_1
X_12036_ net343 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\] net477 vssd1
+ vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16844_ net1388 vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_2
XANTENNA__12430__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16775_ net1319 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_92_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13987_ net1145 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15726_ clknet_leaf_8_wb_clk_i _01866_ _00534_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10112__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ team_02_WB.instance_to_wrap.top.pc\[22\] _06180_ vssd1 vssd1 vccd1 vccd1
+ _07458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15657_ clknet_leaf_120_wb_clk_i _01797_ _00465_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16030__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ _05788_ _05828_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14608_ net1091 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15588_ clknet_leaf_0_wb_clk_i _01728_ _00396_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09805__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14539_ net1202 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ _03771_ _03776_ _03781_ _03759_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16209_ clknet_leaf_22_wb_clk_i _02349_ _01017_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15748__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10179__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12605__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09584__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\] net729 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a22o_1
X_07913_ _03632_ _03634_ _03621_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a21oi_4
XANTENNA__15898__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08893_ net33 net1029 net987 net1741 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_127_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07844_ _03530_ _03559_ _03532_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__a21boi_1
XANTENNA__12340__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ _03474_ _03496_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout363_A _07107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09514_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\] net908 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__a22o_1
XANTENNA__13960__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08847__B2 net1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09445_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\] net739 _04952_ _04955_
+ _04961_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_91_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15278__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16865__1409 vssd1 vssd1 vccd1 vccd1 _16865__1409/HI net1409 sky130_fd_sc_hd__conb_1
XFILLER_0_93_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09376_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\] net922 net886 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08327_ _04038_ _04031_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08258_ _03910_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_116_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12515__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08189_ _03876_ _03896_ _03867_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13200__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ net422 net501 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09575__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10151_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] _04330_ vssd1 vssd1
+ vccd1 vccd1 _05668_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09327__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\] net912 net892 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a22o_1
X_13910_ net1213 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
XANTENNA__12250__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14890_ net1170 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13841_ net1222 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
XANTENNA__07571__C net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16053__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13772_ _03267_ _03268_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__nor2_1
X_16560_ clknet_leaf_94_wb_clk_i _02684_ _01367_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ net974 _06493_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15511_ clknet_leaf_13_wb_clk_i _01651_ _00319_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12723_ _06283_ _07246_ _06375_ _05961_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__or4b_1
X_16491_ clknet_leaf_67_wb_clk_i net1459 _01299_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08683__B team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15442_ clknet_leaf_6_wb_clk_i _01582_ _00250_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12654_ net292 net2148 net434 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _07092_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ net288 net2258 net438 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__mux2_1
X_15373_ clknet_leaf_80_wb_clk_i _01513_ _00186_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10948__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11536_ net1000 _07027_ net947 vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14324_ net1074 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14255_ net1115 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12425__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11467_ net413 _06549_ net424 vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _04774_ net936 net1021 net1678 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_110_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10418_ _05294_ _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and2_1
XANTENNA__08470__A_N team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14186_ net1167 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
X_11398_ _06305_ _06307_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__or2_1
XANTENNA__07577__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13137_ _06911_ net232 net228 _02903_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__a2bb2o_1
X_10349_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\] net709 net705 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09318__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13068_ _07361_ _07362_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__and2b_1
X_12019_ net282 net2007 net476 vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__mux2_1
XANTENNA__12160__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10333__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_45 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16827_ net1371 vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__buf_2
XANTENNA_wire429_A _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07560_ net1240 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16758_ net1302 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15420__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16546__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15709_ clknet_leaf_51_wb_clk_i _01849_ _00517_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16689_ clknet_leaf_77_wb_clk_i _02806_ _01413_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09230_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\] net727 _04736_ _04739_
+ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09161_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\] net885 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\]
+ _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ _03792_ _03830_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_20_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12794__D1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09092_ _04588_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__nor2_1
X_08043_ _03763_ _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12335__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold900 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold911 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12010__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold933 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09557__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold944 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold955 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10363__B _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold966 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13955__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1020_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold988 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _05491_ _05510_ net969 vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__mux2_2
XFILLER_0_25_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold999 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1118_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09309__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ _04458_ _04460_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout480_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12070__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ net20 net1031 _04431_ team_02_WB.instance_to_wrap.ramload\[26\] vssd1 vssd1
+ vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10324__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ _03549_ _03547_ _03536_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__and3b_1
XFILLER_0_135_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14786__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07758_ _03416_ _03479_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_101_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07689_ _03393_ _03394_ _03377_ _03384_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout912_A _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\] net915 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\]
+ _04932_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16840__1384 vssd1 vssd1 vccd1 vccd1 _16840__1384/HI net1384 sky130_fd_sc_hd__conb_1
XFILLER_0_137_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10538__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\] net766 _04874_ _04875_
+ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12370_ net358 net2243 net561 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11321_ net412 _06107_ net418 vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__o21a_1
XANTENNA__12245__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14040_ net1195 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09548__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ _05123_ net661 _06753_ _06037_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__a22o_1
XANTENNA__08024__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16419__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\] net722 _05718_ _05719_
+ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11355__A2 _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ _06688_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input41_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\] net777 net764 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15991_ clknet_leaf_13_wb_clk_i _02131_ _00799_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11385__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14942_ net1189 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
X_10065_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] net792 net652 _05581_
+ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_76_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16569__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09720__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14873_ net1137 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12068__A0 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16612_ clknet_leaf_94_wb_clk_i _02731_ _01405_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[15\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_67_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ net1234 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16543_ clknet_leaf_66_wb_clk_i _00015_ _01350_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_63_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13755_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\] vssd1 vssd1 vccd1
+ vccd1 _03256_ sky130_fd_sc_hd__or3_1
X_10967_ net408 _06479_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13280__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ net72 team_02_WB.EN_VAL_REG _07230_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__mux2_1
XANTENNA__10094__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11291__A1 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16474_ clknet_leaf_74_wb_clk_i net1648 _01282_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13686_ _03200_ _03204_ net1691 vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10898_ _06032_ _06373_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_14_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15425_ clknet_leaf_117_wb_clk_i _01565_ _00233_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12637_ net1786 net351 net555 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12568_ net356 net1976 net442 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09787__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15356_ clknet_leaf_84_wb_clk_i _01496_ _00169_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ net1133 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
X_11519_ net952 _07010_ _07011_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__or3_1
XANTENNA__12155__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15287_ clknet_leaf_78_wb_clk_i _01431_ _00100_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12499_ net331 net1802 net559 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__mux2_1
XANTENNA__10464__A _04885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold207 team_02_WB.instance_to_wrap.ramload\[27\] vssd1 vssd1 vccd1 vccd1 net1665
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09539__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold229 team_02_WB.instance_to_wrap.top.a1.row2\[2\] vssd1 vssd1 vccd1 vccd1 net1687
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ net1191 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11346__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11994__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14169_ net1136 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
Xfanout709 _04387_ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16864__1408 vssd1 vssd1 vccd1 vccd1 _16864__1408/HI net1408 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_33_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] net931 vssd1 vssd1 vccd1
+ vccd1 _04359_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09172__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09711__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08661_ net1058 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] _04286_ vssd1
+ vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07612_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] _03331_ _03333_ vssd1 vssd1
+ vccd1 vccd1 _03335_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08592_ net50 net39 net64 _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09213_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\] net926 net809 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\]
+ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__a221o_1
XANTENNA__13023__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12854__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_A _06975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09144_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\] net846 _04654_ _04658_
+ _04660_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1068_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09075_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\] net907 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a22o_1
XANTENNA__12065__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1235_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ _03720_ _03728_ _03731_ _03748_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold730 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout695_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold752 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold774 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15466__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout862_A _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\] net835 net807 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\]
+ _05493_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ _04173_ _04218_ _04232_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a22o_1
XANTENNA__09163__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09702__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10848__A1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08859_ net1642 net1039 net1036 team_02_WB.instance_to_wrap.ramstore\[5\] vssd1 vssd1
+ vccd1 vccd1 _02567_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ net349 net1863 net493 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10821_ _05017_ net404 _06336_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11652__B _04488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10752_ team_02_WB.instance_to_wrap.top.pc\[26\] _06268_ vssd1 vssd1 vccd1 vccd1
+ _06269_ sky130_fd_sc_hd__and2_1
X_13540_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\] _03061_ _03097_ _03098_
+ net1067 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__o221a_1
XANTENNA__10076__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ team_02_WB.START_ADDR_VAL_REG\[11\] net1069 net1004 vssd1 vssd1 vccd1 vccd1
+ net194 sky130_fd_sc_hd__a21o_1
XFILLER_0_125_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10683_ net790 _05785_ _06127_ _06199_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__o22a_2
XFILLER_0_137_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15210_ clknet_leaf_66_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[1\]
+ _00023_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] sky130_fd_sc_hd__dfrtp_4
X_12422_ net284 net2448 net455 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09769__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16190_ clknet_leaf_118_wb_clk_i _02330_ _00998_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input89_A wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16241__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15141_ net1243 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
X_12353_ net276 net2142 net562 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11304_ net671 _06792_ _06805_ net838 vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__o2bb2a_1
X_15072_ net1261 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
XANTENNA__15809__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12284_ net260 net2218 net570 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14023_ net1117 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11235_ net606 _06732_ _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__and3_4
XANTENNA__12703__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10000__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ _06401_ _06665_ net415 vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10117_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\] net885 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__a22o_1
XANTENNA__15959__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15974_ clknet_leaf_50_wb_clk_i _02114_ _00782_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11097_ _06479_ _06605_ net399 vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_69_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10048_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\] net680 net676 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a22o_1
X_14925_ net1156 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold90 net179 vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11500__A2 _06989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08901__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14856_ net1177 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ net1231 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13253__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14787_ net1147 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11054__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11999_ net335 net2135 net480 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16526_ clknet_leaf_36_wb_clk_i _00016_ _01333_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10067__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13738_ net2578 _03244_ net949 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11989__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15339__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16457_ clknet_leaf_64_wb_clk_i net1482 _01265_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13669_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15408_ clknet_leaf_39_wb_clk_i _01548_ _00216_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16388_ clknet_leaf_91_wb_clk_i _02523_ _01196_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15339_ clknet_leaf_64_wb_clk_i _01482_ _00152_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15489__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\] net914 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\]
+ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12613__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09393__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09932__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\] net750 _05338_ _05341_
+ _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_123_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09762_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\] net814 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\]
+ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09145__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__inv_2
X_09693_ net523 _05206_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__nand2_1
XANTENNA__08499__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08644_ net1058 _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_29_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08575_ team_02_WB.instance_to_wrap.top.a1.hexop\[4\] _04231_ _04228_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_7_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout443_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10058__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09999__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11899__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout708_A _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10816__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08959__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\] net821 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\]
+ _04643_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_105_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09058_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\] net751 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a22o_1
XANTENNA__10230__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08009_ _03726_ _03727_ _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__nor3_1
XFILLER_0_102_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold560 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12523__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11020_ _05970_ _05971_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__nand2b_2
Xhold582 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold593 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12971_ team_02_WB.instance_to_wrap.top.pc\[4\] _05742_ vssd1 vssd1 vccd1 vccd1 _07491_
+ sky130_fd_sc_hd__or2_1
XANTENNA__13483__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1260 team_02_WB.START_ADDR_VAL_REG\[2\] vssd1 vssd1 vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15135__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1271 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
X_14710_ net1092 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1282 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ net292 net2604 net482 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__mux2_1
XANTENNA__10297__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1293 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ clknet_leaf_0_wb_clk_i _01830_ _00498_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14641_ net1117 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11853_ net287 net1979 net492 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10049__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10804_ _04886_ net387 vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__nor2_1
X_11784_ net275 net2747 net593 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__mux2_1
X_14572_ net1080 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08972__A _04482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16311_ clknet_leaf_116_wb_clk_i _02451_ _01119_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13523_ _03077_ _03081_ _03083_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__o21bai_1
X_10735_ _06161_ _06251_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16863__1407 vssd1 vssd1 vccd1 vccd1 _16863__1407/HI net1407 sky130_fd_sc_hd__conb_1
XFILLER_0_126_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16242_ clknet_leaf_6_wb_clk_i _02382_ _01050_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15631__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10666_ net995 _05441_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__nand2_1
X_13454_ _03032_ _02763_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12405_ net362 net2157 net460 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__mux2_1
X_13385_ net2763 net1011 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[14\]
+ sky130_fd_sc_hd__and2_1
X_16173_ clknet_leaf_24_wb_clk_i _02313_ _00981_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10597_ _04464_ _04467_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__or2_2
XFILLER_0_134_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15124_ net1231 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12336_ net342 net2421 net568 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__mux2_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08911__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12941__B _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15055_ net1261 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XANTENNA__12433__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ net335 net2667 net575 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08178__B2 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__inv_2
X_14006_ net1093 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
XANTENNA__09375__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12198_ net317 net2570 net577 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__mux2_1
X_11149_ net607 _06649_ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__and3_2
XFILLER_0_37_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09127__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15957_ clknet_leaf_50_wb_clk_i _02097_ _00765_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15045__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ net1148 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
XANTENNA__10288__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15888_ clknet_leaf_41_wb_clk_i _02028_ _00696_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire509_A _05578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14839_ net1173 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08360_ _04034_ _04041_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16509_ clknet_leaf_29_wb_clk_i _02643_ _01316_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08291_ _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__inv_2
XANTENNA__12608__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10212__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12851__B _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12343__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09366__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 _06815_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09905__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_1
Xfanout325 _06975_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_2
Xfanout336 _06994_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_1
X_09814_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\] net833 net817 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\]
+ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__a221o_1
Xfanout347 _07187_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_103_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout369 net372 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1100_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\] net695 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout560_A _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15504__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout658_A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10279__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\] net830 net826 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\]
+ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08627_ net99 net1652 net956 vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08892__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14794__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15654__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ _03292_ _04226_ _04180_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12518__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ team_02_WB.instance_to_wrap.top.a1.state\[1\] _04184_ net850 net1769 vssd1
+ vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10520_ _04461_ _05963_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__nor2_4
XFILLER_0_110_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10451_ net615 _04733_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13170_ _07487_ _07488_ _07501_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__nand3b_1
XANTENNA__10203__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ net971 net648 vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12121_ net278 net2047 net468 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12253__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10562__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09357__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ net269 net1871 net470 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__mux2_1
Xhold390 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _06349_ _06512_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__nand2_1
X_16860_ net1404 vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_73_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09109__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net873 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_8
X_15811_ clknet_leaf_12_wb_clk_i _01951_ _00619_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout881 _04538_ vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__buf_4
Xfanout892 _04533_ vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__buf_6
X_16791_ net1335 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__08686__B team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15742_ clknet_leaf_118_wb_clk_i _01882_ _00550_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12664__A0 _07013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ team_02_WB.instance_to_wrap.top.pc\[13\] _06205_ vssd1 vssd1 vccd1 vccd1
+ _07474_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1090 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11905_ net347 net2347 net486 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15673_ clknet_leaf_111_wb_clk_i _01813_ _00481_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12885_ net509 _05582_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12416__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14624_ net1155 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11836_ net350 net2126 net592 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14555_ net1156 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
X_11767_ net355 net1679 net599 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__mux2_1
XANTENNA__12428__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14209__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10718_ _06148_ _06234_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14486_ net1093 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
XANTENNA__10456__B _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11698_ net952 _07183_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16225_ clknet_leaf_121_wb_clk_i _02365_ _01033_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13437_ _03036_ _03038_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__xor2_1
XFILLER_0_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ _04350_ _06165_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09596__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16156_ clknet_leaf_47_wb_clk_i _02296_ _00964_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13368_ team_02_WB.instance_to_wrap.ramload\[30\] net1016 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[30\] sky130_fd_sc_hd__and2_1
XANTENNA__09060__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ net1104 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12319_ net281 net2288 net566 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__mux2_1
XANTENNA__12163__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16087_ clknet_leaf_13_wb_clk_i _02227_ _00895_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13299_ team_02_WB.instance_to_wrap.top.pc\[10\] net1051 _06950_ net933 vssd1 vssd1
+ vccd1 vccd1 _02999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13144__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ net1223 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15527__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _03572_ _03582_ _03540_ net329 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_wire626_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07791_ _03490_ net364 vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08596__B net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09530_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\] net706 _05045_ _05046_
+ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15677__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09520__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09461_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\] net915 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\]
+ _04977_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08412_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04106_ vssd1 vssd1 vccd1
+ vccd1 _04120_ sky130_fd_sc_hd__or2_1
X_09392_ _04908_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12846__B _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08343_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12338__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08274_ _03962_ _03988_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13958__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12862__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09587__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1148_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12850__A_N net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11478__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12073__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout775_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1116 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_4
XANTENNA__16452__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12801__S _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16862__1406 vssd1 vssd1 vccd1 vccd1 _16862__1406/HI net1406 sky130_fd_sc_hd__conb_1
X_07989_ _03706_ _03711_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11417__S net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\] net834 net900 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09511__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09659_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\] net687 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12670_ net350 net2233 net437 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09411__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__C _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11621_ net393 _07035_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12248__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08672__D team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14340_ net1130 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11552_ _05916_ _06110_ _07042_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__a21oi_1
Xwire501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09290__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire523 net524 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_4
XFILLER_0_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire534 _04841_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_2
X_10503_ _05208_ _05979_ _05978_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14271_ net1169 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XANTENNA__10991__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11483_ net411 _06579_ net418 vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ clknet_leaf_128_wb_clk_i _02150_ _00818_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09578__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input71_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ net624 net937 net1018 net1525 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__a2bb2o_1
X_10434_ net535 _04822_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10365_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\] net898 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\]
+ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__a221o_1
X_13153_ _07505_ _07506_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13126__A1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12104_ net2606 net357 net581 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
X_13084_ _06683_ net233 _02860_ net978 _02858_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10296_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\] net752 net736 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\]
+ _05812_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12035_ net339 net1676 net477 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08697__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09750__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16843_ net1387 vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_2
XFILLER_0_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16774_ net1318 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
X_13986_ net1151 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09502__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15725_ clknet_leaf_32_wb_clk_i _01865_ _00533_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12937_ team_02_WB.instance_to_wrap.top.pc\[23\] _06177_ vssd1 vssd1 vccd1 vccd1
+ _07457_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15656_ clknet_leaf_14_wb_clk_i _01796_ _00464_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12868_ _05742_ _05782_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__nand2_2
XFILLER_0_29_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14607_ net1111 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
X_11819_ net286 net2671 net591 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__mux2_1
XANTENNA__12158__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15587_ clknet_leaf_2_wb_clk_i _01727_ _00395_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12799_ _04325_ _04355_ _06161_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__nor3_1
XFILLER_0_12_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14538_ net1143 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
XANTENNA__16325__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11997__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14469_ net1087 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16208_ clknet_leaf_38_wb_clk_i _02348_ _01016_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09569__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ clknet_leaf_16_wb_clk_i _02279_ _00947_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16809__1353 vssd1 vssd1 vccd1 vccd1 _16809__1353/HI net1353 sky130_fd_sc_hd__conb_1
XFILLER_0_126_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13117__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08792__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\] net764 net733 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07912_ _03632_ _03633_ _03621_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12621__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08892_ net3 net1031 net989 net2197 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09741__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ _03561_ _03563_ _03564_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__and3b_1
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07774_ net364 vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13319__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09513_ _05023_ _05025_ _05027_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12857__A _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1098_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09444_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\] net771 _04957_ _04958_
+ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12068__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09375_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\] net821 net906 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\]
+ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08326_ _04015_ _04017_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09272__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08257_ _03925_ _03953_ _03960_ _03927_ _03913_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_116_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08188_ _03888_ _03893_ _03862_ _03868_ _03877_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_127_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout892_A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_103_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ _05660_ _05662_ _05664_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nor4_2
XANTENNA__09980__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10081_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\] net835 net799 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\]
+ _05585_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__a221o_1
XANTENNA__12531__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10840__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15992__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ net1224 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
XANTENNA__10893__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13771_ net1749 _03265_ net961 vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10986__S net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10983_ net999 _06494_ _06495_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15510_ clknet_leaf_47_wb_clk_i _01650_ _00318_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12722_ _06469_ _06500_ _07245_ _06426_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__or4b_1
X_16490_ clknet_leaf_71_wb_clk_i net1511 _01298_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16348__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__C team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15441_ clknet_leaf_22_wb_clk_i _01581_ _00249_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ net287 net2693 net436 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ net375 _06940_ _07090_ _07091_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_33_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09799__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15372_ clknet_leaf_76_wb_clk_i _01512_ _00185_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12584_ net276 net2359 net439 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15372__CLK clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14323_ net1165 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11535_ team_02_WB.instance_to_wrap.top.pc\[6\] _06255_ vssd1 vssd1 vccd1 vccd1 _07027_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14254_ net1113 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
X_11466_ _06869_ _06960_ net394 vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13205_ net636 net937 net1018 net1532 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__a2bb2o_1
X_10417_ _05931_ _05933_ _05335_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__o21a_1
X_14185_ net1109 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
X_11397_ _05931_ _06894_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10030__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ _07377_ _07414_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__xnor2_1
X_10348_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\] net721 net701 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__a22o_1
X_13067_ team_02_WB.instance_to_wrap.top.pc\[24\] _07349_ _02845_ _02846_ vssd1 vssd1
+ vccd1 vccd1 _01505_ sky130_fd_sc_hd__o22a_1
X_10279_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\] net928 net799 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\]
+ _05789_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12018_ net269 net2232 net474 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16826_ net1370 vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__buf_2
XFILLER_0_136_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16757_ net1301 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XANTENNA__08829__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ net1253 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
XANTENNA__13283__B1 _06759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10097__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15708_ clknet_leaf_49_wb_clk_i _01848_ _00516_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16688_ clknet_leaf_77_wb_clk_i _02805_ _01412_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09051__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ clknet_leaf_116_wb_clk_i _01779_ _00447_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10197__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15715__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09160_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\] net913 net889 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09254__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ _03792_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_17_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11597__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09091_ net972 net638 net545 vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__o21a_1
X_16861__1405 vssd1 vssd1 vccd1 vccd1 _16861__1405/HI net1405 sky130_fd_sc_hd__conb_1
XANTENNA__12616__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08462__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08042_ _03721_ _03760_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15865__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold901 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold923 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold934 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold956 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10021__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09962__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold978 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _05505_ _05509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__or2_1
Xhold989 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08944_ _04309_ _04459_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__or2_2
XANTENNA__12351__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1013_A _03014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ net21 net1030 net988 net1665 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A _07208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13971__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07826_ _03509_ _03538_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07757_ _03452_ _03477_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13274__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A _04379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10088__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__C1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07688_ _03393_ _03394_ _03377_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_36_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09493__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09427_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\] net802 _04930_ _04943_
+ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15395__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout905_A _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09358_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\] net770 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09245__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08309_ _03992_ _04000_ _04007_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__nand3_1
X_09289_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\] net923 net939 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a22o_1
XANTENNA__12526__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10835__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10260__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ net376 _06606_ _06820_ net383 vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11251_ _05126_ net659 vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08024__B team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10202_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\] net734 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__a22o_1
XANTENNA__09953__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11182_ _05016_ net386 _06338_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_73_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10133_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\] net768 net752 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12261__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15990_ clknet_leaf_57_wb_clk_i _02130_ _00798_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10570__A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09705__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A gpio_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _05441_ _05580_ net551 vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__mux2_1
X_14941_ net1081 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
XANTENNA__09136__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__B _06883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13881__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14872_ net1186 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16611_ clknet_leaf_80_wb_clk_i _02730_ _01404_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_13823_ net1234 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08694__B _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15738__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10079__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16542_ clknet_leaf_66_wb_clk_i _00014_ _01349_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11276__C1 _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13754_ net2092 _03254_ _03255_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10966_ _06399_ _06478_ net369 vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16808__1352 vssd1 vssd1 vccd1 vccd1 _16808__1352/HI net1352 sky130_fd_sc_hd__conb_1
XANTENNA__09484__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__B _06244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12705_ net1003 net1069 _04249_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__or3b_1
X_16473_ clknet_leaf_78_wb_clk_i net1661 _01281_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
X_13685_ _03200_ _03204_ _03213_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11291__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10897_ net668 _06398_ _06407_ net796 _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15424_ clknet_leaf_107_wb_clk_i _01564_ _00232_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ net2247 net361 net555 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__mux2_1
XANTENNA__15888__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09236__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12944__B _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15355_ clknet_leaf_88_wb_clk_i _01495_ _00168_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_12567_ net342 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\] net445 vssd1
+ vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12436__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11340__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10251__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ net1208 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
X_11518_ team_02_WB.instance_to_wrap.top.pc\[7\] net973 _04347_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15286_ clknet_leaf_81_wb_clk_i _01430_ _00099_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12498_ net334 net2590 net559 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__mux2_1
Xhold208 team_02_WB.instance_to_wrap.ramstore\[1\] vssd1 vssd1 vccd1 vccd1 net1666
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 team_02_WB.START_ADDR_VAL_REG\[3\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ net1081 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
X_11449_ _05469_ net664 _06943_ net795 _06944_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__o221a_1
XANTENNA__09944__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14168_ net1193 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _07418_ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12171__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15268__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14099_ net1169 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ net1059 net1057 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1
+ vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07611_ _03331_ _03333_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__or2_1
X_16809_ net1353 vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__buf_2
XANTENNA__13256__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08591_ net66 net65 net68 net67 vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09475__A2 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09212_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\] net910 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__a22o_1
XANTENNA__10490__B1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09227__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09143_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\] net765 net729 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\]
+ _04659_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12346__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10242__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\] net894 net939 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16043__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08025_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] _03746_ _03747_ vssd1 vssd1
+ vccd1 vccd1 _03748_ sky130_fd_sc_hd__or3_1
XANTENNA__13966__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1130_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold731 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold753 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10390__A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12081__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\] net864 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16193__CLK clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08927_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] net959 vssd1 vssd1 vccd1
+ vccd1 _04447_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout855_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08858_ net167 net1039 net1035 net1596 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08795__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08910__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ _03512_ _03524_ _03531_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__a21o_2
XANTENNA__08910__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08789_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] net997 _04329_ team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10820_ _05061_ net387 vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__or2_1
XANTENNA__11652__C _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09466__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10751_ team_02_WB.instance_to_wrap.top.pc\[25\] team_02_WB.instance_to_wrap.top.pc\[24\]
+ _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_98_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ team_02_WB.START_ADDR_VAL_REG\[10\] net1068 net1002 vssd1 vssd1 vccd1 vccd1
+ net193 sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_27_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10682_ net995 _04419_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ net273 net2041 net454 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12256__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14037__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10233__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ net1245 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12352_ net281 net2242 net562 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11303_ _05941_ _06804_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_56_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15071_ net1250 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ net264 net2267 net570 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14022_ net1072 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
X_11234_ net974 _06733_ _06738_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ _06669_ _06670_ _06671_ net667 vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10116_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\] net889 net869 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__a22o_1
X_15973_ clknet_leaf_34_wb_clk_i _02113_ _00781_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11096_ _06542_ _06604_ net370 vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__mux2_1
XANTENNA__13486__B1 _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15560__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14924_ net1080 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
X_10047_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\] net732 _05562_ _05563_
+ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_69_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16860__1404 vssd1 vssd1 vccd1 vccd1 _16860__1404/HI net1404 sky130_fd_sc_hd__conb_1
XANTENNA__08909__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 team_02_WB.instance_to_wrap.ramstore\[0\] vssd1 vssd1 vccd1 vccd1 net1538
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 team_02_WB.instance_to_wrap.ramaddr\[8\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
X_14855_ net1101 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
X_13806_ net1231 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14786_ net1210 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09457__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ net327 net2372 net480 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
X_16525_ clknet_leaf_35_wb_clk_i _02659_ _01332_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13737_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\]
+ _03242_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__and3_1
X_10949_ _06141_ _06145_ _06237_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16456_ clknet_leaf_104_wb_clk_i net1616 _01264_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
X_13668_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__or4bb_1
XANTENNA__09209__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15407_ clknet_leaf_36_wb_clk_i _01547_ _00215_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16066__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11016__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ net2669 net274 net554 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__mux2_1
XANTENNA__12166__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16387_ clknet_leaf_80_wb_clk_i _02522_ _01195_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13599_ team_02_WB.instance_to_wrap.top.a1.row1\[58\] _03117_ _03125_ team_02_WB.instance_to_wrap.top.a1.row2\[34\]
+ _03151_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__a221o_1
XANTENNA__10224__A0 _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13275__A1_N _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15338_ clknet_leaf_63_wb_clk_i _01481_ _00151_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15269_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[28\]
+ _00082_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09830_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\] net839 _05342_ _05343_
+ _05346_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15903__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09761_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\] net818 net883 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__a22o_1
XANTENNA__13213__A1_N net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ _04289_ _04311_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__or2_1
X_09692_ net523 _05206_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09696__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ _03298_ team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _04272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13229__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout269_A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08574_ net2399 _04238_ _04225_ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
XANTENNA__09448__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13228__A1_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1080_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12865__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout436_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1178_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11007__A2 _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout603_A _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09126_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\] net926 net813 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a22o_1
XANTENNA__09081__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10766__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09057_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\] net782 net747 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a22o_1
X_08008_ _03692_ net255 _03729_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__a31o_1
XANTENNA__09908__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold550 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
X_16807__1351 vssd1 vssd1 vccd1 vccd1 _16807__1351/HI net1351 sky130_fd_sc_hd__conb_1
XFILLER_0_64_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold583 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
X_09959_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\] net780 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a22o_1
X_12970_ team_02_WB.instance_to_wrap.top.pc\[4\] _05742_ vssd1 vssd1 vccd1 vccd1 _07490_
+ sky130_fd_sc_hd__nand2_1
Xhold1250 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09687__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1261 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11921_ net286 net2434 net484 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__mux2_1
Xhold1272 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 team_02_WB.instance_to_wrap.top.a1.row2\[15\] vssd1 vssd1 vccd1 vccd1 net2741
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14640_ net1092 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
X_11852_ net272 net2476 net490 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09439__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ net390 _06315_ _06316_ _06318_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__a22o_1
XANTENNA__16089__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14571_ net1201 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ net290 net2075 net595 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__mux2_1
XANTENNA__08972__B _04488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16310_ clknet_leaf_46_wb_clk_i _02450_ _01118_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13522_ _03078_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nor2_1
X_10734_ _04344_ _04349_ _04354_ net849 vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16241_ clknet_leaf_23_wb_clk_i _02381_ _01049_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13453_ _03038_ _03055_ _02768_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10665_ team_02_WB.instance_to_wrap.top.pc\[21\] _06180_ vssd1 vssd1 vccd1 vccd1
+ _06182_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12404_ net354 net2331 net460 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__mux2_1
XANTENNA__10206__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16172_ clknet_leaf_24_wb_clk_i _02312_ _00980_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13384_ net2758 net1012 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[13\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13089__A2_N net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10596_ _04460_ _04468_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__nand2_4
XANTENNA__09611__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output188_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15123_ net1227 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12335_ net339 net2391 net567 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15054_ net1261 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12266_ net327 net2414 net575 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14005_ net1184 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11217_ net373 _06472_ _06721_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12197_ net312 net2574 net577 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__mux2_1
XANTENNA__11182__A1 _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11148_ net974 _06651_ _06654_ _06655_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__a211o_1
X_11079_ net953 _06588_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__nand2_1
X_15956_ clknet_leaf_10_wb_clk_i _02096_ _00764_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09678__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ net1159 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15887_ clknet_leaf_38_wb_clk_i _02027_ _00695_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14838_ net1095 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14769_ net1118 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16508_ clknet_leaf_37_wb_clk_i _02642_ _01315_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_08290_ _04003_ _04004_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09850__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16439_ clknet_leaf_104_wb_clk_i net1593 _01247_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09602__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12624__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08810__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout304 net305 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_2
Xfanout315 _06914_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_2
Xfanout326 _06975_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout337 net340 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_2
X_09813_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\] net918 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__a22o_1
XANTENNA__13152__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout348 net351 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout359 _07069_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_103_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09744_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\] net735 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\]
+ _05260_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a221o_1
XANTENNA__14140__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09675_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\] net875 net856 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout553_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16231__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08626_ net100 net1605 net954 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout720_A _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04174_ vssd1 vssd1 vccd1
+ vccd1 _04226_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout818_A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08488_ team_02_WB.instance_to_wrap.top.a1.row1\[13\] _04185_ vssd1 vssd1 vccd1 vccd1
+ _02697_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09841__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15949__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09054__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ _04630_ _04652_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09109_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\] net758 net718 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07604__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12534__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08801__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _05882_ _05892_ _05895_ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__nor4_2
XFILLER_0_108_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14315__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12120_ net281 net1932 net466 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ net262 net2618 net471 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold380 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold391 team_02_WB.instance_to_wrap.top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1 net1849
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ net415 _06513_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout860 net861 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_6
XFILLER_0_99_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout871 net873 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_4
X_15810_ clknet_leaf_122_wb_clk_i _01950_ _00618_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout882 _04537_ vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_6
X_16790_ net1334 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
Xfanout893 _04533_ vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14050__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15741_ clknet_leaf_51_wb_clk_i _01881_ _00549_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11467__A2 _06549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12664__A1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ team_02_WB.instance_to_wrap.top.pc\[13\] _06205_ vssd1 vssd1 vccd1 vccd1
+ _07473_ sky130_fd_sc_hd__nand2_1
Xhold1080 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1091 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11904_ net350 net1881 net489 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15672_ clknet_leaf_53_wb_clk_i _01812_ _00480_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12884_ net428 _05627_ _07403_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08983__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14623_ net1190 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11219__A2 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11835_ net363 net2038 net592 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14554_ net1181 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
XANTENNA__09293__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11766_ net358 net2383 net597 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09832__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13505_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10717_ _06151_ _06233_ _06152_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__o21bai_1
X_14485_ net1216 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11697_ _07180_ _07182_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16224_ clknet_leaf_105_wb_clk_i _02364_ _01032_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13436_ _03032_ _03042_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__and2_1
XANTENNA__09045__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648_ _06154_ _06163_ _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08922__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16155_ clknet_leaf_127_wb_clk_i _02295_ _00963_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13367_ team_02_WB.instance_to_wrap.ramload\[29\] net1016 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[29\] sky130_fd_sc_hd__and2_1
XFILLER_0_106_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12444__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14225__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10579_ _04970_ net387 _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15106_ net1078 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
X_12318_ net269 net2390 net565 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__mux2_1
X_16086_ clknet_leaf_48_wb_clk_i _02226_ _00894_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13298_ net2619 net983 net964 _02998_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15037_ net1221 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
X_12249_ net256 net1889 net574 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11155__A1 _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09899__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07790_ _03494_ _03485_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_39_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08859__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15939_ clknet_leaf_13_wb_clk_i _02079_ _00747_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11458__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14895__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09460_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\] net887 net875 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08411_ _04105_ _04111_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__xor2_4
XFILLER_0_87_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09391_ _04886_ _04905_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12619__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16806__1350 vssd1 vssd1 vccd1 vccd1 _16806__1350/HI net1350 sky130_fd_sc_hd__conb_1
X_08342_ _04035_ _04053_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09823__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08273_ _03962_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09036__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12862__B _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12354__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1043_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__B1 _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10382__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1210_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13540__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout670_A _05965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A _04372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07988_ _03707_ _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15621__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09727_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\] net820 net907 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\]
+ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__a221o_1
XANTENNA__11449__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout935_A _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09658_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\] net715 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\]
+ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10121__A2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08609_ net87 net1739 net956 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12529__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\] net912 net884 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a22o_1
XANTENNA__15771__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11620_ net1906 net363 net644 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09275__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09814__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11551_ _05915_ _06116_ net661 _05691_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_53_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10502_ _04950_ _05982_ _05981_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a21o_1
Xwire524 _05186_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_2
X_14270_ net1191 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11482_ _05559_ _06006_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__xor2_1
X_13221_ net625 net937 net1019 net1575 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__a2bb2o_1
X_10433_ _04865_ _05949_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__and2_1
XANTENNA__12264__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14045__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input64_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ net1026 _02917_ net1023 team_02_WB.instance_to_wrap.top.pc\[10\] vssd1 vssd1
+ vccd1 vccd1 _01491_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10364_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\] net825 net821 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12103_ net2370 net343 net584 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
XANTENNA__16277__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13884__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13083_ _07427_ _02859_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12334__A0 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10295_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\] net776 net697 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__a22o_1
XANTENNA__11137__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08002__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12034_ net331 net2056 net475 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__mux2_1
XANTENNA__11688__A2 _07161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08697__B net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__A2 _04215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16842_ net1386 vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_2
XFILLER_0_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout690 _04397_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_8
X_16773_ net1317 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
X_13985_ net1184 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
X_12936_ team_02_WB.instance_to_wrap.top.pc\[24\] _04494_ vssd1 vssd1 vccd1 vccd1
+ _07456_ sky130_fd_sc_hd__or2_1
X_15724_ clknet_leaf_25_wb_clk_i _01864_ _00532_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10112__A2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08917__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12947__B _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15655_ clknet_leaf_29_wb_clk_i _01795_ _00463_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12439__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12867_ net507 _05671_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11818_ net273 net2208 net589 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__mux2_1
X_14606_ net1138 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
X_15586_ clknet_leaf_116_wb_clk_i _01726_ _00394_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08449__A2_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12798_ _07321_ _07258_ _07247_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__or3b_2
XFILLER_0_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09805__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14537_ net1099 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11749_ net278 net1973 net597 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468_ net1127 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16207_ clknet_leaf_38_wb_clk_i _02347_ _01015_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13419_ _03030_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12174__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14399_ net1183 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10179__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11376__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16138_ clknet_leaf_130_wb_clk_i _02278_ _00946_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09049__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13117__A2 _07332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08960_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\] net773 net760 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\]
+ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16069_ clknet_leaf_33_wb_clk_i _02209_ _00877_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15644__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ _03614_ _03615_ _03617_ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__a31o_2
X_08891_ net4 net1029 net987 net1688 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_55_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07842_ _03563_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__nand2_1
XANTENNA__10351__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ _03482_ _03494_ _03495_ _03485_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15794__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\] net811 net896 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\]
+ _05028_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10103__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09443_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\] net715 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\]
+ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a221o_1
XANTENNA__12349__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16719__1447 vssd1 vssd1 vccd1 vccd1 net1447 _16719__1447/LO sky130_fd_sc_hd__conb_1
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09374_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\] net902 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13053__B2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08325_ _04038_ _03321_ net1006 net1785 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13969__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1160_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1258_A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07967__A team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08256_ _03966_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_116_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08480__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12084__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08187_ _03875_ _03904_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_132_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout885_A _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12316__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\] net928 _05584_ _05596_
+ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__a211o_1
XANTENNA__10840__B net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10878__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13770_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\]
+ _03263_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__and3_1
X_10982_ _06143_ net655 net495 team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] net497
+ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__a221o_1
XANTENNA__09496__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13292__B2 _02995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ _06533_ _06566_ _06596_ _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_84_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12259__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15440_ clknet_leaf_38_wb_clk_i _01580_ _00248_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__D team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ net273 net2077 net434 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09248__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11603_ net395 _07016_ net381 vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15371_ clknet_leaf_76_wb_clk_i _01511_ _00184_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13879__A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15517__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ net283 net2020 net439 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14322_ net1122 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
X_11534_ net671 _07014_ _07025_ net673 _07024_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__a221o_2
XFILLER_0_136_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ net1154 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
X_11465_ _06919_ _06959_ net366 vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13204_ _04691_ net936 net1020 net2682 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_111_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15667__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ _05378_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__or2_1
X_14184_ net1178 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09420__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output170_A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11396_ _05381_ _05930_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13135_ _07511_ _02902_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10347_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\] net697 net842 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\]
+ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13066_ _06590_ net234 net230 _02843_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_40_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10278_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\] _04529_ _05791_ _05792_
+ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__a2111o_1
X_12017_ net262 net2535 net476 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__mux2_1
XANTENNA__10333__A2 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11530__A1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16825_ net1369 vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_122_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16756_ net1300 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XANTENNA__09487__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13968_ net1251 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__inv_2
XANTENNA__13283__B2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15707_ clknet_leaf_126_wb_clk_i _01847_ _00515_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12919_ net542 _06139_ _07355_ _07438_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12169__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13899_ net1234 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
X_16687_ clknet_leaf_74_wb_clk_i _02804_ _01411_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10478__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09051__B _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15638_ clknet_leaf_48_wb_clk_i _01778_ _00446_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09239__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10197__B net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16442__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15569_ clknet_leaf_21_wb_clk_i _01709_ _00377_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08110_ _03795_ _03800_ _03815_ _03816_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a22oi_4
XANTENNA__11801__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11597__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09090_ _04593_ _04601_ _04604_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_20_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08041_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _03760_ _03761_ vssd1 vssd1
+ vccd1 vccd1 _03763_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold902 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold913 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold924 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 team_02_WB.instance_to_wrap.ramload\[3\] vssd1 vssd1 vccd1 vccd1 net2393
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold946 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold968 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12632__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ _05494_ _05496_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__or3_1
Xhold979 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08943_ _04309_ _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__nor2_1
XANTENNA__13496__A_N net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout299_A _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08874_ net22 net1030 net988 net1726 vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10324__A2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1006_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ _03536_ _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09190__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout466_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12868__A _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07756_ _03449_ _03451_ _03477_ _03445_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13274__A1 team_02_WB.instance_to_wrap.ramaddr\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07687_ _03403_ _03409_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__nand2_1
XANTENNA__12079__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09426_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\] net834 net919 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\]
+ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09357_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\] net782 net718 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12807__S _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_A _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11711__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ _04020_ _04021_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09288_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\] net887 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08239_ _03942_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ net421 _06749_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09402__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08024__C team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10201_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\] net750 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12542__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11181_ _05041_ _05945_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_73_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07964__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10132_ _05647_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__nor2_2
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10063_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] _04330_ net650 team_02_WB.instance_to_wrap.top.a1.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a22o_2
X_14940_ net1148 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11512__A1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16315__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ net1174 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16610_ clknet_leaf_80_wb_clk_i _02729_ _01403_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13822_ net1234 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09469__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16541_ clknet_leaf_66_wb_clk_i _00013_ _01348_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_13753_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\] _03254_ net949 vssd1
+ vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_15_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10965_ _06076_ _06079_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__or2_1
XANTENNA__16465__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12704_ net345 net2150 net432 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16472_ clknet_leaf_78_wb_clk_i net1623 _01280_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
X_13684_ net1516 _03199_ net1065 vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10896_ net657 _06402_ _06409_ _06410_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12635_ net2454 net353 net555 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__mux2_1
X_15423_ clknet_leaf_86_wb_clk_i _01563_ _00231_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15354_ clknet_leaf_84_wb_clk_i _01494_ _00167_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_130_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ net337 net2417 net444 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09641__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14305_ net1209 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
X_11517_ net998 _07009_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15285_ clknet_leaf_90_wb_clk_i _01429_ _00098_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12497_ net325 net1736 net559 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__mux2_1
Xhold209 _02563_ vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14236_ net1148 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11448_ _05465_ net661 _06116_ _05466_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12960__B _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14167_ net1172 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12452__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ net422 _06037_ _06388_ _06110_ _06014_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_128_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap529_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16718__1446 vssd1 vssd1 vccd1 vccd1 net1446 _16718__1446/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_52_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _07372_ _07373_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__and2b_1
X_14098_ net1121 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ net1027 _02831_ net1025 team_02_WB.instance_to_wrap.top.pc\[27\] vssd1 vssd1
+ vccd1 vccd1 _01508_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_33_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1260 net1264 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09172__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07610_ team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] _03324_ _03328_ vssd1 vssd1
+ vccd1 vccd1 _03333_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16808_ net1352 vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__buf_2
X_08590_ net70 net69 net41 net40 vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__or4_1
XFILLER_0_117_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16739_ net1284 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09997__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09211_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\] net866 _04715_ _04727_
+ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_27_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10490__B2 _05556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12627__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09142_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\] net737 net693 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09632__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09073_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\] net818 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_92_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08024_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] team_02_WB.instance_to_wrap.top.a1.dataIn\[6\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold710 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold721 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold743 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12362__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold754 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold765 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold776 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16338__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold787 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\] net896 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10390__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ net1495 _04446_ net930 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XANTENNA__09699__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09163__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ net168 net1038 net1033 net1602 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout750_A _04376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11706__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08795__B _04422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ _03530_ _03527_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_1166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08788_ net1058 net650 _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07739_ _03422_ _03459_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__xnor2_4
XANTENNA__12748__D _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10750_ team_02_WB.instance_to_wrap.top.pc\[23\] _06266_ vssd1 vssd1 vccd1 vccd1
+ _06267_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09871__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09409_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\] net763 _04923_ _04924_
+ _04925_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_48_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10681_ team_02_WB.instance_to_wrap.top.pc\[14\] _06197_ vssd1 vssd1 vccd1 vccd1
+ _06198_ sky130_fd_sc_hd__nand2_1
XANTENNA__12537__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12420_ net288 net2183 net455 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12351_ net268 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\] net561 vssd1
+ vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_67_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11302_ _05212_ _05940_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__nor2_1
X_15070_ net1264 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
X_12282_ net259 net2315 net572 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ net1128 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11233_ _06186_ net654 _06737_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15149__A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12272__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10581__A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ net378 _06396_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\] _04529_ net873 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__a22o_1
XANTENNA__15705__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13892__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15972_ clknet_leaf_2_wb_clk_i _02112_ _00780_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11095_ _06072_ _06098_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__or2_1
XANTENNA__08986__A team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09154__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ net1150 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
X_10046_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\] net708 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold70 net108 vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 _02562_ vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08901__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 _02602_ vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ net1082 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15855__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13805_ net1257 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11997_ net322 net2684 net480 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
X_14785_ net1209 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16524_ clknet_leaf_29_wb_clk_i _02658_ _01331_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10948_ _06140_ net655 net495 team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] net497
+ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13736_ _03244_ net949 _03243_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__and3b_1
XFILLER_0_15_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16455_ clknet_leaf_46_wb_clk_i _02590_ _01263_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12447__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__or4b_1
X_10879_ _06066_ _06090_ net366 vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15406_ clknet_leaf_9_wb_clk_i _01546_ _00214_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ net1834 net289 net555 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__mux2_1
X_16386_ clknet_leaf_92_wb_clk_i _02521_ _01194_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13598_ team_02_WB.instance_to_wrap.top.a1.row1\[114\] _03121_ _03123_ team_02_WB.instance_to_wrap.top.a1.row2\[42\]
+ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__a22o_1
XANTENNA__09614__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10224__A1 _05740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08968__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15337_ clknet_leaf_104_wb_clk_i _01480_ _00150_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12549_ net270 net1980 net444 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _06626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ clknet_leaf_67_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[27\]
+ _00081_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14219_ net1201 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12182__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15199_ net1260 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09393__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14898__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15385__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09760_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\] net919 net810 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\]
+ _05276_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__a221o_1
XANTENNA__16630__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ net1061 _04309_ _04339_ _04316_ _04268_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__o32a_1
XANTENNA__09145__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ _05187_ _05206_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__and2_1
Xfanout1090 net1097 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_2
X_08642_ net1057 _04270_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10160__B1 _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13229__B2 _05760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08573_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] _04228_ _04230_ _02812_
+ _04227_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12865__B _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout331_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12357__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1073_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09605__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09125_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\] _04529_ _04530_
+ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\] _04641_ vssd1 vssd1 vccd1
+ vccd1 _04642_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08959__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1240_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09056_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\] net763 _04570_ _04572_
+ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08007_ net255 _03691_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout798_A _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15728__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12092__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold540 team_02_WB.instance_to_wrap.top.a1.row1\[15\] vssd1 vssd1 vccd1 vccd1 net1998
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold551 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold562 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold573 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold584 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout965_A _02957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\] net736 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a22o_1
XANTENNA__15878__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08909_ net1514 _04436_ net930 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
XANTENNA__11479__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\] net805 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\]
+ _05401_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1240 team_02_WB.instance_to_wrap.top.a1.row2\[41\] vssd1 vssd1 vccd1 vccd1 net2698
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11920_ net272 net2509 net482 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__mux2_1
Xhold1262 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
X_11851_ net290 net2317 net492 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ net390 _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14570_ net1167 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ net277 net2052 net594 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09844__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10733_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _06161_ _06248_ net953 vssd1
+ vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__a31o_1
X_13521_ team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[1\] team_02_WB.instance_to_wrap.top.pad.keyCode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__or4b_2
XFILLER_0_3_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12267__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14048__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16240_ clknet_leaf_41_wb_clk_i _02380_ _01048_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13452_ _02764_ _02765_ _03036_ _02763_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__or4_1
X_10664_ team_02_WB.instance_to_wrap.top.pc\[21\] _06180_ vssd1 vssd1 vccd1 vccd1
+ _06181_ sky130_fd_sc_hd__and2_1
XANTENNA_input94_A wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12403_ net358 net1867 net458 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13383_ net1683 net1012 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[12\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_24_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16171_ clknet_leaf_117_wb_clk_i _02311_ _00979_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10595_ _04460_ _04468_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15122_ net1227 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12334_ net332 net2533 net567 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15053_ net1261 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
X_12265_ net322 net2689 net575 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16653__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11613__A2_N net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14004_ net1074 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11216_ net424 _06475_ _06638_ _06471_ net376 vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__a221o_1
XANTENNA__09375__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ net306 net2263 net577 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ _06177_ net654 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] net496
+ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09127__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15955_ clknet_leaf_55_wb_clk_i _02095_ _00763_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11078_ _06580_ _06584_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_76_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14906_ net1183 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
X_10029_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\] net815 net799 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\]
+ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__a221o_1
X_15886_ clknet_leaf_9_wb_clk_i _02026_ _00694_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14837_ net1215 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
XANTENNA__16033__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09835__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14768_ net1091 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16507_ clknet_leaf_7_wb_clk_i _02641_ _01314_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13719_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14699_ net1150 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16438_ clknet_leaf_103_wb_clk_i net1576 _01246_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16183__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16369_ clknet_leaf_23_wb_clk_i _02509_ _01177_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09366__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _06891_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_26_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09812_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\] net821 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\]
+ _05316_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__a221o_1
Xfanout327 _06975_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12640__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout338 net340 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
Xfanout349 net351 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09118__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\] net779 net775 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout379_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09674_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\] net911 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\]
+ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__a221o_1
XANTENNA__10133__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11881__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08625_ net101 net2249 net955 vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__mux2_1
XANTENNA__11692__C_N _07177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1190_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12876__A _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout546_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ net1045 _04183_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__nor2_2
XANTENNA__16526__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15400__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_122_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12087__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08487_ _04168_ _04179_ _04183_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__or3_2
XFILLER_0_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout713_A _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13500__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\] net750 net722 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\]
+ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10380_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\] net833 net894 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\]
+ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a221o_1
XANTENNA__08801__B2 team_02_WB.instance_to_wrap.ramaddr\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09039_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\] net888 net877 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\]
+ _04553_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12050_ net266 net2613 net471 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09357__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold370 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 team_02_WB.instance_to_wrap.top.a1.row2\[10\] vssd1 vssd1 vccd1 vccd1 net1850
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net398 _06346_ _06512_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12550__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10372__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 _04186_ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 _04544_ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_4
XANTENNA__09109__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_6
Xfanout883 _04537_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16056__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout894 net897 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11166__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15740_ clknet_leaf_44_wb_clk_i _01880_ _00548_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12952_ team_02_WB.instance_to_wrap.top.pc\[14\] _06200_ vssd1 vssd1 vccd1 vccd1
+ _07472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1070 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1081 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1092 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11903_ net360 net1844 net487 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__mux2_1
X_15671_ clknet_leaf_116_wb_clk_i _01811_ _00479_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12883_ _07387_ _07401_ _07402_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14622_ net1194 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11834_ net353 net2620 net591 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11765_ net342 net2629 net600 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__mux2_1
X_14553_ net1140 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_82_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13504_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__or4_1
X_10716_ team_02_WB.instance_to_wrap.top.pc\[24\] _06172_ _06232_ vssd1 vssd1 vccd1
+ vccd1 _06233_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14484_ net1089 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_11_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11696_ _04458_ _04468_ _07177_ _07181_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16223_ clknet_leaf_86_wb_clk_i _02363_ _01031_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ _04344_ _04349_ _06161_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__and3_1
X_13435_ _03030_ _02765_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13212__A1_N net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13366_ team_02_WB.instance_to_wrap.ramload\[28\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[28\] sky130_fd_sc_hd__and2_1
XFILLER_0_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09596__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16154_ clknet_leaf_120_wb_clk_i _02294_ _00962_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10578_ _05017_ net387 vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15105_ net1098 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12317_ net261 net2046 net566 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__mux2_1
X_16085_ clknet_leaf_43_wb_clk_i _02225_ _00893_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13297_ team_02_WB.instance_to_wrap.top.pc\[11\] net1051 _06931_ net933 vssd1 vssd1
+ vccd1 vccd1 _02998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ net1219 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
X_12248_ net250 net2348 net573 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13144__A3 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12179_ net247 net2601 net578 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__mux2_1
XANTENNA__12460__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap609_A _05781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11560__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13301__B1 _06970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15938_ clknet_leaf_117_wb_clk_i _02078_ _00746_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10115__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09520__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15869_ clknet_leaf_51_wb_clk_i _02009_ _00677_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08410_ _04105_ _04111_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__nand2b_1
X_09390_ _04886_ _04905_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08341_ _04030_ _04040_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15573__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08272_ _03981_ _03986_ _03964_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12635__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09587__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1036_A _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09339__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16079__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12370__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07987_ _03645_ _03695_ _03696_ _03703_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_138_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09726_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\] net893 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11854__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09511__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\] net775 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout830_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout928_A _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08608_ net88 net1551 net957 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
X_09588_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\] net823 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a22o_1
X_08539_ _03313_ _04184_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11015__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11082__A1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11550_ net381 _06382_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire503 net504 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ _05985_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__nor2_1
X_11481_ net2026 net325 net643 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
Xwire525 net527 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_46_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12545__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_4
XFILLER_0_123_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ _05375_ net937 net1018 net1592 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09578__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ _04907_ _05948_ _04908_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13151_ _06952_ net232 _02916_ net977 _02915_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10363_ net368 _05876_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ net1898 net340 net584 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13082_ _04970_ _06180_ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input57_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\] net684 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\]
+ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__a221o_1
XANTENNA__11137__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12033_ net336 net2564 net475 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12280__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15446__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16841_ net1385 vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_2
XANTENNA__09750__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10896__A1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15307__D team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 net681 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_6
XFILLER_0_75_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout691 _04397_ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__buf_4
X_16772_ net1316 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
X_13984_ net1158 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15723_ clknet_leaf_117_wb_clk_i _01863_ _00531_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09502__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12935_ team_02_WB.instance_to_wrap.top.pc\[24\] _04491_ _04493_ vssd1 vssd1 vccd1
+ vccd1 _07455_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15654_ clknet_leaf_49_wb_clk_i _01794_ _00462_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12866_ net509 _05582_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14605_ net1154 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11817_ net289 net2608 net591 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__mux2_1
X_15585_ clknet_leaf_123_wb_clk_i _01725_ _00393_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12797_ _07311_ _07312_ _07320_ _07306_ _07294_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__a311o_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14536_ net1175 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ net280 net2580 net598 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08933__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12963__B _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12455__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14467_ net1145 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11679_ _07163_ _07164_ _06021_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_133_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16206_ clknet_leaf_24_wb_clk_i _02346_ _01014_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09569__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13418_ net1066 _03029_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__nand2_2
XFILLER_0_109_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14398_ net1192 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16221__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16137_ clknet_leaf_104_wb_clk_i _02277_ _00945_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13349_ net1688 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[11\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09049__B _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16068_ clknet_leaf_0_wb_clk_i _02208_ _00876_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07910_ _03571_ _03601_ _03626_ _03605_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__or4b_1
XANTENNA__12190__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15019_ net1203 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
X_08890_ net5 net1030 net988 net1683 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10336__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire631_A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07841_ _03517_ _03521_ _03523_ _03553_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__or4_1
XANTENNA__09741__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07772_ _03448_ _03460_ _03483_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__and3_1
X_09511_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\] net827 net920 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09442_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\] net779 net844 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09373_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\] net833 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\]
+ _04889_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout244_A _06372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08324_ _04031_ _04036_ _04014_ _04017_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_30_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08255_ _03947_ _03967_ _03968_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__or3_1
XFILLER_0_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12365__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1153_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08186_ _03888_ _03893_ _03862_ _03871_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15469__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09980__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout878_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11709__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10327__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09709_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\] net787 _05224_ _05225_
+ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__a211o_1
X_10981_ team_02_WB.instance_to_wrap.top.pc\[27\] _06269_ vssd1 vssd1 vccd1 vccd1
+ _06494_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13292__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ _07243_ _06687_ _06658_ _06627_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_84_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ net288 net2727 net436 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08066__A1_N _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ net388 _07089_ _07088_ net392 vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_61_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15370_ clknet_leaf_75_wb_clk_i _01510_ _00183_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[29\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__09799__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ net269 net2622 net439 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08980__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14321_ net1105 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11533_ _05649_ _05917_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12275__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16244__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11464_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__nand2_1
X_14252_ net1071 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08759__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13203_ net1684 net1018 net938 _04650_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__a22o_1
X_10415_ net519 _05334_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14183_ net1120 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
X_11395_ _06013_ _06892_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10346_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\] net689 net846 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10030__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13134_ _07476_ _07478_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__nand2_1
XANTENNA__09971__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13065_ net979 _07432_ _02844_ net1028 vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__o31ai_1
X_10277_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\] net823 net900 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\]
+ _05793_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12016_ net265 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\] net476 vssd1
+ vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
XANTENNA__09184__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11530__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16824_ net1368 vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_122_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16755_ net1299 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13967_ net1254 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
XANTENNA__13283__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10097__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15706_ clknet_leaf_118_wb_clk_i _01846_ _00514_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11294__A1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ _07356_ _07436_ _07357_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__o21a_1
X_16686_ clknet_leaf_77_wb_clk_i _02803_ _01410_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13898_ net1234 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10478__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15637_ clknet_leaf_41_wb_clk_i _01777_ _00445_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12849_ _06190_ net526 vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_48_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ clknet_leaf_41_wb_clk_i _01708_ _00376_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11597__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14519_ net1173 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12185__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15499_ clknet_leaf_116_wb_clk_i _01639_ _00307_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08040_ _03760_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15611__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold903 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold925 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold936 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold947 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10021__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09962__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold958 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\] net884 _05492_ _05507_
+ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a211o_1
X_08942_ _04270_ _04288_ _04318_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__and3_1
XANTENNA__09175__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08873_ net23 net1030 net988 net2463 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_4_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07824_ _03510_ _03534_ _03502_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16117__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09523__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07755_ _03449_ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13274__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout459_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_07686_ _03406_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__nor2_1
XANTENNA__11285__B2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\] net825 net907 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09356_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\] net750 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\]
+ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_118_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08307_ _03997_ _04018_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__xnor2_4
X_09287_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\] _04529_ net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12095__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08238_ _03914_ _03927_ _03905_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10260__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08169_ _03865_ _03867_ _03876_ _03882_ _03887_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__o311a_2
XFILLER_0_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10200_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\] net758 net730 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a22o_1
XANTENNA__10012__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11180_ net1577 net278 net641 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09953__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10131_ net427 _05646_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09166__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09705__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ net508 vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13654__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870_ net1096 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ net1233 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09433__A _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10079__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16540_ clknet_leaf_93_wb_clk_i _02667_ _01347_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[63\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_67_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13752_ _03254_ net949 _03253_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__and3b_1
XFILLER_0_39_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10964_ net376 _06475_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__a21oi_2
X_12703_ net349 net2753 net433 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__mux2_1
X_16471_ clknet_leaf_78_wb_clk_i net1681 _01279_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ _03206_ _03212_ net1241 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10895_ _06122_ _06357_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11902__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15170__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15422_ clknet_leaf_108_wb_clk_i _01562_ _00230_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_14_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ net2556 net357 net554 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11579__A2 _07064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15353_ clknet_leaf_84_wb_clk_i _01493_ _00166_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12565_ net330 net2228 net443 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14304_ net1155 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10251__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11516_ _06256_ _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__or2_1
X_15284_ clknet_leaf_78_wb_clk_i _01428_ _00097_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ net321 net1799 net559 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14235_ net1180 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
X_11447_ net418 _06514_ _06941_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09608__A _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10003__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11378_ _05932_ net661 net658 _05335_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__a22o_1
X_14166_ net1136 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\] net897 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__a22o_1
X_13117_ net791 _07332_ _07515_ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_52_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ net1117 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _06494_ net234 _02828_ net979 _02830_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_33_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1250 net1265 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__clkbuf_4
Xfanout1261 net1263 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16807_ net1351 vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__buf_2
XANTENNA_wire427_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14999_ net1228 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
XANTENNA__13256__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16738_ net1283 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_117_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16669_ clknet_leaf_73_wb_clk_i _02786_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11812__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15080__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09210_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\] net825 net805 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\]
+ _04726_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\] net741 net725 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\]
+ _04657_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11414__A1_N net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10242__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09072_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08023_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] team_02_WB.instance_to_wrap.top.a1.dataIn\[2\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] team_02_WB.instance_to_wrap.top.a1.dataIn\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12643__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold700 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14424__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold711 team_02_WB.instance_to_wrap.ramaddr\[9\] vssd1 vssd1 vccd1 vccd1 net2169
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold722 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold733 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold744 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold755 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold766 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold799 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] net792 _04331_ _05490_
+ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__a22o_2
XFILLER_0_99_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09148__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1116_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08925_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] net1008 _04444_ _04445_ vssd1
+ vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12879__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08856_ net169 net1040 net1036 net1701 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07807_ _03484_ _03528_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08787_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] _04275_ _04329_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout743_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07738_ _03443_ _03447_ _03452_ _03457_ _03460_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a311o_4
XFILLER_0_135_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09320__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout910_A _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07669_ _03345_ net948 _03361_ _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11722__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\] net703 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ net790 _05740_ _06127_ _06196_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__o22a_2
XANTENNA__10481__A2 _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09339_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\] net798 _04843_ _04855_
+ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11023__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12350_ net260 net2739 net561 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10233__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11301_ _06584_ _06798_ _06802_ _06037_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12281_ net249 net2523 net569 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__mux2_1
XANTENNA__12553__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11232_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] net494 _06736_ _04263_ net496
+ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__a221o_1
X_14020_ net1128 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13183__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13183__B2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11163_ net373 _06386_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09139__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10114_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\] net925 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15971_ clknet_leaf_125_wb_clk_i _02111_ _00779_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11094_ _05983_ _06602_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13486__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16432__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\] net772 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__a22o_1
X_14922_ net1143 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold60 team_02_WB.instance_to_wrap.ramaddr\[7\] vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 _02605_ vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 net159 vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ net1136 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
Xhold93 team_02_WB.START_ADDR_VAL_REG\[24\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13804_ net1483 _03288_ net960 vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14784_ net1148 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11996_ net318 net2505 net478 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
XANTENNA__09311__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16729__1453 vssd1 vssd1 vccd1 vccd1 net1453 _16729__1453/LO sky130_fd_sc_hd__conb_1
XANTENNA__16582__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16523_ clknet_leaf_37_wb_clk_i _02657_ _01330_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08325__A2_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13735_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ _03240_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__and3_1
X_10947_ net999 _06460_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16454_ clknet_leaf_104_wb_clk_i net1533 _01262_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfrtp_1
X_13666_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[5\] _03199_ vssd1 vssd1 vccd1
+ vccd1 _03200_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10878_ net398 _06390_ net383 vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15405_ clknet_leaf_33_wb_clk_i _01545_ _00213_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12617_ net1759 net279 net556 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16385_ clknet_leaf_91_wb_clk_i _02520_ _01193_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13597_ team_02_WB.instance_to_wrap.top.a1.row2\[18\] _03124_ _03126_ team_02_WB.instance_to_wrap.top.a1.row2\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15336_ clknet_leaf_64_wb_clk_i _01479_ _00149_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12548_ net262 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\] net444 vssd1
+ vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__mux2_1
XANTENNA__12971__B _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15267_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[26\]
+ _00080_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12463__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 _06626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net250 net2323 net557 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09378__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14218_ net1168 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15198_ net1260 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14149_ net1086 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11807__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ _04278_ _04289_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__nand2_1
XANTENNA__15075__A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ net523 _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1080 net1088 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09550__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08641_ team_02_WB.instance_to_wrap.top.a1.instruction\[14\] net1058 vssd1 vssd1
+ vccd1 vccd1 _04270_ sky130_fd_sc_hd__nand2b_1
Xfanout1091 net1097 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_4
XFILLER_0_77_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08572_ net1728 _04236_ _04225_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09302__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10947__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12638__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14419__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10666__B _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09605__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout324_A _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1066_A _00018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10215__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09947__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a22o_1
XANTENNA__16305__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09081__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09055_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\] net683 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12373__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ _03648_ _03690_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold530 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09908__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout693_A _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold541 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold574 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold585 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09957_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\] net776 _05472_ _05473_
+ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout860_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08908_ net1045 _04193_ _04205_ net1008 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__a32o_1
XANTENNA__11479__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09888_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\] net829 net825 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\]
+ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a221o_1
Xhold1230 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1241 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ net156 net1039 net1035 net1474 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1263 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1285 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1296 team_02_WB.instance_to_wrap.ramstore\[8\] vssd1 vssd1 vccd1 vccd1 net2754
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11850_ net277 net2328 net491 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__mux2_1
XANTENNA__13625__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _04589_ net405 vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12548__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ net280 net2499 net594 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[5\] team_02_WB.instance_to_wrap.top.pad.keyCode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__or4b_2
XFILLER_0_83_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10732_ _04349_ _04354_ _04344_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_67_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11651__B2 _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13451_ _02765_ _03049_ _03054_ _03041_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10663_ _06128_ _06179_ _04490_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_3_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12402_ net342 net2510 net460 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__mux2_1
XANTENNA__10206__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16170_ clknet_leaf_128_wb_clk_i _02310_ _00978_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13382_ net1688 net1010 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[11\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10594_ _04462_ _06109_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__or2_2
XANTENNA_input87_A wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15121_ net1231 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12333_ net335 net1838 net567 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__mux2_1
XANTENNA__12283__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10592__A _04463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15052_ net1219 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12264_ net318 net2488 net573 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14003_ net1169 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11215_ net417 _06719_ _06355_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__o21a_1
X_12195_ net298 net2221 net578 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09780__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11146_ net999 _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11077_ net673 _06566_ _06585_ net672 _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__a221o_1
X_15954_ clknet_leaf_3_wb_clk_i _02094_ _00762_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09532__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14905_ net1129 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
X_10028_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\] net827 net920 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__a22o_1
X_15885_ clknet_leaf_32_wb_clk_i _02025_ _00693_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15972__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14836_ net1076 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12458__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14767_ net1110 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
X_11979_ net253 net2654 net480 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16506_ clknet_leaf_28_wb_clk_i _02640_ _01313_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13718_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\] net949 vssd1 vssd1 vccd1
+ vccd1 _02769_ sky130_fd_sc_hd__and2b_1
XANTENNA__16328__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14698_ net1142 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16437_ clknet_leaf_120_wb_clk_i net1526 _01245_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13649_ _00018_ net1009 _07339_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09599__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16368_ clknet_leaf_33_wb_clk_i _02508_ _01176_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09063__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15319_ clknet_leaf_103_wb_clk_i _01462_ _00132_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15352__CLK clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12193__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16299_ clknet_leaf_116_wb_clk_i _02439_ _01107_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08810__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout306 _06891_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09771__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout317 net320 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_2
X_09811_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\] net858 _05315_ _05327_
+ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout328 _06975_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_1
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_2
X_16785__1329 vssd1 vssd1 vccd1 vccd1 _16785__1329/HI net1329 sky130_fd_sc_hd__conb_1
X_09742_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\] net683 _05256_ _05257_
+ _05258_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09673_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\] net927 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__a22o_1
X_08624_ net102 net1535 net957 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12876__B net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08555_ _04220_ _04221_ net653 net794 net1621 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a32o_1
XANTENNA__12368__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08486_ _04168_ _04184_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__and2b_2
XANTENNA__10396__B _05690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_A _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09054__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09107_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\] net746 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08801__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13138__A1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09038_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\] net812 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\]
+ _04547_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__a221o_1
XANTENNA__15845__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16728__1452 vssd1 vssd1 vccd1 vccd1 net1452 _16728__1452/LO sky130_fd_sc_hd__conb_1
Xhold360 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold371 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold382 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 team_02_WB.instance_to_wrap.ramstore\[5\] vssd1 vssd1 vccd1 vccd1 net1851
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net398 _06511_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__nand2_1
XANTENNA__09762__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout840 net842 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15995__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout851 net852 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_4
Xfanout862 _04543_ vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_8
Xfanout873 _04540_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__buf_4
Xfanout884 _04537_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09514__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 net897 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__buf_4
XANTENNA__13310__B2 _03004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12951_ team_02_WB.instance_to_wrap.top.pc\[14\] _06200_ vssd1 vssd1 vccd1 vccd1
+ _07471_ sky130_fd_sc_hd__nor2_1
Xhold1060 team_02_WB.instance_to_wrap.top.pad.keyCode\[1\] vssd1 vssd1 vccd1 vccd1
+ net2518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13662__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11902_ net353 net2661 net487 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__mux2_1
X_15670_ clknet_leaf_48_wb_clk_i _01810_ _00478_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1082 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12882_ net429 _05627_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__xnor2_1
X_14621_ net1085 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
X_11833_ net356 net2598 net589 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12278__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10587__A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14552_ net1186 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11764_ net339 net2260 net600 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09293__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__nand2_1
X_10715_ _06231_ _06173_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__and2b_1
XANTENNA__15375__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16717__1276 vssd1 vssd1 vccd1 vccd1 _16717__1276/HI net1276 sky130_fd_sc_hd__conb_1
X_14483_ net1168 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11695_ _04569_ _07138_ _07174_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11910__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16222_ clknet_leaf_112_wb_clk_i _02362_ _01030_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13434_ _03036_ _02767_ _02768_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__and3_1
X_10646_ net849 _06161_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09045__A2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ clknet_leaf_16_wb_clk_i _02293_ _00961_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13365_ net1665 net1017 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[27\]
+ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_51_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10577_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__inv_2
XANTENNA__08504__B net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15104_ net1104 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XANTENNA__10060__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12316_ net264 net2592 net566 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16084_ clknet_leaf_12_wb_clk_i _02224_ _00892_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13296_ net1680 net984 net964 _02997_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15035_ net1219 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12247_ net251 net2060 net575 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ net243 net1796 net579 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__mux2_1
X_11129_ net417 _06636_ _06355_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09505__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13301__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15937_ clknet_leaf_117_wb_clk_i _02077_ _00745_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15868_ clknet_leaf_45_wb_clk_i _02008_ _00676_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire507_A _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14819_ net1131 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
XANTENNA__13065__B1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12188__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15718__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15799_ clknet_leaf_116_wb_clk_i _01939_ _00607_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11615__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08340_ _04040_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ _03981_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11820__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15868__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09036__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11379__B1 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08244__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10051__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12651__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09744__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13540__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout391_A _05856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11551__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_A _07198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07986_ _03696_ _03708_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09725_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\] _04529_ _04530_
+ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\] _05241_ vssd1 vssd1 vccd1
+ vccd1 _05242_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout656_A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09656_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\] net683 _05171_ _05172_
+ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09261__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ net89 net1556 net954 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
XANTENNA__15398__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12098__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout823_A _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09587_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\] net896 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__a22o_1
XANTENNA__16643__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08538_ _04222_ net1654 _04186_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XANTENNA__09275__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08469_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11730__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire504 _05735_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_2
X_10500_ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__dlymetal6s2s_1
X_11480_ _06837_ _06974_ _06971_ net605 vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__o211a_2
XFILLER_0_123_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire537 _04801_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_2
X_10431_ _04951_ _05947_ _04948_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_1615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09983__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ _07383_ _07411_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10362_ _05878_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12101_ net2284 net330 net582 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__mux2_1
XANTENNA__16023__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12561__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10293_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\] net772 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__a22o_1
X_13081_ net229 _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12032_ net325 net1790 net475 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__mux2_1
Xhold190 _02609_ vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16840_ net1384 vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_2
XFILLER_0_79_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout670 _05965_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout681 _04407_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_4
X_16771_ net1315 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
Xfanout692 _04397_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_6
XFILLER_0_137_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13983_ net1175 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
XANTENNA__13295__B1 _06908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15722_ clknet_leaf_0_wb_clk_i _01862_ _00530_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11905__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ team_02_WB.instance_to_wrap.top.pc\[25\] _06171_ vssd1 vssd1 vccd1 vccd1
+ _07454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15653_ clknet_leaf_31_wb_clk_i _01793_ _00461_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12865_ _05489_ _05491_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__and2_1
X_14604_ net1080 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11816_ net279 net1797 net590 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15584_ clknet_leaf_108_wb_clk_i _01724_ _00392_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12796_ _07313_ _07315_ _07319_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14535_ net1107 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11747_ net268 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\] net597 vssd1
+ vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11640__S net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16784__1328 vssd1 vssd1 vccd1 vccd1 _16784__1328/HI net1328 sky130_fd_sc_hd__conb_1
XFILLER_0_84_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13421__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10281__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14466_ net1206 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _05016_ _05037_ _05972_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_133_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16205_ clknet_leaf_23_wb_clk_i _02345_ _01013_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13417_ team_02_WB.instance_to_wrap.top.lcd.currentState\[1\] net1050 net962 vssd1
+ vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__mux2_1
X_10629_ team_02_WB.instance_to_wrap.top.a1.instruction\[26\] net996 vssd1 vssd1 vccd1
+ vccd1 _06146_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14397_ net1083 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10033__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16136_ clknet_leaf_14_wb_clk_i _02276_ _00944_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13348_ net2197 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[10\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_80_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16067_ clknet_leaf_127_wb_clk_i _02207_ _00875_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12471__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13279_ team_02_WB.instance_to_wrap.top.pc\[20\] net1052 _06705_ net934 vssd1 vssd1
+ vccd1 vccd1 _02989_ sky130_fd_sc_hd__a22o_1
X_15018_ net1235 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
XANTENNA__09726__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09346__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07840_ _03521_ _03523_ _03553_ _03517_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__o31ai_1
X_07771_ _03474_ _03489_ _03493_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__a21bo_1
XANTENNA__13286__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11815__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\] net831 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\]
+ _05026_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09441_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\] net783 net747 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16727__1451 vssd1 vssd1 vccd1 vccd1 net1451 _16727__1451/LO sky130_fd_sc_hd__conb_1
XFILLER_0_34_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10020__A _05536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\] net914 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08323_ _04031_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__nand2_1
XANTENNA__12646__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10272__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08254_ _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__inv_2
XANTENNA__10674__B _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13210__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08185_ _03901_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1146_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10024__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10575__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12381__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09717__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout773_A _04371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16716__1275 vssd1 vssd1 vccd1 vccd1 _16716__1275/HI net1275 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07969_ _03690_ _03691_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout940_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13277__B1 _06679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13211__A1_N _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11725__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09708_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\] net753 net737 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__a22o_1
X_10980_ _06236_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09496__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09639_ _05149_ _05151_ _05153_ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_84_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11551__A2_N _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ net277 net2465 net435 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__mux2_1
XANTENNA_input104_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13226__A1_N net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09248__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11601_ net498 net385 _06289_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12581_ net262 net2451 net439 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__mux2_1
XANTENNA__12556__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__S net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13241__A _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14320_ net1076 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11532_ net657 _07019_ _07023_ net795 _07022_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ net1150 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11463_ _05514_ net658 _06113_ _05512_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_22_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13202_ net639 _02955_ net1021 net1481 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09956__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ _05381_ _05930_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14182_ net1073 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
X_11394_ _05380_ _06012_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__nor2_1
XANTENNA__11763__A0 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09420__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15168__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13133_ net1026 _02901_ net1023 team_02_WB.instance_to_wrap.top.pc\[13\] vssd1 vssd1
+ vccd1 vccd1 _01494_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10345_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\] net737 net693 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__a22o_1
XANTENNA__12291__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09708__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13064_ _07360_ _07431_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10276_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\] net908 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15563__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ net256 net1822 net476 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08931__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16823_ net1367 vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13966_ net1254 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__inv_2
X_16754_ net1298 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09487__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12917_ _07356_ _07436_ _07357_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__o21ai_1
X_15705_ clknet_leaf_112_wb_clk_i _01845_ _00513_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_16685_ clknet_leaf_73_wb_clk_i _02802_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_13897_ net1251 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12848_ net529 _06188_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__xor2_1
X_15636_ clknet_leaf_11_wb_clk_i _01776_ _00444_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09239__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16069__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15567_ clknet_leaf_36_wb_clk_i _01707_ _00375_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12466__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ _07019_ _07095_ _07112_ _07136_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10254__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ net1092 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15498_ clknet_leaf_128_wb_clk_i _01638_ _00306_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14449_ net1106 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09947__A0 _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10006__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold904 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold915 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold926 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold937 team_02_WB.instance_to_wrap.ramaddr\[13\] vssd1 vssd1 vccd1 vccd1 net2395
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16119_ clknet_leaf_13_wb_clk_i _02259_ _00927_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15078__A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold948 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold959 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09990_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\] net831 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\]
+ _05506_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08941_ _04336_ _04457_ _04309_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_23_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09175__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ net25 net1031 net989 team_02_WB.instance_to_wrap.ramload\[30\] vssd1 vssd1
+ vccd1 vccd1 _02558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07823_ _03544_ _03545_ _03540_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07754_ _03461_ _03462_ _03443_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11285__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07685_ _03363_ _03395_ _03404_ _03407_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout354_A _07087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1096_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _04935_ _04937_ _04938_ _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08438__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\] net742 net698 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a22o_1
XANTENNA__12376__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13431__B1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1263_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08306_ _04019_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_111_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12785__A2 _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09286_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\] net874 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08237_ _03823_ _03926_ _03951_ _03911_ _03924_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_133_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09938__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16855__1399 vssd1 vssd1 vccd1 vccd1 _16855__1399/HI net1399 sky130_fd_sc_hd__conb_1
XFILLER_0_127_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08168_ _03880_ _03883_ _03885_ _03879_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout890_A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_108_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15586__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08099_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] _03762_ _03796_ vssd1 vssd1
+ vccd1 vccd1 _03819_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_73_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10130_ net427 _05646_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10061_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\] net752 _05572_ _05576_
+ _05577_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a2111oi_2
XANTENNA__12170__A0 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16783__1327 vssd1 vssd1 vccd1 vccd1 _16783__1327/HI net1327 sky130_fd_sc_hd__conb_1
XFILLER_0_76_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13820_ net1229 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09469__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13751_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10963_ net378 _06474_ _06473_ net416 vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_67_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12702_ net360 net2274 net432 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16470_ clknet_leaf_79_wb_clk_i net1529 _01278_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
X_13682_ _03199_ _03211_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10894_ _06110_ _06373_ _06408_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__a21oi_1
X_15421_ clknet_leaf_48_wb_clk_i _01561_ _00229_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12633_ net2205 _07051_ net556 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12286__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10236__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15352_ clknet_leaf_84_wb_clk_i _01492_ _00165_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_12564_ net335 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\] net443 vssd1
+ vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09641__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11984__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14303_ net1183 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11515_ team_02_WB.instance_to_wrap.top.pc\[6\] _06255_ team_02_WB.instance_to_wrap.top.pc\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15283_ clknet_leaf_77_wb_clk_i _01427_ _00096_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12495_ net319 net2469 net557 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__mux2_1
XANTENNA__15929__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14234_ net1167 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
XANTENNA__09929__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11446_ net418 _06356_ _06516_ _06941_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13103__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14165_ net1214 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11377_ _06872_ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13116_ _07470_ _07514_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__and2_1
X_10328_ _05838_ _05840_ _05842_ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14096_ net1095 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
X_16726__1450 vssd1 vssd1 vccd1 vccd1 net1450 _16726__1450/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_52_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ net791 _07332_ _07534_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10259_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\] net780 _05772_ _05773_
+ _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_33_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12969__B _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1240 net1242 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08904__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08904__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1251 net1254 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_4
Xfanout1262 net1263 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_2
XANTENNA__15309__CLK clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16806_ net1350 vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__buf_2
X_14998_ net1222 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
X_16737_ team_02_WB.instance_to_wrap.top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1 net177
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13949_ net1210 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15459__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16668_ clknet_leaf_74_wb_clk_i net1460 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.debounce_dly
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09880__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15619_ clknet_leaf_125_wb_clk_i _01759_ _00427_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12196__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16599_ clknet_leaf_96_wb_clk_i _02718_ _01392_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10227__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09140_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\] net721 net689 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16715__1274 vssd1 vssd1 vccd1 vccd1 _16715__1274/HI net1274 sky130_fd_sc_hd__conb_1
XFILLER_0_31_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09632__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09071_ _04581_ _04587_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__nor2_8
XFILLER_0_60_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08022_ _03698_ _03702_ _03705_ _03701_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold701 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold723 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 team_02_WB.instance_to_wrap.top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1 net2214
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold778 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _05442_ _04421_ net551 vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold789 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ net1045 _04215_ _04232_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1011_A _03014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ net170 net1037 net1033 net1472 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout471_A _07208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout569_A _07217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ _03528_ _03484_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08786_ _04406_ _04409_ _04411_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__nor4_2
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07737_ _03424_ _03458_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_81_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout736_A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07668_ _03380_ _03382_ _03354_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_62_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09871__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09407_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\] net679 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__a22o_1
X_07599_ team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] team_02_WB.instance_to_wrap.top.a1.dataIn\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout903_A _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09338_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\] net927 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\]
+ _04854_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__a221o_1
XANTENNA__11415__C1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11966__A0 _07013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09623__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09269_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\] net770 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08831__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14615__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11300_ net373 _06568_ _06801_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_75_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12280_ net251 net2340 net572 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11231_ _06735_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11162_ _06382_ _06638_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10941__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10113_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\] net893 net881 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ clknet_leaf_122_wb_clk_i _02110_ _00778_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11093_ _04951_ _06601_ _04950_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__a21oi_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14921_ net1110 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
X_10044_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\] net748 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_76_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold50 team_02_WB.instance_to_wrap.top.a1.data\[6\] vssd1 vssd1 vccd1 vccd1 net1508
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 _02601_ vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 team_02_WB.START_ADDR_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 team_02_WB.START_ADDR_VAL_REG\[0\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ net1129 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
Xhold94 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\] vssd1 vssd1
+ vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15601__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13803_ _03288_ net960 _03287_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__and3b_1
XFILLER_0_98_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14783_ net1186 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
X_11995_ net315 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\] net478 vssd1
+ vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11913__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15181__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16522_ clknet_leaf_30_wb_clk_i _02656_ _01329_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13734_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] _03242_ vssd1 vssd1 vccd1
+ vccd1 _03243_ sky130_fd_sc_hd__or2_1
X_10946_ _06270_ _06459_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16453_ clknet_leaf_65_wb_clk_i net1568 _01261_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dfrtp_1
X_13665_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\]
+ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__and3_1
X_10877_ net369 _06077_ _06391_ net399 vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08507__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ net2001 net283 net553 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15404_ clknet_leaf_25_wb_clk_i _01544_ _00212_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09075__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16384_ clknet_leaf_80_wb_clk_i _02519_ _01192_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ net1490 net963 _03148_ net1066 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09614__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15335_ clknet_leaf_104_wb_clk_i _01478_ _00148_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12547_ net266 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\] net444 vssd1
+ vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__mux2_1
XANTENNA__08822__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16107__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15266_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[25\]
+ _00079_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_12478_ net254 net2493 net560 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 _06626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13174__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14217_ net1099 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
X_11429_ net795 _06924_ _06917_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_39_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15197_ net1262 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14148_ net1126 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16257__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14079_ net1182 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
XANTENNA__07573__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire537_A _04801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1070 net61 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_2
X_08640_ _04268_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__inv_2
Xfanout1081 net1088 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__buf_2
XFILLER_0_83_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1092 net1097 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_2
XANTENNA__15281__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10160__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08571_ team_02_WB.instance_to_wrap.top.a1.row1\[61\] _04237_ _04225_ vssd1 vssd1
+ vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
X_16854__1398 vssd1 vssd1 vccd1 vccd1 _16854__1398/HI net1398 sky130_fd_sc_hd__conb_1
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11823__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15091__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09066__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09123_ _04633_ _04635_ _04637_ _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08813__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12654__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16782__1326 vssd1 vssd1 vccd1 vccd1 _16782__1326/HI net1326 sky130_fd_sc_hd__conb_1
XFILLER_0_5_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09054_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\] net758 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08005_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03689_ _03721_ vssd1 vssd1
+ vccd1 vccd1 _03728_ sky130_fd_sc_hd__nand3_1
XFILLER_0_124_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold520 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold531 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1226_A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold542 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold564 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold597 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09956_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\] net748 net712 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a22o_1
XANTENNA__12125__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08907_ net1527 _04435_ _04433_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__mux2_1
X_09887_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\] net886 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a22o_1
XANTENNA__11479__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ net1567 net1040 net1036 team_02_WB.instance_to_wrap.ramstore\[26\] vssd1
+ vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a22o_1
Xhold1242 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1275 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1286 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1297 team_02_WB.instance_to_wrap.ramload\[27\] vssd1 vssd1 vccd1 vccd1 net2755
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08769_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\] net742 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__a22o_1
XANTENNA__11733__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10800_ _04630_ net405 vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11780_ net270 net1967 net594 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09844__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ _04349_ _04354_ _04344_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__and3b_1
XANTENNA__07855__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13450_ _03044_ _03049_ _02768_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09057__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10662_ net996 _04421_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12401_ net337 net2170 net461 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_123_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08804__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ net2197 net1010 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[10\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12564__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ _04462_ _06109_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__nor2_4
X_15120_ net1230 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12332_ net327 net2182 net567 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10592__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15051_ net1220 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12263_ net314 net2333 net573 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__mux2_1
X_14002_ net1123 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11214_ _06351_ _06718_ _06717_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12194_ net308 net1830 net580 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11908__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ _06266_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15953_ clknet_leaf_22_wb_clk_i _02093_ _00761_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11076_ _06574_ _06581_ _06582_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__or3_1
X_16714__1273 vssd1 vssd1 vccd1 vccd1 _16714__1273/HI net1273 sky130_fd_sc_hd__conb_1
X_14904_ net1195 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
X_10027_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\] net831 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\]
+ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__a221o_1
X_15884_ clknet_leaf_20_wb_clk_i _02024_ _00692_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10142__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14835_ net1165 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09296__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14766_ net1114 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
X_11978_ net237 net2280 net478 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09835__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16505_ clknet_leaf_30_wb_clk_i _02639_ _01312_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13717_ _03204_ _03023_ net1065 _03200_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__and4b_1
X_10929_ net369 _06326_ net399 vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__o21ai_1
X_14697_ net1101 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09048__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16436_ clknet_leaf_103_wb_clk_i _02571_ _01244_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__dfrtp_1
X_13648_ team_02_WB.instance_to_wrap.top.lcd.lcd_rs net1066 _03023_ _03194_ vssd1
+ vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16367_ clknet_leaf_36_wb_clk_i _02507_ _01175_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13579_ team_02_WB.instance_to_wrap.top.a1.row1\[8\] _03110_ _03128_ team_02_WB.instance_to_wrap.top.a1.row1\[104\]
+ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15318_ clknet_leaf_120_wb_clk_i _01461_ _00131_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16298_ clknet_leaf_1_wb_clk_i _02438_ _01106_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15249_ clknet_leaf_63_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[8\]
+ _00062_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09220__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10905__A1 _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11818__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\] net926 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\]
+ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a221o_1
Xfanout307 _06891_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_1
XANTENNA__15086__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 net320 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_22_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout329 _03568_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_2
X_09741_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\] net707 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\]
+ _05254_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15797__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09672_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\] net810 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__a22o_1
XANTENNA__10133__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08623_ net103 net1572 net955 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__mux2_1
XANTENNA__12649__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout267_A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08554_ _04217_ _04218_ net653 net793 net1534 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09287__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08485_ _04179_ _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout434_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09039__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout601_A _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12384__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16422__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09106_ _04613_ _04614_ _04615_ _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09037_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\] net816 net897 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\]
+ _04548_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold350 team_02_WB.instance_to_wrap.ramload\[4\] vssd1 vssd1 vccd1 vccd1 net1808
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11728__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold394 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout830 net832 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_4
XANTENNA__10372__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout841 net842 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_6
Xfanout852 _03195_ vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09939_ _05449_ _05451_ _05453_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__or4_1
Xfanout863 _04543_ vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
Xfanout874 _04539_ vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_8
Xfanout885 _04537_ vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_4
Xfanout896 net897 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13310__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ team_02_WB.instance_to_wrap.top.pc\[15\] _06197_ vssd1 vssd1 vccd1 vccd1
+ _07470_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10124__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1050 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1
+ net2508 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__A1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11901_ net357 net2685 net486 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__mux2_1
Xhold1061 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ _07398_ _07400_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1094 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12559__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13244__A _06415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12786__C _06770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11832_ net342 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\] net591 vssd1
+ vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
X_14620_ net1146 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09278__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11690__C _07161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10587__B _04464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551_ net1172 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11763_ net332 net1947 net599 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13502_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__or2_1
X_10714_ _06174_ _06230_ _06175_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14482_ net1121 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11694_ _07130_ _07137_ _07179_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__nand3_1
XFILLER_0_125_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16221_ clknet_leaf_51_wb_clk_i _02361_ _01029_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13433_ _03040_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__inv_2
X_10645_ _06161_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__inv_2
XANTENNA__12294__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16152_ clknet_leaf_54_wb_clk_i _02292_ _00960_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13364_ team_02_WB.instance_to_wrap.ramload\[26\] net1016 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[26\] sky130_fd_sc_hd__and2_1
XFILLER_0_84_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10576_ _06090_ _06092_ net371 vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__mux2_1
XANTENNA__09450__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12315_ net257 net1946 net566 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__mux2_1
X_15103_ net1078 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
X_16083_ clknet_leaf_56_wb_clk_i _02223_ _00891_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13295_ team_02_WB.instance_to_wrap.top.pc\[12\] net1052 _06908_ net933 vssd1 vssd1
+ vccd1 vccd1 _02997_ sky130_fd_sc_hd__a22o_2
XFILLER_0_107_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16853__1397 vssd1 vssd1 vccd1 vccd1 _16853__1397/HI net1397 sky130_fd_sc_hd__conb_1
XFILLER_0_62_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15034_ net1200 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
X_12246_ net237 net2597 net573 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09202__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12177_ net646 _06278_ _06280_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_20_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11560__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ _06353_ _06633_ _06632_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13301__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ _06567_ _06568_ net415 vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__mux2_1
X_15936_ clknet_leaf_109_wb_clk_i _02076_ _00744_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10115__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11312__A1 _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16781__1325 vssd1 vssd1 vccd1 vccd1 _16781__1325/HI net1325 sky130_fd_sc_hd__conb_1
X_15867_ clknet_leaf_127_wb_clk_i _02007_ _00675_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12469__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13154__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13065__A1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14818_ net1205 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
XANTENNA__09269__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15798_ clknet_leaf_47_wb_clk_i _01938_ _00606_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12812__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14749_ net1084 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12812__B2 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ _03983_ _03985_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16419_ clknet_leaf_67_wb_clk_i _02554_ _01227_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09441__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10354__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07985_ _03695_ _03703_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__and2b_1
XFILLER_0_129_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout384_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\] net895 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10106__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__A0 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\] net763 net707 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12379__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08606_ net90 net1564 net955 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09261__B _04733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09586_ net529 vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08537_ _04171_ _04220_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout816_A _04521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08468_ net1606 net1006 net981 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1
+ vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a22o_1
XANTENNA__09680__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15812__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire516 _05439_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_2
X_08399_ _04090_ _04105_ _04106_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__or3_2
XFILLER_0_68_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire538 net540 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_85_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire549 net550 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
X_10430_ _04997_ _05946_ _04993_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__a21oi_1
X_16713__1272 vssd1 vssd1 vccd1 vccd1 _16713__1272/HI net1272 sky130_fd_sc_hd__conb_1
XFILLER_0_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10361_ net389 _05877_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__nor2_1
X_12100_ net1800 net334 net582 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__mux2_1
X_13080_ _07460_ _07524_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10292_ _05787_ _05807_ net968 vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__mux2_1
X_12031_ net322 net2690 net475 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold180 team_02_WB.instance_to_wrap.top.a1.row1\[9\] vssd1 vssd1 vccd1 vccd1 net1638
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10345__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16318__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout660 _06115_ vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__buf_2
Xfanout671 _05964_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16770_ net1314 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
Xfanout682 net685 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_4
Xfanout693 _04397_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_4
X_13982_ net1189 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XANTENNA__13295__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15721_ clknet_leaf_106_wb_clk_i _01861_ _00529_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12933_ team_02_WB.instance_to_wrap.top.pc\[26\] _06150_ vssd1 vssd1 vccd1 vccd1
+ _07453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12289__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13047__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15652_ clknet_leaf_1_wb_clk_i _01792_ _00460_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12864_ _05489_ _05491_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14603_ net1203 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
X_11815_ net280 net2146 net590 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12795_ _06102_ _07099_ _07317_ _07318_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__and4_1
X_15583_ clknet_leaf_55_wb_clk_i _01723_ _00391_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11921__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11746_ net260 net2531 net598 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14534_ net1074 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
XANTENNA__15492__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09671__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08735__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ _05125_ _05978_ _07162_ _05973_ _05124_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__a311o_1
X_14465_ net1211 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08515__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16204_ clknet_leaf_25_wb_clk_i _02344_ _01012_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10628_ team_02_WB.instance_to_wrap.top.pc\[27\] _06143_ vssd1 vssd1 vccd1 vccd1
+ _06145_ sky130_fd_sc_hd__and2_1
X_13416_ team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] team_02_WB.instance_to_wrap.top.lcd.currentState\[0\]
+ _03023_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__mux2_1
XANTENNA__09423__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14396_ net1149 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10569__C1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13347_ net1741 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[9\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09974__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16135_ clknet_leaf_27_wb_clk_i _02275_ _00943_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08777__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10559_ _04714_ net404 vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13278_ net1703 net986 net967 _02988_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__a22o_1
X_16066_ clknet_leaf_121_wb_clk_i _02206_ _00874_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15017_ net1233 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
X_12229_ net1874 net306 net616 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__mux2_1
XANTENNA__13149__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10336__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07770_ _03451_ _03491_ _03492_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__and3_1
XANTENNA__13286__A1 net1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13286__B2 _02992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15919_ clknet_leaf_36_wb_clk_i _02059_ _00727_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12199__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09440_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\] net766 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\]
+ _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09371_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\] net919 net891 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11831__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08322_ _04015_ _04028_ _04032_ _04024_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07610__A team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08253_ _03967_ _03968_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15985__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12549__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08184_ _03892_ _03894_ _03895_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_116_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13210__B2 _04946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12662__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10971__A _06084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1041_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10575__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout599_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10327__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09193__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_A _04372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07968_ _03648_ _03687_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__xor2_1
XANTENNA__10910__S net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13277__B2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09707_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\] net785 net713 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__a22o_1
X_07899_ _03595_ _03619_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout933_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_134_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09638_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\] net920 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\]
+ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16852__1396 vssd1 vssd1 vccd1 vccd1 _16852__1396/HI net1396 sky130_fd_sc_hd__conb_1
XFILLER_0_116_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09569_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\] net784 net760 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ net388 _07052_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11741__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12580_ net267 net2086 net439 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09653__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11531_ net417 _06635_ _06849_ net375 _07018_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14250_ net1138 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
X_11462_ _06007_ _06956_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_22_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09405__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13201_ _04564_ net936 net1020 net1561 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_123_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16780__1324 vssd1 vssd1 vccd1 vccd1 _16780__1324/HI net1324 sky130_fd_sc_hd__conb_1
X_10413_ _05927_ _05929_ _05420_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__o21a_1
XANTENNA__08759__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ net1093 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11393_ net2122 net304 net642 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XANTENNA__12572__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ net228 _02897_ _02900_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a21boi_1
XANTENNA_input62_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\] net765 _05859_ _05860_
+ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15708__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13063_ _07529_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10275_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\] net836 net881 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__a22o_1
XANTENNA__08070__B _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ net250 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\] net474 vssd1
+ vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
XANTENNA__09184__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16290__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11916__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16822_ net1366 vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__buf_2
XANTENNA__15184__A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 _07196_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_6
XFILLER_0_79_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16753_ net1297 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13965_ net1236 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15704_ clknet_leaf_19_wb_clk_i _01844_ _00512_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12916_ _04755_ _06147_ _07435_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16684_ clknet_leaf_73_wb_clk_i _02801_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_13896_ net1251 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09892__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15635_ clknet_leaf_56_wb_clk_i _01775_ _00443_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12847_ _05061_ _06186_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15566_ clknet_leaf_27_wb_clk_i _01706_ _00374_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12778_ _06720_ _06902_ _07299_ _07301_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09644__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14517_ net1216 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11729_ net331 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\] net602 vssd1
+ vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15497_ clknet_leaf_104_wb_clk_i _01637_ _00305_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14448_ net1077 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09947__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12482__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10791__A _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold905 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14379_ net1151 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold916 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
X_16118_ clknet_leaf_52_wb_clk_i _02258_ _00926_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold938 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold949 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15388__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ team_02_WB.instance_to_wrap.top.a1.instruction\[13\] _04278_ _04315_ vssd1
+ vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16049_ clknet_leaf_21_wb_clk_i _02189_ _00857_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16633__CLK clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10309__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__A2 _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ net26 net1030 net988 net1944 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07822_ _03506_ _03541_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__xor2_2
XANTENNA__15094__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11826__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10190__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09092__A _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _03457_ _03475_ _03460_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_105_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16712__1271 vssd1 vssd1 vccd1 vccd1 _16712__1271/HI net1271 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_101_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07684_ _03363_ _03368_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_101_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09423_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\] net863 net856 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\]
+ _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a221o_1
XANTENNA__16013__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10882__A2_N _06388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11561__S net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_A _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1089_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\] net840 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09635__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10245__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08305_ _03976_ _03993_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_60_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1197_A team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09285_ net536 vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__inv_2
XANTENNA__12785__A3 _06388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1256_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08236_ _03952_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__inv_2
XANTENNA__13195__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12392__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ _03879_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__nor2_2
XFILLER_0_71_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08098_ _03815_ _03816_ _03800_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a21boi_1
XANTENNA_fanout883_A _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09166__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10060_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\] net760 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11736__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13750_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] _03251_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__a21o_1
X_10962_ _06068_ _06094_ net393 vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09874__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ net352 net2512 net432 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12567__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13681_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\] _03198_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__a21oi_1
X_10893_ _05957_ net663 net659 _04653_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15420_ clknet_leaf_45_wb_clk_i _01560_ _00228_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12632_ net1891 net338 net553 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09626__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ net326 net1939 net443 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__mux2_1
X_15351_ clknet_leaf_87_wb_clk_i _01491_ _00164_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14302_ net1190 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _05604_ _06113_ _07006_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_81_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12494_ net312 net1984 net557 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__mux2_1
X_15282_ clknet_leaf_90_wb_clk_i _01426_ _00095_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ net374 _06747_ _06940_ net381 vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__a2bb2o_1
X_14233_ net1128 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
XANTENNA__15179__A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14164_ net1076 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11376_ net415 _06401_ _06853_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13115_ team_02_WB.instance_to_wrap.top.pc\[16\] net1024 _02886_ _07337_ vssd1 vssd1
+ vccd1 vccd1 _01497_ sky130_fd_sc_hd__a22o_1
X_10327_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\] net820 net808 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\]
+ _05843_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_128_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14095_ net1115 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _07451_ _07533_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__and2_1
XANTENNA__09157__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\] net841 net676 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\]
+ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_124_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1230 net1237 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1241 net1242 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__clkbuf_4
Xfanout1252 net1253 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__buf_4
X_10189_ _05699_ _05701_ _05703_ _05705_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__or4_1
Xfanout1263 net1264 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__buf_2
X_16805_ net1349 vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_2
X_14997_ net1221 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16736_ net1282 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13948_ net1210 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09865__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16667_ clknet_leaf_74_wb_clk_i _00017_ _01409_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.noisy
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12477__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ net1256 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15618_ clknet_leaf_124_wb_clk_i _01758_ _00426_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09617__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16598_ clknet_leaf_96_wb_clk_i _02717_ _01391_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15549_ clknet_leaf_51_wb_clk_i _01689_ _00357_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\] net770 _04583_ _04585_
+ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a2111o_2
XTAP_TAPCELL_ROW_96_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08021_ _03733_ _03737_ _03742_ _03712_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__a31o_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold702 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold724 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold735 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold746 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold768 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
X_16851__1395 vssd1 vssd1 vccd1 vccd1 _16851__1395/HI net1395 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold779 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__inv_2
XANTENNA__09148__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\] net958 vssd1 vssd1 vccd1
+ vccd1 _04444_ sky130_fd_sc_hd__or2_1
XANTENNA__08047__A2_N _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ net140 net1037 net1033 net1525 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10163__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1004_A _04259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07805_ _03481_ _03494_ net364 vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13056__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08785_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\] net726 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\]
+ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout464_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07736_ _03424_ _03458_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__nand2b_2
XANTENNA__11112__C1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07667_ _03388_ _03389_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__or2_1
XANTENNA__12387__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09406_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\] net739 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\]
+ _04922_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07598_ net2741 net1009 _03321_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09337_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\] net822 net875 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a22o_1
XANTENNA__15553__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09268_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\] net767 net747 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08219_ _03916_ _03918_ _03919_ _03926_ _03934_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__o41ai_1
XFILLER_0_16_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16533__D net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11331__A_N net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\] net833 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11179__C1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11230_ _06264_ _06734_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _04993_ net662 net659 _04995_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__a22oi_1
X_10112_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\] net901 net800 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\]
+ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a221o_1
XANTENNA__09139__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ _05976_ _06600_ _06022_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_8_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16059__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14920_ net1178 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10043_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\] net756 net744 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12789__C _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold40 team_02_WB.START_ADDR_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_02_WB.START_ADDR_VAL_REG\[22\] vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_02_WB.instance_to_wrap.ramaddr\[27\] vssd1 vssd1 vccd1 vccd1 net1520
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 net137 vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ net1145 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold84 team_02_WB.instance_to_wrap.top.a1.data\[8\] vssd1 vssd1 vccd1 vccd1 net1542
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1
+ net1553 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\]
+ _03284_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__and3_1
X_14782_ net1189 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
XANTENNA__09847__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11994_ net305 net2519 net478 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
XANTENNA__09311__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16521_ clknet_leaf_7_wb_clk_i _02655_ _01328_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13733_ _03242_ net949 _03241_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__and3b_1
X_10945_ team_02_WB.instance_to_wrap.top.pc\[27\] _06269_ team_02_WB.instance_to_wrap.top.pc\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12297__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ clknet_leaf_64_wb_clk_i net1475 _01260_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13664_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[2\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _03198_
+ sky130_fd_sc_hd__and3_1
X_16875__1419 vssd1 vssd1 vccd1 vccd1 _16875__1419/HI net1419 sky130_fd_sc_hd__conb_1
XFILLER_0_27_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10876_ net390 _06079_ _06080_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15403_ clknet_leaf_115_wb_clk_i _01543_ _00211_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12615_ net1746 net269 net553 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16383_ clknet_leaf_80_wb_clk_i _02518_ _01191_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _03112_ _03135_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15334_ clknet_leaf_64_wb_clk_i _01477_ _00147_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12546_ net256 net1778 net444 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15265_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[24\]
+ _00078_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_12477_ net239 net2133 net557 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__mux2_1
X_16711__1270 vssd1 vssd1 vccd1 vccd1 _16711__1270/HI net1270 sky130_fd_sc_hd__conb_1
XANTENNA__08523__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_4 _06657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14216_ net1176 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09378__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ net419 _06481_ _06922_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__a21o_1
X_15196_ net1260 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ _06201_ _06206_ _06208_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__nand3_1
X_14147_ net1131 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
XANTENNA_max_cap527_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14078_ net1189 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13029_ _07352_ _07440_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10145__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15426__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 net1061 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_2
XFILLER_0_98_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1071 net1079 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_4
XANTENNA__11893__A0 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1082 net1088 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__buf_4
Xfanout1093 net1097 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_4
XFILLER_0_117_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08570_ net1009 _04236_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09302__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11645__B1 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16719_ net1447 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15576__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11405__A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12000__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\] net809 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\]
+ _04638_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08813__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09053_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\] net754 net731 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08004_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03689_ _03721_ vssd1 vssd1
+ vccd1 vccd1 _03727_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold532 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12670__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold554 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1121_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1219_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09955_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\] net756 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout581_A _07209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout679_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08906_ net1045 _04190_ _04202_ net1008 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__a32o_1
XANTENNA__10136__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\] net918 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a22o_1
Xhold1210 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09541__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1232 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ net158 net1037 net1033 net1532 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
Xhold1243 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1254 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15919__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1265 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1287 team_02_WB.instance_to_wrap.top.a1.row1\[17\] vssd1 vssd1 vccd1 vccd1 net2745
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08768_ net847 _04365_ _04370_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__and3_4
Xhold1298 team_02_WB.instance_to_wrap.ramstore\[17\] vssd1 vssd1 vccd1 vccd1 net2756
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold257_A team_02_WB.instance_to_wrap.ramstore\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_135_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07719_ _03440_ _03441_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08699_ _04276_ _04320_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10730_ net994 net849 vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ team_02_WB.instance_to_wrap.top.pc\[22\] _06177_ vssd1 vssd1 vccd1 vccd1
+ _06178_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14626__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12400_ net332 net2600 net460 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13380_ net1741 net1010 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[9\]
+ sky130_fd_sc_hd__and2_1
X_10592_ _04463_ _04467_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ net322 net2388 net567 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11050__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15050_ net1200 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
X_12262_ net305 net2286 net573 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14001_ net1105 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
X_11213_ net410 _06480_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12580__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12193_ net302 net2112 net578 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15449__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ team_02_WB.instance_to_wrap.top.pc\[21\] _06265_ team_02_WB.instance_to_wrap.top.pc\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09780__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13313__B1 _07083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15952_ clknet_leaf_34_wb_clk_i _02092_ _00760_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11075_ _04865_ _06026_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10127__B1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14903_ net1174 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
X_10026_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\] net904 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09532__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15599__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ clknet_leaf_117_wb_clk_i _02023_ _00691_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11924__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14834_ net1121 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14765_ net1147 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11977_ net247 net2742 net478 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ clknet_leaf_5_wb_clk_i _02638_ _01311_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13716_ net1695 _03231_ _03232_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10928_ net390 _06315_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__nor2_1
X_16850__1394 vssd1 vssd1 vccd1 vccd1 _16850__1394/HI net1394 sky130_fd_sc_hd__conb_1
XFILLER_0_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14696_ net1176 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16435_ clknet_leaf_64_wb_clk_i net1702 _01243_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09048__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13647_ _03289_ _03114_ _03115_ _03193_ _03023_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__a311oi_1
X_10859_ _04693_ _05956_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09599__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16366_ clknet_leaf_27_wb_clk_i _02506_ _01174_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13578_ team_02_WB.instance_to_wrap.top.a1.row1\[56\] _03117_ _03119_ team_02_WB.instance_to_wrap.top.a1.row1\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15317_ clknet_leaf_105_wb_clk_i _01460_ _00130_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12529_ net323 net2187 net448 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__mux2_1
XANTENNA__10602__B2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16297_ clknet_leaf_119_wb_clk_i _02437_ _01105_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15248_ clknet_leaf_61_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[7\]
+ _00061_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08079__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12490__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10366__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ net1238 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XANTENNA__10905__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout308 net311 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_2
XANTENNA__09771__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15204__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13304__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09740_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\] net755 net727 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__a22o_1
XANTENNA__10118__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
.ends

