* NGSPICE file created from SRAM_1024x32_wb_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for EF_SRAM_1024x32 abstract view
.subckt EF_SRAM_1024x32 DO[16] BEN[16] DO[17] BEN[17] DO[18] BEN[18] DO[19] BEN[19]
+ DO[20] BEN[20] DO[21] BEN[21] DO[22] BEN[22] DO[23] BEN[23] DO[24] BEN[24] DO[25]
+ BEN[25] DO[26] BEN[26] DO[27] BEN[27] DO[28] BEN[28] DO[29] BEN[29] DO[30] BEN[30]
+ DO[31] BEN[31] AD[0] AD[1] AD[2] WLBI WLOFF CLKin EN R_WB SM TM ScanInDR ScanOutCC
+ ScanInDL DO[9] BEN[9] DO[10] BEN[10] DO[11] BEN[11] DO[12] BEN[12] DO[13] BEN[13]
+ DO[14] BEN[14] DO[15] BEN[15] BEN[8] AD[3] AD[4] AD[5] AD[6] AD[7] AD[8] AD[9] ScanInCC
+ DO[0] BEN[0] DO[1] BEN[1] DO[2] BEN[2] DO[3] BEN[3] DO[4] BEN[4] DO[5] BEN[5] DO[6]
+ BEN[6] DO[7] BEN[7] DO[8] DI[3] DI[12] DI[0] DI[4] DI[14] DI[11] DI[5] DI[1] DI[9]
+ DI[6] DI[15] DI[2] DI[7] DI[13] DI[10] DI[8] DI[23] DI[27] DI[19] DI[21] DI[28]
+ DI[24] DI[18] DI[29] DI[16] DI[25] DI[30] DI[22] DI[20] DI[26] DI[17] DI[31] vnb
+ vpwrm vpwra vpwrp vgnd vpb vpwrpc vpwrac
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt SRAM_1024x32_wb_wrapper VGND VPWR wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XPHY_EDGE_ROW_95_2_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_127_2_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_2_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_2_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_2_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_2_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_2_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_136_2_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_2_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_2_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold30 net36 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 net25 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 net201 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 net224 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 net7 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 wbs_sel_i[3] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 net179 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_2_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput75 net75 VGND VGND VPWR VPWR wbs_dat_o[30] sky130_fd_sc_hd__buf_12
Xoutput64 net64 VGND VGND VPWR VPWR wbs_dat_o[20] sky130_fd_sc_hd__buf_12
Xoutput53 net53 VGND VGND VPWR VPWR wbs_dat_o[10] sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_144_2_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_25_2_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_2_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_108_2_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_2_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_152_2_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_2_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_153_2_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold42 net22 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 wbs_cyc_i VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 net222 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 net208 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 net228 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 net46 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_12
Xhold20 net44 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 net10 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_154_2_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_2_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput76 net76 VGND VGND VPWR VPWR wbs_dat_o[31] sky130_fd_sc_hd__buf_12
Xoutput65 net65 VGND VGND VPWR VPWR wbs_dat_o[21] sky130_fd_sc_hd__buf_12
Xoutput54 net54 VGND VGND VPWR VPWR wbs_dat_o[11] sky130_fd_sc_hd__buf_12
XFILLER_0_129_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_2_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_155_2_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_2_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_2_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_2_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_2_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_2_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_2_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_2_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_2_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold32 net37 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 net32 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 net26 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 net204 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 net214 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 net192 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 wbs_we_i VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 wbs_sel_i[1] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 net6 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_2_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_2_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_2_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_2_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_154_2_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_2_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_2_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput66 net66 VGND VGND VPWR VPWR wbs_dat_o[22] sky130_fd_sc_hd__buf_12
Xoutput55 net55 VGND VGND VPWR VPWR wbs_dat_o[12] sky130_fd_sc_hd__buf_12
Xoutput77 net77 VGND VGND VPWR VPWR wbs_dat_o[3] sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_12_2_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_2_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_2_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_2_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_2_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_2_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold140 wbs_adr_i[0] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_2_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_2_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_2_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_2_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_2_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_2_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_2_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_2_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSRAM_0 net59 net184 net60 net184 net61 net184 net62 net184 net64 net184 net65 net184
+ net66 net184 net67 net184 net68 net187 net69 net187 net70 net187 net71 net187 net72
+ net187 net73 net187 net75 net187 net76 net187 net176 net174 net172 net84 net85 clknet_1_1__leaf_wb_clk_i
+ ram_controller.EN ram_controller.R_WB net86 net87 net88 SRAM_0/ScanOutCC net89 net83
+ net178 net53 net178 net54 net178 net55 net178 net56 net178 net57 net178 net58 net178
+ net178 net170 net168 net166 net164 net160 net156 net150 net90 net52 net181 net63
+ net181 net74 net181 net77 net181 net78 net181 net79 net181 net80 net181 net81 net181
+ net82 net158 net128 net110 net140 net114 net94 net132 net106 net112 net130 net96
+ net100 net126 net118 net104 net120 net152 net102 net138 net146 net108 net154 net134
+ net116 net142 net162 net122 net148 net144 net98 net136 net124 VGND VPWR VPWR VPWR
+ VGND VPWR net91 net92 EF_SRAM_1024x32
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_2_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_2_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_2_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_2_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_2_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold11 net196 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 net18 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_37_2_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold44 net21 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 net206 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 net182 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 wbs_dat_i[15] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 net229 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 net199 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 net38 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_33_2_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_2_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_2_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_2_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput67 net67 VGND VGND VPWR VPWR wbs_dat_o[23] sky130_fd_sc_hd__buf_12
Xoutput56 net56 VGND VGND VPWR VPWR wbs_dat_o[13] sky130_fd_sc_hd__buf_12
Xoutput78 net78 VGND VGND VPWR VPWR wbs_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_0_152_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_2_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_2_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_2_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold130 wbs_dat_i[31] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_2_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_2_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 clknet_1_0__leaf_wb_clk_i VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_100_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_2_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold56 net27 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 net220 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 net205 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 net42 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 net14 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 net225 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 net5 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 net45 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_12
XFILLER_0_39_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput57 net57 VGND VGND VPWR VPWR wbs_dat_o[14] sky130_fd_sc_hd__buf_12
Xoutput68 net68 VGND VGND VPWR VPWR wbs_dat_o[24] sky130_fd_sc_hd__buf_12
Xoutput79 net79 VGND VGND VPWR VPWR wbs_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_0_35_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_2_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_153_2_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold131 wbs_adr_i[9] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 wbs_dat_i[2] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_2_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_2_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_94_2_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_140_2_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold24 net34 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 net23 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 net230 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 net194 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 net223 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 net217 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 net9 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_102_2_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_141_2_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput69 net69 VGND VGND VPWR VPWR wbs_dat_o[25] sky130_fd_sc_hd__buf_12
Xoutput58 net58 VGND VGND VPWR VPWR wbs_dat_o[15] sky130_fd_sc_hd__buf_12
XFILLER_0_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_106_2_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_2_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_2_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_2_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_2_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold110 wbs_dat_i[5] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold132 wbs_adr_i[8] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 wbs_dat_i[26] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_2_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_2_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_106_2_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold69 net215 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 net193 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 net209 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 net24 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 net16 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 net11 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_107_2_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput59 net59 VGND VGND VPWR VPWR wbs_dat_o[16] sky130_fd_sc_hd__buf_12
XFILLER_0_67_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_108_2_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_2_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold100 wbs_dat_i[14] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 wbs_dat_i[20] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 wbs_adr_i[7] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 wbs_dat_i[3] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_2_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_2_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_152_2_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_2_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold15 net218 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 net210 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 net200 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 net39 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 net17 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_2_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_2_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_2_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold123 wbs_dat_i[25] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 wbs_dat_i[17] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 wbs_dat_i[13] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 wbs_adr_i[6] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_105_2_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_2_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_91_2_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold16 net33 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 net198 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold38 net41 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 net207 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold102 wbs_dat_i[12] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 wbs_dat_i[27] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold113 wbs_dat_i[19] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 wbs_adr_i[5] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_1_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_2_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_2_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_2_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_2_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold17 net219 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 net202 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 net43 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_2_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Left_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_2_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_2_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold114 wbs_dat_i[22] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 wbs_adr_i[4] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 wbs_dat_i[11] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 wbs_dat_i[1] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_2_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_36_2_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold29 net221 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 net13 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_90_2_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_2_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold115 wbs_dat_i[16] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 wbs_dat_i[10] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 wbs_dat_i[28] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold137 wbs_adr_i[3] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_2_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold19 net197 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_2_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_2_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_150_2_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_2_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_150_2_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_2_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_2_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_2_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold127 wbs_dat_i[0] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 wbs_dat_i[21] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 wbs_dat_i[9] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 wbs_adr_i[2] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_151_2_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_2_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_2_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_2_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_2_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_2_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_2_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_2_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_2_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_2_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_2_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_115_2_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_2_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 wb_rst_i VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_2_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_2_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_2_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_2_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_2_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_2_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_2_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_2_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_2_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_2_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_2_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_2_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_2_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold117 wbs_dat_i[4] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 wbs_dat_i[29] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 wbs_dat_i[8] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 wbs_adr_i[1] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_2_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_2_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_2_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_2_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_2_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_119_2_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_2_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_2_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_2_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_2_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 net175 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_68_2_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_2_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_2_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_2_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_2_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_2_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_2_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold107 wbs_dat_i[7] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 wbs_dat_i[30] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 wbs_dat_i[23] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_144_2_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_2_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_2_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_2_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput3 net173 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XFILLER_0_47_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_90_2_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput50 net190 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_2_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold108 wbs_dat_i[6] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold119 wbs_dat_i[24] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_2_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_2_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 net171 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_4
XFILLER_0_149_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6_ clknet_1_0__leaf_wb_clk_i _0_ _1_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput40 net131 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_2_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_2_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_2_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold109 wbs_dat_i[18] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_2_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_2_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_143_2_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_2_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_2_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 net169 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_0_70_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5_ net51 net12 net49 VGND VGND VPWR VPWR _0_ sky130_fd_sc_hd__and3b_1
XFILLER_0_139_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_89_2_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 net161 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
Xinput41 net129 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_2_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_2_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 net167 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_4
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4_ net12 net49 VGND VGND VPWR VPWR ram_controller.EN sky130_fd_sc_hd__and2_4
XFILLER_0_84_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_124_2_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_2_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_2_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput20 net141 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput31 net97 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_4
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 net125 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_2_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_2_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_2_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_2_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_123_2_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 net165 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_4
XFILLER_0_55_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSRAM_0_90 VGND VGND VPWR VPWR SRAM_0_90/HI net90 sky130_fd_sc_hd__conb_1
X_3_ net1 VGND VGND VPWR VPWR _1_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_142_2_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_124_2_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_79_2_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_2_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput32 net101 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
Xinput21 net135 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_4
Xinput43 net119 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
Xinput10 net155 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_4
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_2_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_2_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_2_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_88_2_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_127_2_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_2_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_2_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_2_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 net163 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_4
XFILLER_0_47_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_2_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_2_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XSRAM_0_91 VGND VGND VPWR VPWR net91 SRAM_0_91/LO sky130_fd_sc_hd__conb_1
X_2_ net50 VGND VGND VPWR VPWR ram_controller.R_WB sky130_fd_sc_hd__clkinv_4
XFILLER_0_52_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput22 net133 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
Xinput11 net149 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_4
Xinput33 net107 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_4
Xinput44 net111 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_123_2_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_2_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_148_2_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_2_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_2_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 net159 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_4
XFILLER_0_87_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XSRAM_0_92 VGND VGND VPWR VPWR net92 SRAM_0_92/LO sky130_fd_sc_hd__conb_1
XFILLER_0_154_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput34 net115 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_4
Xinput23 net137 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
Xinput45 net180 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_12
Xinput12 net189 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_21_2_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_141_2_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_2_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_2_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1 net195 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_104_2_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_2_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_2_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_2_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_2_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_2_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 net109 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_4
XFILLER_0_142_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput35 net99 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_4
Xinput46 net177 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_12
Xinput24 net105 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_4
XFILLER_0_25_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_2_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2 net15 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_62_2_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_2_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_2_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_2_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_2_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_2_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_147_2_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_2_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_111_2_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_79_2_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_2_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_2_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_2_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput36 net121 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_4
Xinput25 net143 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
Xinput14 net103 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_2_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput47 net183 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_12
XFILLER_0_118_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_2_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_2_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_2_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_88_2_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_140_2_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 net191 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_62_2_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_2_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_2_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_2_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XSRAM_0_84 VGND VGND VPWR VPWR SRAM_0_84/HI net84 sky130_fd_sc_hd__conb_1
XFILLER_0_139_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_2_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_2_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_86_2_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput37 net123 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_4
Xinput26 net145 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
Xinput48 net186 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_12
Xinput15 net93 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_112_2_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_2_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_2_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold4 net19 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_2_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_121_2_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_2_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_2_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XSRAM_0_85 VGND VGND VPWR VPWR SRAM_0_85/HI net85 sky130_fd_sc_hd__conb_1
XFILLER_0_139_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_2_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput16 net127 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
Xinput49 wbs_stb_i VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_1
Xinput27 net147 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
Xinput38 net157 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_2_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_134_2_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_2_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_130_2_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_2_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_2_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_0_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_2_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold5 net213 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_2_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_155_2_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_87_2_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_2_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_2_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSRAM_0_86 VGND VGND VPWR VPWR SRAM_0_86/HI net86 sky130_fd_sc_hd__conb_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_2_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_2_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_102_2_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput28 net151 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
Xinput17 net117 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
Xinput39 net139 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_2_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_139_2_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_2_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_96_2_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_85_2_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 net31 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_2_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_111_2_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_2_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_2_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_2_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_2_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSRAM_0_87 VGND VGND VPWR VPWR SRAM_0_87/HI net87 sky130_fd_sc_hd__conb_1
XFILLER_0_139_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_2_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_2_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_2_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_2_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 net113 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
Xinput29 net153 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_2_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 net212 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_145_2_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_2_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_2_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSRAM_0_88 VGND VGND VPWR VPWR SRAM_0_88/HI net88 sky130_fd_sc_hd__conb_1
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_2_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_2_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_2_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_2_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput19 net95 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_2_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_101_2_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_2_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 net35 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_33_2_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_95_2_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_2_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_2_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_110_2_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSRAM_0_89 VGND VGND VPWR VPWR SRAM_0_89/HI net89 sky130_fd_sc_hd__conb_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_2_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_2_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_2_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_2_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_2_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_121_2_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_2_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_2_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold9 net216 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_7_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_2_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_139_2_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_2_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_2_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_2_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_2_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_2_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_2_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_2_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_2_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_2_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_2_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_2_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_2_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold90 wbs_sel_i[0] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput80 net80 VGND VGND VPWR VPWR wbs_dat_o[6] sky130_fd_sc_hd__buf_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_2_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_142_2_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_2_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_2_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_143_2_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_2_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_2_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_2_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_55_2_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_2_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_145_2_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold80 net4 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 net185 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_2_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_2_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput70 net70 VGND VGND VPWR VPWR wbs_dat_o[26] sky130_fd_sc_hd__buf_12
Xoutput81 net81 VGND VGND VPWR VPWR wbs_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_0_144_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_2_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_2_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_138_2_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_2_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_147_2_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_2_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_1_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_2_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_2_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_2_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_2_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_2_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_2_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold70 net30 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 net47 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_12
Xhold81 net231 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_2_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput71 net71 VGND VGND VPWR VPWR wbs_dat_o[27] sky130_fd_sc_hd__buf_12
Xoutput60 net60 VGND VGND VPWR VPWR wbs_dat_o[17] sky130_fd_sc_hd__buf_12
Xoutput82 net82 VGND VGND VPWR VPWR wbs_dat_o[8] sky130_fd_sc_hd__buf_12
XPHY_EDGE_ROW_36_2_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_2_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_2_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_1_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_150_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_119_2_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_56_2_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_2_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_2_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold60 net28 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 net3 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 net226 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 wbs_sel_i[2] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_2_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_65_2_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_2_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput72 net72 VGND VGND VPWR VPWR wbs_dat_o[28] sky130_fd_sc_hd__buf_12
Xoutput61 net61 VGND VGND VPWR VPWR wbs_dat_o[18] sky130_fd_sc_hd__buf_12
Xoutput83 net83 VGND VGND VPWR VPWR wbs_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_0_144_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_2_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_137_2_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_2_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_63_2_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_26_2_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold50 net20 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 net211 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 net232 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 net188 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_21_2_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold72 net8 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_2_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput73 net73 VGND VGND VPWR VPWR wbs_dat_o[29] sky130_fd_sc_hd__buf_12
Xoutput62 net62 VGND VGND VPWR VPWR wbs_dat_o[19] sky130_fd_sc_hd__buf_12
Xoutput51 net51 VGND VGND VPWR VPWR wbs_ack_o sky130_fd_sc_hd__buf_12
XFILLER_0_129_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_2_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_2_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_2_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_2_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_130_2_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_2_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_2_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_2_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_2_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_2_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_44_2_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold40 net40 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 net48 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_12
Xhold62 net29 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 net203 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 net227 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 net2 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_94_2_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput52 net52 VGND VGND VPWR VPWR wbs_dat_o[0] sky130_fd_sc_hd__buf_12
XPHY_EDGE_ROW_4_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput63 net63 VGND VGND VPWR VPWR wbs_dat_o[1] sky130_fd_sc_hd__buf_12
Xoutput74 net74 VGND VGND VPWR VPWR wbs_dat_o[2] sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_152_2_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

