magic
tech sky130A
magscale 1 2
timestamp 1720829860
<< viali >>
rect 38853 37417 38887 37451
rect 45569 37417 45603 37451
rect 46673 37417 46707 37451
rect 44189 37349 44223 37383
rect 36277 37213 36311 37247
rect 40509 37213 40543 37247
rect 40785 37213 40819 37247
rect 39129 37145 39163 37179
rect 44005 37145 44039 37179
rect 45293 37145 45327 37179
rect 46581 37145 46615 37179
rect 35725 37077 35759 37111
rect 35633 36873 35667 36907
rect 40325 36873 40359 36907
rect 40693 36873 40727 36907
rect 41153 36873 41187 36907
rect 41797 36873 41831 36907
rect 42625 36873 42659 36907
rect 42901 36873 42935 36907
rect 45201 36873 45235 36907
rect 45661 36873 45695 36907
rect 46121 36873 46155 36907
rect 46949 36873 46983 36907
rect 47685 36873 47719 36907
rect 48237 36873 48271 36907
rect 48973 36873 49007 36907
rect 49433 36873 49467 36907
rect 50169 36873 50203 36907
rect 50813 36873 50847 36907
rect 51457 36873 51491 36907
rect 52101 36873 52135 36907
rect 52837 36873 52871 36907
rect 53481 36873 53515 36907
rect 53941 36873 53975 36907
rect 54585 36873 54619 36907
rect 55229 36873 55263 36907
rect 55873 36873 55907 36907
rect 56609 36873 56643 36907
rect 57253 36873 57287 36907
rect 57989 36873 58023 36907
rect 58541 36873 58575 36907
rect 59185 36873 59219 36907
rect 59921 36873 59955 36907
rect 60473 36873 60507 36907
rect 61209 36873 61243 36907
rect 61669 36873 61703 36907
rect 62405 36873 62439 36907
rect 63233 36873 63267 36907
rect 63693 36873 63727 36907
rect 64337 36873 64371 36907
rect 64981 36873 65015 36907
rect 65625 36873 65659 36907
rect 66269 36873 66303 36907
rect 66913 36873 66947 36907
rect 67557 36873 67591 36907
rect 68385 36873 68419 36907
rect 68845 36873 68879 36907
rect 69489 36873 69523 36907
rect 70133 36873 70167 36907
rect 70777 36873 70811 36907
rect 71421 36873 71455 36907
rect 72065 36873 72099 36907
rect 72525 36873 72559 36907
rect 72893 36873 72927 36907
rect 36705 36805 36739 36839
rect 36921 36805 36955 36839
rect 45385 36805 45419 36839
rect 32873 36737 32907 36771
rect 33149 36737 33183 36771
rect 35725 36737 35759 36771
rect 35909 36737 35943 36771
rect 40509 36737 40543 36771
rect 40877 36737 40911 36771
rect 41337 36737 41371 36771
rect 41429 36737 41463 36771
rect 41981 36737 42015 36771
rect 42073 36737 42107 36771
rect 42441 36737 42475 36771
rect 43085 36737 43119 36771
rect 45017 36737 45051 36771
rect 45845 36737 45879 36771
rect 45937 36737 45971 36771
rect 47133 36737 47167 36771
rect 47225 36737 47259 36771
rect 47869 36737 47903 36771
rect 48421 36737 48455 36771
rect 48513 36737 48547 36771
rect 48789 36737 48823 36771
rect 49617 36737 49651 36771
rect 49709 36737 49743 36771
rect 50353 36737 50387 36771
rect 50445 36737 50479 36771
rect 50997 36737 51031 36771
rect 51089 36737 51123 36771
rect 51641 36737 51675 36771
rect 51733 36737 51767 36771
rect 52285 36737 52319 36771
rect 52377 36737 52411 36771
rect 53021 36737 53055 36771
rect 53297 36737 53331 36771
rect 54125 36737 54159 36771
rect 54217 36737 54251 36771
rect 54769 36737 54803 36771
rect 54861 36737 54895 36771
rect 55413 36737 55447 36771
rect 55505 36737 55539 36771
rect 56057 36737 56091 36771
rect 56149 36737 56183 36771
rect 56793 36737 56827 36771
rect 56885 36737 56919 36771
rect 57437 36737 57471 36771
rect 57529 36737 57563 36771
rect 58173 36737 58207 36771
rect 58725 36737 58759 36771
rect 58817 36737 58851 36771
rect 59369 36737 59403 36771
rect 59461 36737 59495 36771
rect 60105 36737 60139 36771
rect 60657 36737 60691 36771
rect 61025 36737 61059 36771
rect 61853 36737 61887 36771
rect 61945 36737 61979 36771
rect 62589 36737 62623 36771
rect 62681 36737 62715 36771
rect 63049 36737 63083 36771
rect 63877 36737 63911 36771
rect 63969 36737 64003 36771
rect 64521 36737 64555 36771
rect 64613 36737 64647 36771
rect 65165 36737 65199 36771
rect 65257 36737 65291 36771
rect 65809 36737 65843 36771
rect 65901 36737 65935 36771
rect 66453 36737 66487 36771
rect 66545 36737 66579 36771
rect 67097 36737 67131 36771
rect 67189 36737 67223 36771
rect 67741 36737 67775 36771
rect 67833 36737 67867 36771
rect 68201 36737 68235 36771
rect 69029 36737 69063 36771
rect 69121 36737 69155 36771
rect 69673 36737 69707 36771
rect 69765 36737 69799 36771
rect 70317 36737 70351 36771
rect 70409 36737 70443 36771
rect 70961 36737 70995 36771
rect 71053 36737 71087 36771
rect 71605 36737 71639 36771
rect 71697 36737 71731 36771
rect 72249 36737 72283 36771
rect 72709 36737 72743 36771
rect 73077 36737 73111 36771
rect 73629 36737 73663 36771
rect 2053 36669 2087 36703
rect 32229 36669 32263 36703
rect 33241 36669 33275 36703
rect 33885 36669 33919 36703
rect 34161 36669 34195 36703
rect 38209 36669 38243 36703
rect 38485 36669 38519 36703
rect 43177 36669 43211 36703
rect 43453 36669 43487 36703
rect 46213 36669 46247 36703
rect 60749 36669 60783 36703
rect 73353 36669 73387 36703
rect 36553 36601 36587 36635
rect 33425 36533 33459 36567
rect 35909 36533 35943 36567
rect 36737 36533 36771 36567
rect 39957 36533 39991 36567
rect 44925 36533 44959 36567
rect 2329 36329 2363 36363
rect 32045 36329 32079 36363
rect 34989 36329 35023 36363
rect 35633 36329 35667 36363
rect 38761 36329 38795 36363
rect 39681 36329 39715 36363
rect 42533 36329 42567 36363
rect 43085 36329 43119 36363
rect 43545 36329 43579 36363
rect 43729 36329 43763 36363
rect 44373 36329 44407 36363
rect 44649 36329 44683 36363
rect 47777 36329 47811 36363
rect 48789 36329 48823 36363
rect 52929 36329 52963 36363
rect 53297 36329 53331 36363
rect 58081 36329 58115 36363
rect 60657 36329 60691 36363
rect 61025 36329 61059 36363
rect 63141 36329 63175 36363
rect 68293 36329 68327 36363
rect 72249 36329 72283 36363
rect 34713 36261 34747 36295
rect 35909 36261 35943 36295
rect 2513 36193 2547 36227
rect 33517 36193 33551 36227
rect 33793 36193 33827 36227
rect 36185 36193 36219 36227
rect 36461 36193 36495 36227
rect 42257 36193 42291 36227
rect 46305 36193 46339 36227
rect 2053 36125 2087 36159
rect 2145 36125 2179 36159
rect 34989 36125 35023 36159
rect 35173 36125 35207 36159
rect 35909 36125 35943 36159
rect 36093 36125 36127 36159
rect 38577 36125 38611 36159
rect 38945 36125 38979 36159
rect 39221 36125 39255 36159
rect 39313 36125 39347 36159
rect 44097 36125 44131 36159
rect 44189 36125 44223 36159
rect 46121 36125 46155 36159
rect 46397 36125 46431 36159
rect 39497 36057 39531 36091
rect 41981 36057 42015 36091
rect 1869 35989 1903 36023
rect 33977 35989 34011 36023
rect 37933 35989 37967 36023
rect 38025 35989 38059 36023
rect 39129 35989 39163 36023
rect 40509 35989 40543 36023
rect 43729 35989 43763 36023
rect 45937 35989 45971 36023
rect 32781 35785 32815 35819
rect 36093 35785 36127 35819
rect 36369 35785 36403 35819
rect 36829 35785 36863 35819
rect 38393 35785 38427 35819
rect 40785 35785 40819 35819
rect 41537 35785 41571 35819
rect 41705 35785 41739 35819
rect 44373 35785 44407 35819
rect 47317 35785 47351 35819
rect 32321 35717 32355 35751
rect 36645 35717 36679 35751
rect 37013 35717 37047 35751
rect 41337 35717 41371 35751
rect 45845 35717 45879 35751
rect 2053 35649 2087 35683
rect 2145 35649 2179 35683
rect 31769 35649 31803 35683
rect 32137 35649 32171 35683
rect 32505 35649 32539 35683
rect 32597 35649 32631 35683
rect 32781 35649 32815 35683
rect 36277 35649 36311 35683
rect 36461 35649 36495 35683
rect 36737 35649 36771 35683
rect 38209 35649 38243 35683
rect 38393 35649 38427 35683
rect 40601 35649 40635 35683
rect 40785 35649 40819 35683
rect 40877 35649 40911 35683
rect 41061 35649 41095 35683
rect 44557 35649 44591 35683
rect 44741 35649 44775 35683
rect 44833 35649 44867 35683
rect 31953 35581 31987 35615
rect 45569 35581 45603 35615
rect 37013 35513 37047 35547
rect 1869 35445 1903 35479
rect 31585 35445 31619 35479
rect 41245 35445 41279 35479
rect 41521 35445 41555 35479
rect 47685 35445 47719 35479
rect 34713 35241 34747 35275
rect 45201 35241 45235 35275
rect 45845 35241 45879 35275
rect 28457 35105 28491 35139
rect 28733 35105 28767 35139
rect 31493 35105 31527 35139
rect 36277 35105 36311 35139
rect 28365 35037 28399 35071
rect 29561 35037 29595 35071
rect 30113 35037 30147 35071
rect 31217 35037 31251 35071
rect 34989 35037 35023 35071
rect 35173 35037 35207 35071
rect 35541 35037 35575 35071
rect 36553 35037 36587 35071
rect 43361 35037 43395 35071
rect 43545 35037 43579 35071
rect 43637 35037 43671 35071
rect 44005 35037 44039 35071
rect 44557 35037 44591 35071
rect 45661 35037 45695 35071
rect 46029 35037 46063 35071
rect 46121 35037 46155 35071
rect 45385 34969 45419 35003
rect 2053 34901 2087 34935
rect 32965 34901 32999 34935
rect 34897 34901 34931 34935
rect 35449 34901 35483 34935
rect 43177 34901 43211 34935
rect 45017 34901 45051 34935
rect 45185 34901 45219 34935
rect 1869 34697 1903 34731
rect 36277 34697 36311 34731
rect 45115 34697 45149 34731
rect 28733 34629 28767 34663
rect 42717 34629 42751 34663
rect 45201 34629 45235 34663
rect 2053 34561 2087 34595
rect 28457 34561 28491 34595
rect 32413 34561 32447 34595
rect 33517 34561 33551 34595
rect 36185 34561 36219 34595
rect 36369 34561 36403 34595
rect 37933 34561 37967 34595
rect 39037 34561 39071 34595
rect 42441 34561 42475 34595
rect 45017 34561 45051 34595
rect 45293 34561 45327 34595
rect 2145 34493 2179 34527
rect 30849 34493 30883 34527
rect 32321 34493 32355 34527
rect 32505 34493 32539 34527
rect 32597 34493 32631 34527
rect 35265 34493 35299 34527
rect 35449 34493 35483 34527
rect 36093 34493 36127 34527
rect 30297 34425 30331 34459
rect 30205 34357 30239 34391
rect 32137 34357 32171 34391
rect 33780 34357 33814 34391
rect 37289 34357 37323 34391
rect 39300 34357 39334 34391
rect 40785 34357 40819 34391
rect 44189 34357 44223 34391
rect 38117 34153 38151 34187
rect 39313 34153 39347 34187
rect 39497 34153 39531 34187
rect 41337 34153 41371 34187
rect 43361 34153 43395 34187
rect 1869 34085 1903 34119
rect 29101 34085 29135 34119
rect 30205 34017 30239 34051
rect 31953 34017 31987 34051
rect 35725 34017 35759 34051
rect 36277 34017 36311 34051
rect 43177 34017 43211 34051
rect 2053 33949 2087 33983
rect 26985 33949 27019 33983
rect 28825 33949 28859 33983
rect 28917 33949 28951 33983
rect 32321 33949 32355 33983
rect 32413 33949 32447 33983
rect 34897 33949 34931 33983
rect 35081 33949 35115 33983
rect 35541 33949 35575 33983
rect 36001 33949 36035 33983
rect 36093 33949 36127 33983
rect 36369 33949 36403 33983
rect 38945 33949 38979 33983
rect 40233 33949 40267 33983
rect 40877 33949 40911 33983
rect 41153 33949 41187 33983
rect 43637 33949 43671 33983
rect 27261 33881 27295 33915
rect 29101 33881 29135 33915
rect 30481 33881 30515 33915
rect 32597 33881 32631 33915
rect 34989 33881 35023 33915
rect 35265 33881 35299 33915
rect 36277 33881 36311 33915
rect 36645 33881 36679 33915
rect 39313 33881 39347 33915
rect 39865 33881 39899 33915
rect 40049 33881 40083 33915
rect 28733 33813 28767 33847
rect 32045 33813 32079 33847
rect 32229 33813 32263 33847
rect 34713 33813 34747 33847
rect 35357 33813 35391 33847
rect 40969 33813 41003 33847
rect 43545 33813 43579 33847
rect 45109 33813 45143 33847
rect 28365 33609 28399 33643
rect 28825 33609 28859 33643
rect 29561 33609 29595 33643
rect 30389 33609 30423 33643
rect 40325 33609 40359 33643
rect 40493 33609 40527 33643
rect 41981 33609 42015 33643
rect 44465 33609 44499 33643
rect 46121 33609 46155 33643
rect 29724 33541 29758 33575
rect 29929 33541 29963 33575
rect 32781 33541 32815 33575
rect 39833 33541 39867 33575
rect 40049 33541 40083 33575
rect 40693 33541 40727 33575
rect 41153 33541 41187 33575
rect 45109 33541 45143 33575
rect 2053 33473 2087 33507
rect 2145 33473 2179 33507
rect 28273 33473 28307 33507
rect 28457 33473 28491 33507
rect 30849 33473 30883 33507
rect 32321 33473 32355 33507
rect 32505 33473 32539 33507
rect 35449 33473 35483 33507
rect 35633 33473 35667 33507
rect 36369 33473 36403 33507
rect 36553 33473 36587 33507
rect 38117 33473 38151 33507
rect 38393 33473 38427 33507
rect 38577 33473 38611 33507
rect 38945 33473 38979 33507
rect 40785 33473 40819 33507
rect 41521 33473 41555 33507
rect 41797 33473 41831 33507
rect 42165 33473 42199 33507
rect 42441 33473 42475 33507
rect 42717 33473 42751 33507
rect 44281 33473 44315 33507
rect 44649 33473 44683 33507
rect 44833 33473 44867 33507
rect 46305 33473 46339 33507
rect 46397 33473 46431 33507
rect 46581 33473 46615 33507
rect 46673 33473 46707 33507
rect 46949 33473 46983 33507
rect 29469 33405 29503 33439
rect 35541 33405 35575 33439
rect 39589 33405 39623 33439
rect 42533 33405 42567 33439
rect 45937 33405 45971 33439
rect 47777 33405 47811 33439
rect 48053 33405 48087 33439
rect 1869 33337 1903 33371
rect 30573 33337 30607 33371
rect 41337 33337 41371 33371
rect 42901 33337 42935 33371
rect 29745 33269 29779 33303
rect 32137 33269 32171 33303
rect 32689 33269 32723 33303
rect 36553 33269 36587 33303
rect 37933 33269 37967 33303
rect 39681 33269 39715 33303
rect 39865 33269 39899 33303
rect 40509 33269 40543 33303
rect 41153 33269 41187 33303
rect 41797 33269 41831 33303
rect 42441 33269 42475 33303
rect 44649 33269 44683 33303
rect 47041 33269 47075 33303
rect 49525 33269 49559 33303
rect 49709 33269 49743 33303
rect 32045 33065 32079 33099
rect 33701 33065 33735 33099
rect 37013 33065 37047 33099
rect 37381 33065 37415 33099
rect 39313 33065 39347 33099
rect 40877 33065 40911 33099
rect 43821 33065 43855 33099
rect 45201 33065 45235 33099
rect 46581 33065 46615 33099
rect 47961 33065 47995 33099
rect 32413 32997 32447 33031
rect 39221 32997 39255 33031
rect 45017 32997 45051 33031
rect 46397 32997 46431 33031
rect 30297 32929 30331 32963
rect 33057 32929 33091 32963
rect 33609 32929 33643 32963
rect 37473 32929 37507 32963
rect 37749 32929 37783 32963
rect 39681 32929 39715 32963
rect 42625 32929 42659 32963
rect 44097 32929 44131 32963
rect 46305 32929 46339 32963
rect 48053 32929 48087 32963
rect 49893 32929 49927 32963
rect 2053 32861 2087 32895
rect 2145 32861 2179 32895
rect 28273 32861 28307 32895
rect 28457 32861 28491 32895
rect 28641 32861 28675 32895
rect 29193 32861 29227 32895
rect 32045 32861 32079 32895
rect 32137 32861 32171 32895
rect 33701 32861 33735 32895
rect 33977 32861 34011 32895
rect 34069 32861 34103 32895
rect 35663 32861 35697 32895
rect 35817 32861 35851 32895
rect 37013 32861 37047 32895
rect 37105 32861 37139 32895
rect 39497 32861 39531 32895
rect 44189 32861 44223 32895
rect 44649 32861 44683 32895
rect 45293 32861 45327 32895
rect 45569 32861 45603 32895
rect 45820 32861 45854 32895
rect 47041 32861 47075 32895
rect 47225 32861 47259 32895
rect 47317 32861 47351 32895
rect 47501 32861 47535 32895
rect 47593 32861 47627 32895
rect 47685 32861 47719 32895
rect 29561 32793 29595 32827
rect 42349 32793 42383 32827
rect 43729 32793 43763 32827
rect 45937 32793 45971 32827
rect 46765 32793 46799 32827
rect 47133 32793 47167 32827
rect 48329 32793 48363 32827
rect 1869 32725 1903 32759
rect 28365 32725 28399 32759
rect 33885 32725 33919 32759
rect 34161 32725 34195 32759
rect 35449 32725 35483 32759
rect 39957 32725 39991 32759
rect 44373 32725 44407 32759
rect 44557 32725 44591 32759
rect 45661 32725 45695 32759
rect 46029 32725 46063 32759
rect 46565 32725 46599 32759
rect 49801 32725 49835 32759
rect 30297 32521 30331 32555
rect 32505 32521 32539 32555
rect 45201 32521 45235 32555
rect 46213 32521 46247 32555
rect 47593 32521 47627 32555
rect 18981 32453 19015 32487
rect 33977 32453 34011 32487
rect 45369 32453 45403 32487
rect 45569 32453 45603 32487
rect 45845 32453 45879 32487
rect 46061 32453 46095 32487
rect 48053 32453 48087 32487
rect 17141 32385 17175 32419
rect 26985 32385 27019 32419
rect 29009 32385 29043 32419
rect 29745 32385 29779 32419
rect 30113 32385 30147 32419
rect 31033 32385 31067 32419
rect 31125 32385 31159 32419
rect 31309 32385 31343 32419
rect 34253 32385 34287 32419
rect 34345 32385 34379 32419
rect 43729 32385 43763 32419
rect 44097 32385 44131 32419
rect 44465 32385 44499 32419
rect 44649 32385 44683 32419
rect 47777 32385 47811 32419
rect 48237 32385 48271 32419
rect 48329 32385 48363 32419
rect 2053 32317 2087 32351
rect 17417 32317 17451 32351
rect 27261 32317 27295 32351
rect 28733 32317 28767 32351
rect 29193 32317 29227 32351
rect 29653 32317 29687 32351
rect 30389 32317 30423 32351
rect 34621 32317 34655 32351
rect 36093 32317 36127 32351
rect 36737 32317 36771 32351
rect 47961 32317 47995 32351
rect 48053 32317 48087 32351
rect 43545 32249 43579 32283
rect 18889 32181 18923 32215
rect 28825 32181 28859 32215
rect 29377 32181 29411 32215
rect 30021 32181 30055 32215
rect 31125 32181 31159 32215
rect 36185 32181 36219 32215
rect 45385 32181 45419 32215
rect 46029 32181 46063 32215
rect 1869 31977 1903 32011
rect 17141 31977 17175 32011
rect 27997 31977 28031 32011
rect 29837 31977 29871 32011
rect 31413 31977 31447 32011
rect 34713 31977 34747 32011
rect 35081 31977 35115 32011
rect 44005 31977 44039 32011
rect 46305 31977 46339 32011
rect 46489 31977 46523 32011
rect 43894 31909 43928 31943
rect 44373 31909 44407 31943
rect 16681 31841 16715 31875
rect 21465 31841 21499 31875
rect 31677 31841 31711 31875
rect 35173 31841 35207 31875
rect 44097 31841 44131 31875
rect 2053 31773 2087 31807
rect 12081 31773 12115 31807
rect 15393 31773 15427 31807
rect 15577 31773 15611 31807
rect 16773 31773 16807 31807
rect 17877 31773 17911 31807
rect 18521 31773 18555 31807
rect 27813 31773 27847 31807
rect 27997 31773 28031 31807
rect 29561 31773 29595 31807
rect 29837 31773 29871 31807
rect 34897 31773 34931 31807
rect 37289 31773 37323 31807
rect 43729 31773 43763 31807
rect 12357 31705 12391 31739
rect 14197 31705 14231 31739
rect 20637 31705 20671 31739
rect 21649 31705 21683 31739
rect 29653 31705 29687 31739
rect 46121 31705 46155 31739
rect 46337 31705 46371 31739
rect 2145 31637 2179 31671
rect 13829 31637 13863 31671
rect 15485 31637 15519 31671
rect 29929 31637 29963 31671
rect 37473 31637 37507 31671
rect 1869 31433 1903 31467
rect 12357 31433 12391 31467
rect 17509 31433 17543 31467
rect 29811 31433 29845 31467
rect 30849 31433 30883 31467
rect 40709 31433 40743 31467
rect 41061 31433 41095 31467
rect 15025 31365 15059 31399
rect 30021 31365 30055 31399
rect 36737 31365 36771 31399
rect 36953 31365 36987 31399
rect 40049 31365 40083 31399
rect 40509 31365 40543 31399
rect 45109 31365 45143 31399
rect 45385 31365 45419 31399
rect 45845 31365 45879 31399
rect 46857 31365 46891 31399
rect 2053 31297 2087 31331
rect 14749 31297 14783 31331
rect 17693 31297 17727 31331
rect 27813 31297 27847 31331
rect 28549 31297 28583 31331
rect 29193 31297 29227 31331
rect 39773 31297 39807 31331
rect 39957 31297 39991 31331
rect 40233 31297 40267 31331
rect 40969 31297 41003 31331
rect 41153 31297 41187 31331
rect 41521 31297 41555 31331
rect 41705 31297 41739 31331
rect 42533 31297 42567 31331
rect 44741 31297 44775 31331
rect 45569 31297 45603 31331
rect 45753 31297 45787 31331
rect 46029 31297 46063 31331
rect 46581 31297 46615 31331
rect 46673 31297 46707 31331
rect 46949 31297 46983 31331
rect 47133 31297 47167 31331
rect 9597 31229 9631 31263
rect 9873 31229 9907 31263
rect 11345 31229 11379 31263
rect 12081 31229 12115 31263
rect 13369 31229 13403 31263
rect 14105 31229 14139 31263
rect 17233 31229 17267 31263
rect 17969 31229 18003 31263
rect 19441 31229 19475 31263
rect 20085 31229 20119 31263
rect 27721 31229 27755 31263
rect 31401 31229 31435 31263
rect 38761 31229 38795 31263
rect 39037 31229 39071 31263
rect 46213 31229 46247 31263
rect 46857 31229 46891 31263
rect 29653 31161 29687 31195
rect 37105 31161 37139 31195
rect 39865 31161 39899 31195
rect 41337 31161 41371 31195
rect 11529 31093 11563 31127
rect 12817 31093 12851 31127
rect 13553 31093 13587 31127
rect 16497 31093 16531 31127
rect 16681 31093 16715 31127
rect 19533 31093 19567 31127
rect 20361 31093 20395 31127
rect 27445 31093 27479 31127
rect 29837 31093 29871 31127
rect 36921 31093 36955 31127
rect 37289 31093 37323 31127
rect 40325 31093 40359 31127
rect 40693 31093 40727 31127
rect 40877 31093 40911 31127
rect 43085 31093 43119 31127
rect 45109 31093 45143 31127
rect 45293 31093 45327 31127
rect 46949 31093 46983 31127
rect 10977 30889 11011 30923
rect 12173 30889 12207 30923
rect 15485 30889 15519 30923
rect 18521 30889 18555 30923
rect 29101 30889 29135 30923
rect 31585 30889 31619 30923
rect 37289 30889 37323 30923
rect 37841 30889 37875 30923
rect 40693 30889 40727 30923
rect 41613 30889 41647 30923
rect 46765 30889 46799 30923
rect 48697 30889 48731 30923
rect 17417 30821 17451 30855
rect 31401 30821 31435 30855
rect 11345 30753 11379 30787
rect 11713 30753 11747 30787
rect 17601 30753 17635 30787
rect 27353 30753 27387 30787
rect 27629 30753 27663 30787
rect 43361 30753 43395 30787
rect 45017 30753 45051 30787
rect 46949 30753 46983 30787
rect 47225 30753 47259 30787
rect 2053 30685 2087 30719
rect 2145 30685 2179 30719
rect 10977 30685 11011 30719
rect 11161 30685 11195 30719
rect 11253 30685 11287 30719
rect 11437 30685 11471 30719
rect 11805 30685 11839 30719
rect 15209 30685 15243 30719
rect 15485 30685 15519 30719
rect 17141 30685 17175 30719
rect 17417 30685 17451 30719
rect 18245 30685 18279 30719
rect 18337 30685 18371 30719
rect 18521 30685 18555 30719
rect 31585 30685 31619 30719
rect 31953 30685 31987 30719
rect 32045 30685 32079 30719
rect 34253 30685 34287 30719
rect 37473 30685 37507 30719
rect 37749 30685 37783 30719
rect 37841 30685 37875 30719
rect 38117 30685 38151 30719
rect 40601 30685 40635 30719
rect 33977 30617 34011 30651
rect 36277 30617 36311 30651
rect 36461 30617 36495 30651
rect 37933 30617 37967 30651
rect 43085 30617 43119 30651
rect 45293 30617 45327 30651
rect 1869 30549 1903 30583
rect 15301 30549 15335 30583
rect 17233 30549 17267 30583
rect 30665 30549 30699 30583
rect 32505 30549 32539 30583
rect 36093 30549 36127 30583
rect 37657 30549 37691 30583
rect 43729 30549 43763 30583
rect 48789 30549 48823 30583
rect 13093 30345 13127 30379
rect 15961 30345 15995 30379
rect 17601 30345 17635 30379
rect 43085 30345 43119 30379
rect 44373 30345 44407 30379
rect 12449 30277 12483 30311
rect 12633 30277 12667 30311
rect 13277 30277 13311 30311
rect 14013 30277 14047 30311
rect 15761 30277 15795 30311
rect 17509 30277 17543 30311
rect 30665 30277 30699 30311
rect 32505 30277 32539 30311
rect 36093 30277 36127 30311
rect 36309 30277 36343 30311
rect 36645 30277 36679 30311
rect 37381 30277 37415 30311
rect 37933 30277 37967 30311
rect 40693 30277 40727 30311
rect 44097 30277 44131 30311
rect 44741 30277 44775 30311
rect 2053 30209 2087 30243
rect 2145 30209 2179 30243
rect 11805 30209 11839 30243
rect 11897 30209 11931 30243
rect 12541 30209 12575 30243
rect 13001 30209 13035 30243
rect 13375 30209 13409 30243
rect 13553 30209 13587 30243
rect 17233 30209 17267 30243
rect 17417 30209 17451 30243
rect 18429 30209 18463 30243
rect 18613 30209 18647 30243
rect 18797 30209 18831 30243
rect 29377 30209 29411 30243
rect 29561 30209 29595 30243
rect 29837 30209 29871 30243
rect 30205 30209 30239 30243
rect 31585 30209 31619 30243
rect 32137 30209 32171 30243
rect 32321 30209 32355 30243
rect 33149 30209 33183 30243
rect 34253 30209 34287 30243
rect 36553 30209 36587 30243
rect 36737 30209 36771 30243
rect 42809 30209 42843 30243
rect 42901 30209 42935 30243
rect 43637 30209 43671 30243
rect 44557 30209 44591 30243
rect 14565 30141 14599 30175
rect 19349 30141 19383 30175
rect 29653 30141 29687 30175
rect 31217 30141 31251 30175
rect 31677 30141 31711 30175
rect 32229 30141 32263 30175
rect 34529 30141 34563 30175
rect 39221 30141 39255 30175
rect 40969 30141 41003 30175
rect 42441 30141 42475 30175
rect 43453 30141 43487 30175
rect 11621 30073 11655 30107
rect 12265 30073 12299 30107
rect 12817 30073 12851 30107
rect 13369 30073 13403 30107
rect 16129 30073 16163 30107
rect 30021 30073 30055 30107
rect 1869 30005 1903 30039
rect 13277 30005 13311 30039
rect 15945 30005 15979 30039
rect 17785 30005 17819 30039
rect 18429 30005 18463 30039
rect 29561 30005 29595 30039
rect 30481 30005 30515 30039
rect 31861 30005 31895 30039
rect 36001 30005 36035 30039
rect 36277 30005 36311 30039
rect 36461 30005 36495 30039
rect 37473 30005 37507 30039
rect 43821 30005 43855 30039
rect 44833 30005 44867 30039
rect 46949 30005 46983 30039
rect 11621 29801 11655 29835
rect 15485 29801 15519 29835
rect 15853 29801 15887 29835
rect 17693 29801 17727 29835
rect 17877 29801 17911 29835
rect 18797 29801 18831 29835
rect 22293 29801 22327 29835
rect 31309 29801 31343 29835
rect 34713 29801 34747 29835
rect 37749 29801 37783 29835
rect 18613 29733 18647 29767
rect 34897 29733 34931 29767
rect 8953 29665 8987 29699
rect 10701 29665 10735 29699
rect 11345 29665 11379 29699
rect 15301 29665 15335 29699
rect 19993 29665 20027 29699
rect 20453 29665 20487 29699
rect 20545 29665 20579 29699
rect 29561 29665 29595 29699
rect 32413 29665 32447 29699
rect 35173 29665 35207 29699
rect 36277 29665 36311 29699
rect 42257 29665 42291 29699
rect 15117 29597 15151 29631
rect 15577 29597 15611 29631
rect 16037 29597 16071 29631
rect 16221 29597 16255 29631
rect 18337 29597 18371 29631
rect 18797 29597 18831 29631
rect 18889 29597 18923 29631
rect 19073 29597 19107 29631
rect 19257 29597 19291 29631
rect 19441 29597 19475 29631
rect 20085 29597 20119 29631
rect 36001 29597 36035 29631
rect 9229 29529 9263 29563
rect 17509 29529 17543 29563
rect 17714 29529 17748 29563
rect 17969 29529 18003 29563
rect 18153 29529 18187 29563
rect 20821 29529 20855 29563
rect 29837 29529 29871 29563
rect 37841 29529 37875 29563
rect 38577 29529 38611 29563
rect 42533 29529 42567 29563
rect 44281 29529 44315 29563
rect 2053 29461 2087 29495
rect 10793 29461 10827 29495
rect 14933 29461 14967 29495
rect 18245 29461 18279 29495
rect 18521 29461 18555 29495
rect 19349 29461 19383 29495
rect 31861 29461 31895 29495
rect 38853 29461 38887 29495
rect 1869 29257 1903 29291
rect 10793 29257 10827 29291
rect 12173 29257 12207 29291
rect 14749 29257 14783 29291
rect 18981 29257 19015 29291
rect 21833 29257 21867 29291
rect 30113 29257 30147 29291
rect 32137 29257 32171 29291
rect 39405 29257 39439 29291
rect 42625 29257 42659 29291
rect 42993 29257 43027 29291
rect 13185 29189 13219 29223
rect 20453 29189 20487 29223
rect 41429 29189 41463 29223
rect 43545 29189 43579 29223
rect 2053 29121 2087 29155
rect 10701 29121 10735 29155
rect 10885 29121 10919 29155
rect 10977 29121 11011 29155
rect 11161 29121 11195 29155
rect 11529 29121 11563 29155
rect 11897 29121 11931 29155
rect 11989 29121 12023 29155
rect 15393 29121 15427 29155
rect 15577 29121 15611 29155
rect 16681 29121 16715 29155
rect 20729 29121 20763 29155
rect 22385 29121 22419 29155
rect 30021 29121 30055 29155
rect 30205 29121 30239 29155
rect 31585 29121 31619 29155
rect 33885 29121 33919 29155
rect 38292 29121 38326 29155
rect 40049 29121 40083 29155
rect 40877 29121 40911 29155
rect 40969 29121 41003 29155
rect 44097 29121 44131 29155
rect 45661 29121 45695 29155
rect 46121 29121 46155 29155
rect 46305 29121 46339 29155
rect 48237 29121 48271 29155
rect 48513 29121 48547 29155
rect 2145 29053 2179 29087
rect 11069 29053 11103 29087
rect 12909 29053 12943 29087
rect 14657 29053 14691 29087
rect 20913 29053 20947 29087
rect 31677 29053 31711 29087
rect 31953 29053 31987 29087
rect 33609 29053 33643 29087
rect 38025 29053 38059 29087
rect 41153 29053 41187 29087
rect 43085 29053 43119 29087
rect 43269 29053 43303 29087
rect 44189 29053 44223 29087
rect 45753 29053 45787 29087
rect 46029 29053 46063 29087
rect 44465 28985 44499 29019
rect 11989 28917 12023 28951
rect 15485 28917 15519 28951
rect 16773 28917 16807 28951
rect 39497 28917 39531 28951
rect 40509 28917 40543 28951
rect 46489 28917 46523 28951
rect 48329 28917 48363 28951
rect 48605 28917 48639 28951
rect 10701 28713 10735 28747
rect 10885 28713 10919 28747
rect 11713 28713 11747 28747
rect 14565 28713 14599 28747
rect 15853 28713 15887 28747
rect 16129 28713 16163 28747
rect 20821 28713 20855 28747
rect 38301 28713 38335 28747
rect 39129 28713 39163 28747
rect 1869 28645 1903 28679
rect 11161 28645 11195 28679
rect 13645 28645 13679 28679
rect 20453 28645 20487 28679
rect 20637 28645 20671 28679
rect 42717 28645 42751 28679
rect 46305 28645 46339 28679
rect 46673 28645 46707 28679
rect 13277 28577 13311 28611
rect 36369 28577 36403 28611
rect 39865 28577 39899 28611
rect 40141 28577 40175 28611
rect 41889 28577 41923 28611
rect 47501 28577 47535 28611
rect 49249 28577 49283 28611
rect 2053 28509 2087 28543
rect 9505 28509 9539 28543
rect 11529 28509 11563 28543
rect 12541 28509 12575 28543
rect 14381 28509 14415 28543
rect 14565 28509 14599 28543
rect 15301 28509 15335 28543
rect 15393 28509 15427 28543
rect 15577 28509 15611 28543
rect 17417 28509 17451 28543
rect 20177 28509 20211 28543
rect 36737 28509 36771 28543
rect 38577 28509 38611 28543
rect 38669 28509 38703 28543
rect 38761 28509 38795 28543
rect 38945 28509 38979 28543
rect 42441 28509 42475 28543
rect 42809 28509 42843 28543
rect 42901 28509 42935 28543
rect 43361 28509 43395 28543
rect 43453 28509 43487 28543
rect 46029 28509 46063 28543
rect 46397 28509 46431 28543
rect 46489 28509 46523 28543
rect 49525 28509 49559 28543
rect 10869 28441 10903 28475
rect 11069 28441 11103 28475
rect 11345 28441 11379 28475
rect 15669 28441 15703 28475
rect 15885 28441 15919 28475
rect 16313 28441 16347 28475
rect 16497 28441 16531 28475
rect 20269 28441 20303 28475
rect 20453 28441 20487 28475
rect 20789 28441 20823 28475
rect 21005 28441 21039 28475
rect 46121 28441 46155 28475
rect 46305 28441 46339 28475
rect 46673 28441 46707 28475
rect 10149 28373 10183 28407
rect 11437 28373 11471 28407
rect 14749 28373 14783 28407
rect 16037 28373 16071 28407
rect 16773 28373 16807 28407
rect 38163 28373 38197 28407
rect 42533 28373 42567 28407
rect 43177 28373 43211 28407
rect 49709 28373 49743 28407
rect 8401 28169 8435 28203
rect 18429 28169 18463 28203
rect 20269 28169 20303 28203
rect 20637 28169 20671 28203
rect 41981 28169 42015 28203
rect 45845 28169 45879 28203
rect 48329 28169 48363 28203
rect 9873 28101 9907 28135
rect 10241 28101 10275 28135
rect 11069 28101 11103 28135
rect 14933 28101 14967 28135
rect 16957 28101 16991 28135
rect 19993 28101 20027 28135
rect 45477 28101 45511 28135
rect 46397 28101 46431 28135
rect 2053 28033 2087 28067
rect 2145 28033 2179 28067
rect 10517 28033 10551 28067
rect 10609 28033 10643 28067
rect 10701 28033 10735 28067
rect 10885 28033 10919 28067
rect 10977 28033 11011 28067
rect 13093 28033 13127 28067
rect 15485 28033 15519 28067
rect 15669 28033 15703 28067
rect 15761 28033 15795 28067
rect 15853 28033 15887 28067
rect 20177 28033 20211 28067
rect 20361 28033 20395 28067
rect 21189 28033 21223 28067
rect 41153 28033 41187 28067
rect 43269 28033 43303 28067
rect 44097 28033 44131 28067
rect 44190 28033 44224 28067
rect 45937 28033 45971 28067
rect 47869 28033 47903 28067
rect 47961 28033 47995 28067
rect 10149 27965 10183 27999
rect 13369 27965 13403 27999
rect 16681 27965 16715 27999
rect 32873 27965 32907 27999
rect 33241 27965 33275 27999
rect 34805 27965 34839 27999
rect 35173 27965 35207 27999
rect 41245 27965 41279 27999
rect 43085 27965 43119 27999
rect 43177 27965 43211 27999
rect 44465 27965 44499 27999
rect 47685 27965 47719 27999
rect 1869 27897 1903 27931
rect 45109 27897 45143 27931
rect 45661 27897 45695 27931
rect 46213 27897 46247 27931
rect 14841 27829 14875 27863
rect 16129 27829 16163 27863
rect 18613 27829 18647 27863
rect 20545 27829 20579 27863
rect 34667 27829 34701 27863
rect 36599 27829 36633 27863
rect 43453 27829 43487 27863
rect 45477 27829 45511 27863
rect 46029 27829 46063 27863
rect 46121 27829 46155 27863
rect 47409 27829 47443 27863
rect 10793 27625 10827 27659
rect 16116 27625 16150 27659
rect 17601 27625 17635 27659
rect 33885 27625 33919 27659
rect 35173 27625 35207 27659
rect 36645 27625 36679 27659
rect 43085 27625 43119 27659
rect 12909 27557 12943 27591
rect 35633 27557 35667 27591
rect 44005 27557 44039 27591
rect 12449 27489 12483 27523
rect 15853 27489 15887 27523
rect 20545 27489 20579 27523
rect 34345 27489 34379 27523
rect 37105 27489 37139 27523
rect 37841 27489 37875 27523
rect 42625 27489 42659 27523
rect 2053 27421 2087 27455
rect 2145 27421 2179 27455
rect 10977 27421 11011 27455
rect 11161 27421 11195 27455
rect 12541 27421 12575 27455
rect 14105 27421 14139 27455
rect 14657 27421 14691 27455
rect 19441 27421 19475 27455
rect 19717 27421 19751 27455
rect 19901 27421 19935 27455
rect 19993 27421 20027 27455
rect 22477 27421 22511 27455
rect 34069 27421 34103 27455
rect 34161 27421 34195 27455
rect 34437 27421 34471 27455
rect 35357 27421 35391 27455
rect 35449 27421 35483 27455
rect 35725 27421 35759 27455
rect 36829 27421 36863 27455
rect 36921 27421 36955 27455
rect 37197 27421 37231 27455
rect 38209 27421 38243 27455
rect 42717 27421 42751 27455
rect 43085 27421 43119 27455
rect 43361 27421 43395 27455
rect 43545 27421 43579 27455
rect 43637 27421 43671 27455
rect 43730 27421 43764 27455
rect 45845 27421 45879 27455
rect 22201 27353 22235 27387
rect 1869 27285 1903 27319
rect 17693 27285 17727 27319
rect 19257 27285 19291 27319
rect 20729 27285 20763 27319
rect 22661 27285 22695 27319
rect 36461 27285 36495 27319
rect 39635 27285 39669 27319
rect 43269 27285 43303 27319
rect 45937 27285 45971 27319
rect 10317 27081 10351 27115
rect 10701 27081 10735 27115
rect 19993 27081 20027 27115
rect 20545 27081 20579 27115
rect 31953 27081 31987 27115
rect 35265 27081 35299 27115
rect 36921 27081 36955 27115
rect 38117 27081 38151 27115
rect 46029 27081 46063 27115
rect 10517 27013 10551 27047
rect 18521 27013 18555 27047
rect 36277 27013 36311 27047
rect 36553 27013 36587 27047
rect 42993 27013 43027 27047
rect 10793 26945 10827 26979
rect 11713 26945 11747 26979
rect 12265 26945 12299 26979
rect 12449 26945 12483 26979
rect 12541 26945 12575 26979
rect 12633 26945 12667 26979
rect 14749 26945 14783 26979
rect 20453 26945 20487 26979
rect 20637 26945 20671 26979
rect 35449 26945 35483 26979
rect 35541 26945 35575 26979
rect 35633 26945 35667 26979
rect 35817 26945 35851 26979
rect 36369 26945 36403 26979
rect 36645 26945 36679 26979
rect 36737 26945 36771 26979
rect 38301 26945 38335 26979
rect 38393 26945 38427 26979
rect 38669 26945 38703 26979
rect 39681 26945 39715 26979
rect 42441 26945 42475 26979
rect 42901 26945 42935 26979
rect 43085 26945 43119 26979
rect 43637 26945 43671 26979
rect 44189 26945 44223 26979
rect 45937 26945 45971 26979
rect 2053 26877 2087 26911
rect 11805 26877 11839 26911
rect 11897 26877 11931 26911
rect 11989 26877 12023 26911
rect 12909 26877 12943 26911
rect 14473 26877 14507 26911
rect 18245 26877 18279 26911
rect 32137 26877 32171 26911
rect 32505 26877 32539 26911
rect 36001 26877 36035 26911
rect 39957 26877 39991 26911
rect 41705 26877 41739 26911
rect 42717 26877 42751 26911
rect 43361 26877 43395 26911
rect 44557 26877 44591 26911
rect 44649 26877 44683 26911
rect 44741 26877 44775 26911
rect 44833 26877 44867 26911
rect 45017 26877 45051 26911
rect 48513 26877 48547 26911
rect 48789 26877 48823 26911
rect 50353 26877 50387 26911
rect 50629 26877 50663 26911
rect 54217 26877 54251 26911
rect 54493 26877 54527 26911
rect 11529 26809 11563 26843
rect 42533 26809 42567 26843
rect 44189 26809 44223 26843
rect 10149 26741 10183 26775
rect 10333 26741 10367 26775
rect 13001 26741 13035 26775
rect 18153 26741 18187 26775
rect 33931 26741 33965 26775
rect 35081 26741 35115 26775
rect 38577 26741 38611 26775
rect 42625 26741 42659 26775
rect 50261 26741 50295 26775
rect 52101 26741 52135 26775
rect 52745 26741 52779 26775
rect 1869 26537 1903 26571
rect 11805 26537 11839 26571
rect 11989 26537 12023 26571
rect 12357 26537 12391 26571
rect 20361 26537 20395 26571
rect 31033 26537 31067 26571
rect 32229 26537 32263 26571
rect 32689 26537 32723 26571
rect 34713 26537 34747 26571
rect 40417 26537 40451 26571
rect 41245 26537 41279 26571
rect 45845 26537 45879 26571
rect 49157 26537 49191 26571
rect 49617 26537 49651 26571
rect 53573 26537 53607 26571
rect 54033 26537 54067 26571
rect 45017 26469 45051 26503
rect 45477 26469 45511 26503
rect 9965 26401 9999 26435
rect 11713 26401 11747 26435
rect 20269 26401 20303 26435
rect 35357 26401 35391 26435
rect 41061 26401 41095 26435
rect 46397 26401 46431 26435
rect 48789 26401 48823 26435
rect 50721 26401 50755 26435
rect 52377 26401 52411 26435
rect 2053 26333 2087 26367
rect 12265 26333 12299 26367
rect 12449 26333 12483 26367
rect 20085 26333 20119 26367
rect 21925 26333 21959 26367
rect 30757 26333 30791 26367
rect 30849 26333 30883 26367
rect 31125 26333 31159 26367
rect 32125 26333 32159 26367
rect 32413 26333 32447 26367
rect 32505 26333 32539 26367
rect 34897 26333 34931 26367
rect 35265 26333 35299 26367
rect 40785 26333 40819 26367
rect 44097 26333 44131 26367
rect 44281 26333 44315 26367
rect 44649 26333 44683 26367
rect 44833 26333 44867 26367
rect 45293 26333 45327 26367
rect 45385 26333 45419 26367
rect 45569 26333 45603 26367
rect 45753 26333 45787 26367
rect 45970 26333 46004 26367
rect 46489 26333 46523 26367
rect 49341 26333 49375 26367
rect 49433 26333 49467 26367
rect 49709 26333 49743 26367
rect 50169 26333 50203 26367
rect 50905 26333 50939 26367
rect 51089 26333 51123 26367
rect 51273 26333 51307 26367
rect 52745 26333 52779 26367
rect 53389 26333 53423 26367
rect 53481 26333 53515 26367
rect 53757 26333 53791 26367
rect 53849 26333 53883 26367
rect 10241 26265 10275 26299
rect 11973 26265 12007 26299
rect 12173 26265 12207 26299
rect 20361 26265 20395 26299
rect 34989 26265 35023 26299
rect 35081 26265 35115 26299
rect 44465 26265 44499 26299
rect 46095 26265 46129 26299
rect 46765 26265 46799 26299
rect 48513 26265 48547 26299
rect 51181 26265 51215 26299
rect 51641 26265 51675 26299
rect 19901 26197 19935 26231
rect 21373 26197 21407 26231
rect 30573 26197 30607 26231
rect 40877 26197 40911 26231
rect 44741 26197 44775 26231
rect 51457 26197 51491 26231
rect 1869 25993 1903 26027
rect 15761 25993 15795 26027
rect 17877 25993 17911 26027
rect 31769 25993 31803 26027
rect 32413 25993 32447 26027
rect 37841 25993 37875 26027
rect 38577 25993 38611 26027
rect 40877 25993 40911 26027
rect 42901 25993 42935 26027
rect 46581 25993 46615 26027
rect 47961 25993 47995 26027
rect 48329 25993 48363 26027
rect 49893 25993 49927 26027
rect 51089 25993 51123 26027
rect 53297 25993 53331 26027
rect 15117 25925 15151 25959
rect 19717 25925 19751 25959
rect 31539 25925 31573 25959
rect 32689 25925 32723 25959
rect 38209 25925 38243 25959
rect 46121 25925 46155 25959
rect 53021 25925 53055 25959
rect 2053 25857 2087 25891
rect 2145 25857 2179 25891
rect 17417 25857 17451 25891
rect 17693 25857 17727 25891
rect 19625 25857 19659 25891
rect 19901 25857 19935 25891
rect 20361 25857 20395 25891
rect 20913 25857 20947 25891
rect 21281 25857 21315 25891
rect 32597 25857 32631 25891
rect 32781 25857 32815 25891
rect 32965 25857 32999 25891
rect 34529 25857 34563 25891
rect 37473 25857 37507 25891
rect 37657 25857 37691 25891
rect 37749 25857 37783 25891
rect 38025 25857 38059 25891
rect 38301 25857 38335 25891
rect 38393 25857 38427 25891
rect 40785 25857 40819 25891
rect 42625 25857 42659 25891
rect 42717 25857 42751 25891
rect 44557 25857 44591 25891
rect 44649 25857 44683 25891
rect 44833 25857 44867 25891
rect 44925 25857 44959 25891
rect 49341 25857 49375 25891
rect 49525 25857 49559 25891
rect 49617 25857 49651 25891
rect 49709 25857 49743 25891
rect 51273 25857 51307 25891
rect 51365 25857 51399 25891
rect 51641 25857 51675 25891
rect 52745 25857 52779 25891
rect 52929 25857 52963 25891
rect 53113 25857 53147 25891
rect 15485 25789 15519 25823
rect 17509 25789 17543 25823
rect 21189 25789 21223 25823
rect 21649 25789 21683 25823
rect 23305 25789 23339 25823
rect 23581 25789 23615 25823
rect 29745 25789 29779 25823
rect 30113 25789 30147 25823
rect 34253 25789 34287 25823
rect 47409 25789 47443 25823
rect 47685 25789 47719 25823
rect 47869 25789 47903 25823
rect 51549 25789 51583 25823
rect 15393 25721 15427 25755
rect 17233 25721 17267 25755
rect 21833 25721 21867 25755
rect 23765 25721 23799 25755
rect 46489 25721 46523 25755
rect 53389 25721 53423 25755
rect 15255 25653 15289 25687
rect 17693 25653 17727 25687
rect 19901 25653 19935 25687
rect 37289 25653 37323 25687
rect 44373 25653 44407 25687
rect 51825 25653 51859 25687
rect 13277 25449 13311 25483
rect 14289 25449 14323 25483
rect 14565 25449 14599 25483
rect 21005 25449 21039 25483
rect 26985 25449 27019 25483
rect 31033 25449 31067 25483
rect 42073 25449 42107 25483
rect 51917 25449 51951 25483
rect 53665 25449 53699 25483
rect 13461 25381 13495 25415
rect 18705 25381 18739 25415
rect 42349 25381 42383 25415
rect 12817 25313 12851 25347
rect 14197 25313 14231 25347
rect 15577 25313 15611 25347
rect 19257 25313 19291 25347
rect 34437 25313 34471 25347
rect 37841 25313 37875 25347
rect 41061 25313 41095 25347
rect 41153 25313 41187 25347
rect 43269 25313 43303 25347
rect 55321 25313 55355 25347
rect 2053 25245 2087 25279
rect 2145 25245 2179 25279
rect 12909 25245 12943 25279
rect 13277 25245 13311 25279
rect 14381 25245 14415 25279
rect 14657 25245 14691 25279
rect 14841 25245 14875 25279
rect 17601 25245 17635 25279
rect 17693 25245 17727 25279
rect 17969 25245 18003 25279
rect 18061 25245 18095 25279
rect 18889 25245 18923 25279
rect 19073 25245 19107 25279
rect 27077 25245 27111 25279
rect 31217 25245 31251 25279
rect 31401 25245 31435 25279
rect 31585 25245 31619 25279
rect 34161 25245 34195 25279
rect 34253 25245 34287 25279
rect 34529 25245 34563 25279
rect 34897 25245 34931 25279
rect 35081 25245 35115 25279
rect 35265 25245 35299 25279
rect 35725 25245 35759 25279
rect 36093 25245 36127 25279
rect 38209 25245 38243 25279
rect 40969 25245 41003 25279
rect 41429 25245 41463 25279
rect 41521 25245 41555 25279
rect 41889 25245 41923 25279
rect 42441 25245 42475 25279
rect 42993 25245 43027 25279
rect 43637 25245 43671 25279
rect 51641 25245 51675 25279
rect 51733 25245 51767 25279
rect 52009 25245 52043 25279
rect 53113 25245 53147 25279
rect 53389 25245 53423 25279
rect 53481 25245 53515 25279
rect 53711 25245 53745 25279
rect 14105 25177 14139 25211
rect 15853 25177 15887 25211
rect 18429 25177 18463 25211
rect 18981 25177 19015 25211
rect 19533 25177 19567 25211
rect 27813 25177 27847 25211
rect 31309 25177 31343 25211
rect 34989 25177 35023 25211
rect 41337 25177 41371 25211
rect 41705 25177 41739 25211
rect 41797 25177 41831 25211
rect 43453 25177 43487 25211
rect 55597 25177 55631 25211
rect 1869 25109 1903 25143
rect 14749 25109 14783 25143
rect 17325 25109 17359 25143
rect 17417 25109 17451 25143
rect 17785 25109 17819 25143
rect 18153 25109 18187 25143
rect 18337 25109 18371 25143
rect 18521 25109 18555 25143
rect 21097 25109 21131 25143
rect 33977 25109 34011 25143
rect 34713 25109 34747 25143
rect 37519 25109 37553 25143
rect 39635 25109 39669 25143
rect 51457 25109 51491 25143
rect 53205 25109 53239 25143
rect 57069 25109 57103 25143
rect 13185 24905 13219 24939
rect 17601 24905 17635 24939
rect 17785 24905 17819 24939
rect 20069 24905 20103 24939
rect 31033 24905 31067 24939
rect 35219 24905 35253 24939
rect 36461 24905 36495 24939
rect 38209 24905 38243 24939
rect 43453 24905 43487 24939
rect 43545 24905 43579 24939
rect 44081 24905 44115 24939
rect 44741 24905 44775 24939
rect 51365 24905 51399 24939
rect 51917 24905 51951 24939
rect 54769 24905 54803 24939
rect 55689 24905 55723 24939
rect 13001 24837 13035 24871
rect 15469 24837 15503 24871
rect 15669 24837 15703 24871
rect 20269 24837 20303 24871
rect 41889 24837 41923 24871
rect 44281 24837 44315 24871
rect 51089 24837 51123 24871
rect 53297 24837 53331 24871
rect 2053 24769 2087 24803
rect 2145 24769 2179 24803
rect 10333 24769 10367 24803
rect 10793 24769 10827 24803
rect 12357 24769 12391 24803
rect 12541 24769 12575 24803
rect 13093 24769 13127 24803
rect 14197 24769 14231 24803
rect 14289 24769 14323 24803
rect 14473 24769 14507 24803
rect 14565 24769 14599 24803
rect 15209 24769 15243 24803
rect 16957 24769 16991 24803
rect 17693 24769 17727 24803
rect 28457 24769 28491 24803
rect 30573 24769 30607 24803
rect 30665 24769 30699 24803
rect 30941 24769 30975 24803
rect 33793 24769 33827 24803
rect 36645 24769 36679 24803
rect 36737 24769 36771 24803
rect 37013 24769 37047 24803
rect 37565 24769 37599 24803
rect 37749 24769 37783 24803
rect 37841 24769 37875 24803
rect 37933 24769 37967 24803
rect 38393 24769 38427 24803
rect 38485 24769 38519 24803
rect 38761 24769 38795 24803
rect 42073 24769 42107 24803
rect 42717 24769 42751 24803
rect 42809 24769 42843 24803
rect 42901 24769 42935 24803
rect 43085 24769 43119 24803
rect 43637 24769 43671 24803
rect 44649 24769 44683 24803
rect 45017 24769 45051 24803
rect 45201 24769 45235 24803
rect 50813 24769 50847 24803
rect 50997 24769 51031 24803
rect 51181 24769 51215 24803
rect 53021 24769 53055 24803
rect 55137 24769 55171 24803
rect 55413 24769 55447 24803
rect 55505 24769 55539 24803
rect 7757 24701 7791 24735
rect 8033 24701 8067 24735
rect 9505 24701 9539 24735
rect 10149 24701 10183 24735
rect 11069 24701 11103 24735
rect 12817 24701 12851 24735
rect 13461 24701 13495 24735
rect 17141 24701 17175 24735
rect 17233 24701 17267 24735
rect 28825 24701 28859 24735
rect 30389 24701 30423 24735
rect 30849 24701 30883 24735
rect 33425 24701 33459 24735
rect 47685 24701 47719 24735
rect 47961 24701 47995 24735
rect 50077 24701 50111 24735
rect 52561 24701 52595 24735
rect 55045 24701 55079 24735
rect 11345 24633 11379 24667
rect 13369 24633 13403 24667
rect 14473 24633 14507 24667
rect 30251 24633 30285 24667
rect 38117 24633 38151 24667
rect 43821 24633 43855 24667
rect 1869 24565 1903 24599
rect 9597 24565 9631 24599
rect 10885 24565 10919 24599
rect 12541 24565 12575 24599
rect 14105 24565 14139 24599
rect 15301 24565 15335 24599
rect 15485 24565 15519 24599
rect 19901 24565 19935 24599
rect 20085 24565 20119 24599
rect 36921 24565 36955 24599
rect 38669 24565 38703 24599
rect 42441 24565 42475 24599
rect 43269 24565 43303 24599
rect 43913 24565 43947 24599
rect 44097 24565 44131 24599
rect 49433 24565 49467 24599
rect 49525 24565 49559 24599
rect 55229 24565 55263 24599
rect 9045 24361 9079 24395
rect 9873 24361 9907 24395
rect 10793 24361 10827 24395
rect 13369 24361 13403 24395
rect 13829 24361 13863 24395
rect 16221 24361 16255 24395
rect 31125 24361 31159 24395
rect 43913 24361 43947 24395
rect 48421 24361 48455 24395
rect 49801 24361 49835 24395
rect 53389 24361 53423 24395
rect 55873 24361 55907 24395
rect 10149 24293 10183 24327
rect 48329 24293 48363 24327
rect 9413 24225 9447 24259
rect 11897 24225 11931 24259
rect 13553 24225 13587 24259
rect 14749 24225 14783 24259
rect 45477 24225 45511 24259
rect 47501 24225 47535 24259
rect 48881 24225 48915 24259
rect 50813 24225 50847 24259
rect 9321 24157 9355 24191
rect 10701 24157 10735 24191
rect 10793 24157 10827 24191
rect 10885 24157 10919 24191
rect 11621 24157 11655 24191
rect 13461 24157 13495 24191
rect 13645 24157 13679 24191
rect 14473 24157 14507 24191
rect 17417 24157 17451 24191
rect 17601 24157 17635 24191
rect 21097 24157 21131 24191
rect 31309 24157 31343 24191
rect 31493 24157 31527 24191
rect 31677 24157 31711 24191
rect 33333 24157 33367 24191
rect 34345 24157 34379 24191
rect 42717 24157 42751 24191
rect 43821 24157 43855 24191
rect 44005 24157 44039 24191
rect 44281 24157 44315 24191
rect 44465 24157 44499 24191
rect 48605 24157 48639 24191
rect 48697 24157 48731 24191
rect 48973 24157 49007 24191
rect 49249 24157 49283 24191
rect 49433 24157 49467 24191
rect 49617 24157 49651 24191
rect 49985 24157 50019 24191
rect 52837 24157 52871 24191
rect 53113 24157 53147 24191
rect 53205 24157 53239 24191
rect 55321 24157 55355 24191
rect 55689 24157 55723 24191
rect 9857 24089 9891 24123
rect 10057 24089 10091 24123
rect 10425 24089 10459 24123
rect 10517 24089 10551 24123
rect 11069 24089 11103 24123
rect 31401 24089 31435 24123
rect 34069 24089 34103 24123
rect 36093 24089 36127 24123
rect 40049 24089 40083 24123
rect 40233 24089 40267 24123
rect 42533 24089 42567 24123
rect 45753 24089 45787 24123
rect 49341 24089 49375 24123
rect 51089 24089 51123 24123
rect 53021 24089 53055 24123
rect 55505 24089 55539 24123
rect 55597 24089 55631 24123
rect 2053 24021 2087 24055
rect 9689 24021 9723 24055
rect 10333 24021 10367 24055
rect 16313 24021 16347 24055
rect 17509 24021 17543 24055
rect 20453 24021 20487 24055
rect 36277 24021 36311 24055
rect 39865 24021 39899 24055
rect 40417 24021 40451 24055
rect 42349 24021 42383 24055
rect 44097 24021 44131 24055
rect 49065 24021 49099 24055
rect 52561 24021 52595 24055
rect 1869 23817 1903 23851
rect 14105 23817 14139 23851
rect 19073 23817 19107 23851
rect 21557 23817 21591 23851
rect 35909 23817 35943 23851
rect 37105 23817 37139 23851
rect 38209 23817 38243 23851
rect 41061 23817 41095 23851
rect 45937 23817 45971 23851
rect 49801 23817 49835 23851
rect 9045 23749 9079 23783
rect 10609 23749 10643 23783
rect 17233 23749 17267 23783
rect 17601 23749 17635 23783
rect 20085 23749 20119 23783
rect 21833 23749 21867 23783
rect 35081 23749 35115 23783
rect 35541 23749 35575 23783
rect 35633 23749 35667 23783
rect 36369 23749 36403 23783
rect 36461 23749 36495 23783
rect 37565 23749 37599 23783
rect 37657 23749 37691 23783
rect 39589 23749 39623 23783
rect 39926 23749 39960 23783
rect 42441 23749 42475 23783
rect 42993 23749 43027 23783
rect 46305 23749 46339 23783
rect 50905 23749 50939 23783
rect 2053 23681 2087 23715
rect 8769 23681 8803 23715
rect 10793 23681 10827 23715
rect 10977 23681 11011 23715
rect 11069 23681 11103 23715
rect 16957 23681 16991 23715
rect 17049 23681 17083 23715
rect 19349 23681 19383 23715
rect 30113 23681 30147 23715
rect 31907 23681 31941 23715
rect 34575 23681 34609 23715
rect 34897 23681 34931 23715
rect 34989 23681 35023 23715
rect 35265 23681 35299 23715
rect 35357 23681 35391 23715
rect 35725 23681 35759 23715
rect 36093 23681 36127 23715
rect 36186 23681 36220 23715
rect 36558 23681 36592 23715
rect 37473 23681 37507 23715
rect 37841 23681 37875 23715
rect 38945 23681 38979 23715
rect 39129 23681 39163 23715
rect 39221 23681 39255 23715
rect 39313 23681 39347 23715
rect 42901 23681 42935 23715
rect 43177 23681 43211 23715
rect 44281 23681 44315 23715
rect 44373 23681 44407 23715
rect 44465 23681 44499 23715
rect 46397 23681 46431 23715
rect 47961 23681 47995 23715
rect 48237 23681 48271 23715
rect 48329 23681 48363 23715
rect 48605 23681 48639 23715
rect 48881 23681 48915 23715
rect 49617 23681 49651 23715
rect 49985 23681 50019 23715
rect 50629 23681 50663 23715
rect 50813 23681 50847 23715
rect 51021 23681 51055 23715
rect 54309 23681 54343 23715
rect 54493 23681 54527 23715
rect 54585 23681 54619 23715
rect 54677 23681 54711 23715
rect 77861 23681 77895 23715
rect 78045 23681 78079 23715
rect 2145 23613 2179 23647
rect 10517 23613 10551 23647
rect 14657 23613 14691 23647
rect 17325 23613 17359 23647
rect 19441 23613 19475 23647
rect 19717 23613 19751 23647
rect 19809 23613 19843 23647
rect 30481 23613 30515 23647
rect 32781 23613 32815 23647
rect 33149 23613 33183 23647
rect 39681 23613 39715 23647
rect 44557 23613 44591 23647
rect 45845 23613 45879 23647
rect 46581 23613 46615 23647
rect 48513 23613 48547 23647
rect 49433 23613 49467 23647
rect 50261 23613 50295 23647
rect 17233 23545 17267 23579
rect 32229 23545 32263 23579
rect 36829 23545 36863 23579
rect 38025 23545 38059 23579
rect 43269 23545 43303 23579
rect 50537 23545 50571 23579
rect 34713 23477 34747 23511
rect 36737 23477 36771 23511
rect 37289 23477 37323 23511
rect 44741 23477 44775 23511
rect 48053 23477 48087 23511
rect 51181 23477 51215 23511
rect 54861 23477 54895 23511
rect 78229 23477 78263 23511
rect 17417 23273 17451 23307
rect 17601 23273 17635 23307
rect 18705 23273 18739 23307
rect 29929 23273 29963 23307
rect 30757 23273 30791 23307
rect 31217 23273 31251 23307
rect 33333 23273 33367 23307
rect 40509 23273 40543 23307
rect 42165 23273 42199 23307
rect 49157 23273 49191 23307
rect 53389 23273 53423 23307
rect 53757 23273 53791 23307
rect 55321 23273 55355 23307
rect 58541 23273 58575 23307
rect 2329 23205 2363 23239
rect 35817 23205 35851 23239
rect 2513 23137 2547 23171
rect 10885 23137 10919 23171
rect 11161 23137 11195 23171
rect 17969 23137 18003 23171
rect 33793 23137 33827 23171
rect 41429 23137 41463 23171
rect 43085 23137 43119 23171
rect 44189 23137 44223 23171
rect 44281 23137 44315 23171
rect 44473 23137 44507 23171
rect 45201 23137 45235 23171
rect 45293 23137 45327 23171
rect 45477 23137 45511 23171
rect 47593 23137 47627 23171
rect 49525 23137 49559 23171
rect 2053 23069 2087 23103
rect 2145 23069 2179 23103
rect 10793 23069 10827 23103
rect 14657 23069 14691 23103
rect 16405 23069 16439 23103
rect 29653 23069 29687 23103
rect 29745 23069 29779 23103
rect 30113 23069 30147 23103
rect 30481 23069 30515 23103
rect 30941 23069 30975 23103
rect 31033 23069 31067 23103
rect 31309 23069 31343 23103
rect 33517 23069 33551 23103
rect 33609 23069 33643 23103
rect 33885 23069 33919 23103
rect 35265 23069 35299 23103
rect 35449 23069 35483 23103
rect 35633 23069 35667 23103
rect 36277 23069 36311 23103
rect 36369 23069 36403 23103
rect 36553 23069 36587 23103
rect 36645 23069 36679 23103
rect 36921 23069 36955 23103
rect 39865 23069 39899 23103
rect 39958 23069 39992 23103
rect 40330 23069 40364 23103
rect 41889 23069 41923 23103
rect 42257 23069 42291 23103
rect 43729 23069 43763 23103
rect 43821 23069 43855 23103
rect 43913 23069 43947 23103
rect 44373 23069 44407 23103
rect 45385 23069 45419 23103
rect 46121 23069 46155 23103
rect 46397 23069 46431 23103
rect 47317 23069 47351 23103
rect 49341 23069 49375 23103
rect 51089 23069 51123 23103
rect 51237 23069 51271 23103
rect 51554 23069 51588 23103
rect 53113 23069 53147 23103
rect 53205 23069 53239 23103
rect 53481 23069 53515 23103
rect 54033 23069 54067 23103
rect 54585 23069 54619 23103
rect 57069 23069 57103 23103
rect 57161 23069 57195 23103
rect 17141 23001 17175 23035
rect 17785 23001 17819 23035
rect 18245 23001 18279 23035
rect 18521 23001 18555 23035
rect 30297 23001 30331 23035
rect 30389 23001 30423 23035
rect 35541 23001 35575 23035
rect 36001 23001 36035 23035
rect 40141 23001 40175 23035
rect 40233 23001 40267 23035
rect 41981 23001 42015 23035
rect 43269 23001 43303 23035
rect 46489 23001 46523 23035
rect 50905 23001 50939 23035
rect 51365 23001 51399 23035
rect 51457 23001 51491 23035
rect 53665 23001 53699 23035
rect 56793 23001 56827 23035
rect 57406 23001 57440 23035
rect 1869 22933 1903 22967
rect 14105 22933 14139 22967
rect 17575 22933 17609 22967
rect 19349 22933 19383 22967
rect 30665 22933 30699 22967
rect 36185 22933 36219 22967
rect 36829 22933 36863 22967
rect 40601 22933 40635 22967
rect 44649 22933 44683 22967
rect 45017 22933 45051 22967
rect 49065 22933 49099 22967
rect 49709 22933 49743 22967
rect 50721 22933 50755 22967
rect 51733 22933 51767 22967
rect 52929 22933 52963 22967
rect 10701 22729 10735 22763
rect 13645 22729 13679 22763
rect 18521 22729 18555 22763
rect 19441 22729 19475 22763
rect 30665 22729 30699 22763
rect 32781 22729 32815 22763
rect 38301 22729 38335 22763
rect 38485 22729 38519 22763
rect 39129 22729 39163 22763
rect 39957 22729 39991 22763
rect 43361 22729 43395 22763
rect 49065 22729 49099 22763
rect 51181 22729 51215 22763
rect 51733 22729 51767 22763
rect 56885 22729 56919 22763
rect 58633 22729 58667 22763
rect 9689 22661 9723 22695
rect 10517 22661 10551 22695
rect 11621 22661 11655 22695
rect 15485 22661 15519 22695
rect 19349 22661 19383 22695
rect 19809 22661 19843 22695
rect 33149 22661 33183 22695
rect 35173 22661 35207 22695
rect 35817 22661 35851 22695
rect 37749 22661 37783 22695
rect 37841 22661 37875 22695
rect 39221 22661 39255 22695
rect 50813 22661 50847 22695
rect 50905 22661 50939 22695
rect 51273 22661 51307 22695
rect 53021 22661 53055 22695
rect 55413 22661 55447 22695
rect 56057 22661 56091 22695
rect 13093 22593 13127 22627
rect 27997 22593 28031 22627
rect 30113 22593 30147 22627
rect 30205 22593 30239 22627
rect 30297 22593 30331 22627
rect 30481 22593 30515 22627
rect 32321 22593 32355 22627
rect 32413 22593 32447 22627
rect 32689 22593 32723 22627
rect 32965 22593 32999 22627
rect 33057 22593 33091 22627
rect 33313 22593 33347 22627
rect 34897 22593 34931 22627
rect 35081 22593 35115 22627
rect 35265 22593 35299 22627
rect 36553 22593 36587 22627
rect 37565 22593 37599 22627
rect 37933 22593 37967 22627
rect 38393 22593 38427 22627
rect 39313 22593 39347 22627
rect 39589 22593 39623 22627
rect 39681 22593 39715 22627
rect 42441 22593 42475 22627
rect 42625 22593 42659 22627
rect 42717 22593 42751 22627
rect 43637 22593 43671 22627
rect 43821 22593 43855 22627
rect 48237 22593 48271 22627
rect 48421 22593 48455 22627
rect 48569 22593 48603 22627
rect 48697 22593 48731 22627
rect 48789 22593 48823 22627
rect 48886 22593 48920 22627
rect 49617 22593 49651 22627
rect 49709 22593 49743 22627
rect 49802 22593 49836 22627
rect 49985 22593 50019 22627
rect 50077 22593 50111 22627
rect 50174 22593 50208 22627
rect 50537 22593 50571 22627
rect 50685 22593 50719 22627
rect 51002 22593 51036 22627
rect 51549 22593 51583 22627
rect 54861 22593 54895 22627
rect 55137 22593 55171 22627
rect 55229 22593 55263 22627
rect 56241 22593 56275 22627
rect 56425 22593 56459 22627
rect 56517 22593 56551 22627
rect 56609 22593 56643 22627
rect 57897 22593 57931 22627
rect 58541 22593 58575 22627
rect 11253 22525 11287 22559
rect 13001 22525 13035 22559
rect 15117 22525 15151 22559
rect 15393 22525 15427 22559
rect 16681 22525 16715 22559
rect 16957 22525 16991 22559
rect 18429 22525 18463 22559
rect 19073 22525 19107 22559
rect 28365 22525 28399 22559
rect 36645 22525 36679 22559
rect 43177 22525 43211 22559
rect 43545 22525 43579 22559
rect 43729 22525 43763 22559
rect 51365 22525 51399 22559
rect 52745 22525 52779 22559
rect 13461 22457 13495 22491
rect 29791 22457 29825 22491
rect 35449 22457 35483 22491
rect 36921 22457 36955 22491
rect 38117 22457 38151 22491
rect 38761 22457 38795 22491
rect 38853 22457 38887 22491
rect 39865 22457 39899 22491
rect 50353 22457 50387 22491
rect 54677 22457 54711 22491
rect 29929 22389 29963 22423
rect 32137 22389 32171 22423
rect 32597 22389 32631 22423
rect 35633 22389 35667 22423
rect 36737 22389 36771 22423
rect 38669 22389 38703 22423
rect 40233 22389 40267 22423
rect 48053 22389 48087 22423
rect 49157 22389 49191 22423
rect 49433 22389 49467 22423
rect 51273 22389 51307 22423
rect 54493 22389 54527 22423
rect 54953 22389 54987 22423
rect 11725 22185 11759 22219
rect 14933 22185 14967 22219
rect 16589 22185 16623 22219
rect 29193 22185 29227 22219
rect 30021 22185 30055 22219
rect 45017 22185 45051 22219
rect 45845 22185 45879 22219
rect 49801 22185 49835 22219
rect 53297 22185 53331 22219
rect 13001 22117 13035 22151
rect 30481 22117 30515 22151
rect 31033 22117 31067 22151
rect 46673 22117 46707 22151
rect 11989 22049 12023 22083
rect 12725 22049 12759 22083
rect 14289 22049 14323 22083
rect 17049 22049 17083 22083
rect 18613 22049 18647 22083
rect 29561 22049 29595 22083
rect 32413 22049 32447 22083
rect 33839 22049 33873 22083
rect 46581 22049 46615 22083
rect 47409 22049 47443 22083
rect 49157 22049 49191 22083
rect 50353 22049 50387 22083
rect 54125 22049 54159 22083
rect 1685 21981 1719 22015
rect 16957 21981 16991 22015
rect 29377 21981 29411 22015
rect 29745 21981 29779 22015
rect 29837 21981 29871 22015
rect 30113 21981 30147 22015
rect 30297 21981 30331 22015
rect 31125 21981 31159 22015
rect 31401 21981 31435 22015
rect 32045 21981 32079 22015
rect 42625 21981 42659 22015
rect 45201 21981 45235 22015
rect 45293 21981 45327 22015
rect 46029 21981 46063 22015
rect 46121 21981 46155 22015
rect 46949 21981 46983 22015
rect 49249 21981 49283 22015
rect 49617 21981 49651 22015
rect 52745 21981 52779 22015
rect 53021 21981 53055 22015
rect 53113 21981 53147 22015
rect 30849 21913 30883 21947
rect 37197 21913 37231 21947
rect 37565 21913 37599 21947
rect 37841 21913 37875 21947
rect 41797 21913 41831 21947
rect 42165 21913 42199 21947
rect 42257 21913 42291 21947
rect 42533 21913 42567 21947
rect 42993 21913 43027 21947
rect 43085 21913 43119 21947
rect 43361 21913 43395 21947
rect 45753 21913 45787 21947
rect 46857 21913 46891 21947
rect 48973 21913 49007 21947
rect 49433 21913 49467 21947
rect 49525 21913 49559 21947
rect 52929 21913 52963 21947
rect 53389 21913 53423 21947
rect 1501 21845 1535 21879
rect 10241 21845 10275 21879
rect 13185 21845 13219 21879
rect 38301 21845 38335 21879
rect 39313 21845 39347 21879
rect 42349 21845 42383 21879
rect 43177 21845 43211 21879
rect 50169 21845 50203 21879
rect 12449 21641 12483 21675
rect 31217 21641 31251 21675
rect 51273 21641 51307 21675
rect 53297 21641 53331 21675
rect 13921 21573 13955 21607
rect 30021 21573 30055 21607
rect 30113 21573 30147 21607
rect 37565 21573 37599 21607
rect 45201 21573 45235 21607
rect 45937 21573 45971 21607
rect 50261 21573 50295 21607
rect 54769 21573 54803 21607
rect 1685 21505 1719 21539
rect 7573 21505 7607 21539
rect 29745 21505 29779 21539
rect 29837 21505 29871 21539
rect 30205 21505 30239 21539
rect 30665 21505 30699 21539
rect 30757 21505 30791 21539
rect 31033 21505 31067 21539
rect 31401 21505 31435 21539
rect 33885 21505 33919 21539
rect 37473 21505 37507 21539
rect 37657 21505 37691 21539
rect 37841 21505 37875 21539
rect 40049 21505 40083 21539
rect 45109 21505 45143 21539
rect 45293 21505 45327 21539
rect 45753 21505 45787 21539
rect 46029 21505 46063 21539
rect 47777 21505 47811 21539
rect 47869 21505 47903 21539
rect 49985 21505 50019 21539
rect 50169 21505 50203 21539
rect 50353 21505 50387 21539
rect 50629 21505 50663 21539
rect 50722 21505 50756 21539
rect 50905 21505 50939 21539
rect 50997 21505 51031 21539
rect 51135 21505 51169 21539
rect 54585 21505 54619 21539
rect 54861 21505 54895 21539
rect 54953 21505 54987 21539
rect 56977 21505 57011 21539
rect 7849 21437 7883 21471
rect 14197 21437 14231 21471
rect 30481 21437 30515 21471
rect 34161 21437 34195 21471
rect 35633 21437 35667 21471
rect 36369 21437 36403 21471
rect 39773 21437 39807 21471
rect 44649 21437 44683 21471
rect 56701 21437 56735 21471
rect 29561 21369 29595 21403
rect 30941 21369 30975 21403
rect 35725 21369 35759 21403
rect 49709 21369 49743 21403
rect 50537 21369 50571 21403
rect 1501 21301 1535 21335
rect 9321 21301 9355 21335
rect 30389 21301 30423 21335
rect 31493 21301 31527 21335
rect 37289 21301 37323 21335
rect 38301 21301 38335 21335
rect 46213 21301 46247 21335
rect 47593 21301 47627 21335
rect 48053 21301 48087 21335
rect 49801 21301 49835 21335
rect 55137 21301 55171 21335
rect 55229 21301 55263 21335
rect 7573 21097 7607 21131
rect 14749 21097 14783 21131
rect 39681 21097 39715 21131
rect 50537 21097 50571 21131
rect 51089 21097 51123 21131
rect 53205 21097 53239 21131
rect 56149 21097 56183 21131
rect 56609 21097 56643 21131
rect 50353 21029 50387 21063
rect 7021 20961 7055 20995
rect 8125 20961 8159 20995
rect 9781 20961 9815 20995
rect 29929 20961 29963 20995
rect 37749 20961 37783 20995
rect 39221 20961 39255 20995
rect 39865 20961 39899 20995
rect 52285 20961 52319 20995
rect 54217 20961 54251 20995
rect 55321 20961 55355 20995
rect 1685 20893 1719 20927
rect 7113 20893 7147 20927
rect 7297 20893 7331 20927
rect 8401 20893 8435 20927
rect 11345 20893 11379 20927
rect 11529 20893 11563 20927
rect 14473 20893 14507 20927
rect 29561 20893 29595 20927
rect 34897 20893 34931 20927
rect 35265 20893 35299 20927
rect 38485 20893 38519 20927
rect 39037 20893 39071 20927
rect 39129 20893 39163 20927
rect 39405 20893 39439 20927
rect 39497 20893 39531 20927
rect 42625 20893 42659 20927
rect 44373 20893 44407 20927
rect 45017 20893 45051 20927
rect 48973 20893 49007 20927
rect 49065 20893 49099 20927
rect 49157 20893 49191 20927
rect 49341 20893 49375 20927
rect 50813 20893 50847 20927
rect 50905 20893 50939 20927
rect 51181 20893 51215 20927
rect 51733 20893 51767 20927
rect 52929 20893 52963 20927
rect 53021 20893 53055 20927
rect 53297 20893 53331 20927
rect 53665 20893 53699 20927
rect 54401 20893 54435 20927
rect 54677 20893 54711 20927
rect 54769 20893 54803 20927
rect 55965 20893 55999 20927
rect 56057 20893 56091 20927
rect 56333 20893 56367 20927
rect 56425 20893 56459 20927
rect 8033 20825 8067 20859
rect 8585 20825 8619 20859
rect 8769 20825 8803 20859
rect 31493 20825 31527 20859
rect 35081 20825 35115 20859
rect 35173 20825 35207 20859
rect 37473 20825 37507 20859
rect 40141 20825 40175 20859
rect 42165 20825 42199 20859
rect 42533 20825 42567 20859
rect 42901 20825 42935 20859
rect 44097 20825 44131 20859
rect 44465 20825 44499 20859
rect 44833 20825 44867 20859
rect 54585 20825 54619 20859
rect 1501 20757 1535 20791
rect 7481 20757 7515 20791
rect 7941 20757 7975 20791
rect 10425 20757 10459 20791
rect 11437 20757 11471 20791
rect 14197 20757 14231 20791
rect 31355 20757 31389 20791
rect 35449 20757 35483 20791
rect 36001 20757 36035 20791
rect 41613 20757 41647 20791
rect 42717 20757 42751 20791
rect 44281 20757 44315 20791
rect 45201 20757 45235 20791
rect 48605 20757 48639 20791
rect 48789 20757 48823 20791
rect 50629 20757 50663 20791
rect 52745 20757 52779 20791
rect 54953 20757 54987 20791
rect 56701 20757 56735 20791
rect 7573 20553 7607 20587
rect 34713 20553 34747 20587
rect 38577 20553 38611 20587
rect 39681 20553 39715 20587
rect 41521 20553 41555 20587
rect 43913 20553 43947 20587
rect 55965 20553 55999 20587
rect 8125 20485 8159 20519
rect 12541 20485 12575 20519
rect 38209 20485 38243 20519
rect 43453 20485 43487 20519
rect 47225 20485 47259 20519
rect 50813 20485 50847 20519
rect 53021 20485 53055 20519
rect 56517 20485 56551 20519
rect 7573 20417 7607 20451
rect 7757 20417 7791 20451
rect 7849 20417 7883 20451
rect 9781 20417 9815 20451
rect 9965 20417 9999 20451
rect 10425 20417 10459 20451
rect 23581 20417 23615 20451
rect 27905 20417 27939 20451
rect 32137 20417 32171 20451
rect 34897 20417 34931 20451
rect 34989 20417 35023 20451
rect 35265 20417 35299 20451
rect 36645 20417 36679 20451
rect 36737 20417 36771 20451
rect 37013 20417 37047 20451
rect 37289 20417 37323 20451
rect 38025 20417 38059 20451
rect 38301 20417 38335 20451
rect 38393 20417 38427 20451
rect 39865 20417 39899 20451
rect 39957 20417 39991 20451
rect 40233 20417 40267 20451
rect 40693 20417 40727 20451
rect 41613 20417 41647 20451
rect 46673 20417 46707 20451
rect 46765 20417 46799 20451
rect 48145 20417 48179 20451
rect 50537 20417 50571 20451
rect 52745 20417 52779 20451
rect 54861 20417 54895 20451
rect 55137 20417 55171 20451
rect 55229 20417 55263 20451
rect 55781 20417 55815 20451
rect 56793 20417 56827 20451
rect 9597 20349 9631 20383
rect 10149 20349 10183 20383
rect 10241 20349 10275 20383
rect 12265 20349 12299 20383
rect 14013 20349 14047 20383
rect 14289 20349 14323 20383
rect 28641 20349 28675 20383
rect 32413 20349 32447 20383
rect 33885 20349 33919 20383
rect 34621 20349 34655 20383
rect 36461 20349 36495 20383
rect 37841 20349 37875 20383
rect 41245 20349 41279 20383
rect 46489 20349 46523 20383
rect 48421 20349 48455 20383
rect 52285 20349 52319 20383
rect 23765 20281 23799 20315
rect 43821 20281 43855 20315
rect 54493 20281 54527 20315
rect 55597 20281 55631 20315
rect 9873 20213 9907 20247
rect 10609 20213 10643 20247
rect 14933 20213 14967 20247
rect 22293 20213 22327 20247
rect 27721 20213 27755 20247
rect 33977 20213 34011 20247
rect 35173 20213 35207 20247
rect 36921 20213 36955 20247
rect 39497 20213 39531 20247
rect 40141 20213 40175 20247
rect 41889 20213 41923 20247
rect 49893 20213 49927 20247
rect 54953 20213 54987 20247
rect 55413 20213 55447 20247
rect 56241 20213 56275 20247
rect 56885 20213 56919 20247
rect 7573 20009 7607 20043
rect 7757 20009 7791 20043
rect 9873 20009 9907 20043
rect 10057 20009 10091 20043
rect 11897 20009 11931 20043
rect 28411 20009 28445 20043
rect 31769 20009 31803 20043
rect 33333 20009 33367 20043
rect 34069 20009 34103 20043
rect 36645 20009 36679 20043
rect 46489 20009 46523 20043
rect 47501 20009 47535 20043
rect 48605 20009 48639 20043
rect 49065 20009 49099 20043
rect 50905 20009 50939 20043
rect 51181 20009 51215 20043
rect 52837 20009 52871 20043
rect 55321 20009 55355 20043
rect 45477 19941 45511 19975
rect 48513 19941 48547 19975
rect 10149 19873 10183 19907
rect 12173 19873 12207 19907
rect 12817 19873 12851 19907
rect 14289 19873 14323 19907
rect 14565 19873 14599 19907
rect 33793 19873 33827 19907
rect 45661 19873 45695 19907
rect 56793 19873 56827 19907
rect 57069 19873 57103 19907
rect 1685 19805 1719 19839
rect 7113 19805 7147 19839
rect 7205 19805 7239 19839
rect 7297 19805 7331 19839
rect 9413 19805 9447 19839
rect 9505 19805 9539 19839
rect 9873 19805 9907 19839
rect 12909 19805 12943 19839
rect 13093 19805 13127 19839
rect 18521 19805 18555 19839
rect 26617 19805 26651 19839
rect 26985 19805 27019 19839
rect 33241 19805 33275 19839
rect 33517 19805 33551 19839
rect 33609 19805 33643 19839
rect 33885 19805 33919 19839
rect 34897 19805 34931 19839
rect 34989 19805 35023 19839
rect 35265 19805 35299 19839
rect 42073 19805 42107 19839
rect 42257 19805 42291 19839
rect 46673 19805 46707 19839
rect 46765 19805 46799 19839
rect 48789 19805 48823 19839
rect 48881 19805 48915 19839
rect 49157 19805 49191 19839
rect 49249 19805 49283 19839
rect 50169 19805 50203 19839
rect 50353 19805 50387 19839
rect 50537 19805 50571 19839
rect 50721 19805 50755 19839
rect 50997 19805 51031 19839
rect 51365 19805 51399 19839
rect 52285 19805 52319 19839
rect 52561 19805 52595 19839
rect 52653 19805 52687 19839
rect 7941 19737 7975 19771
rect 10425 19737 10459 19771
rect 28549 19737 28583 19771
rect 35081 19737 35115 19771
rect 42441 19737 42475 19771
rect 45201 19737 45235 19771
rect 47225 19737 47259 19771
rect 47317 19737 47351 19771
rect 50629 19737 50663 19771
rect 52469 19737 52503 19771
rect 1501 19669 1535 19703
rect 7481 19669 7515 19703
rect 7741 19669 7775 19703
rect 13001 19669 13035 19703
rect 16037 19669 16071 19703
rect 17969 19669 18003 19703
rect 34713 19669 34747 19703
rect 36829 19669 36863 19703
rect 41889 19669 41923 19703
rect 42165 19669 42199 19703
rect 47517 19669 47551 19703
rect 47685 19669 47719 19703
rect 12081 19465 12115 19499
rect 14473 19465 14507 19499
rect 37105 19465 37139 19499
rect 38393 19465 38427 19499
rect 40049 19465 40083 19499
rect 41429 19465 41463 19499
rect 43269 19465 43303 19499
rect 43545 19465 43579 19499
rect 44281 19465 44315 19499
rect 44465 19465 44499 19499
rect 47317 19465 47351 19499
rect 47593 19465 47627 19499
rect 13001 19397 13035 19431
rect 17868 19397 17902 19431
rect 37933 19397 37967 19431
rect 40509 19397 40543 19431
rect 41613 19397 41647 19431
rect 47869 19397 47903 19431
rect 47961 19397 47995 19431
rect 7573 19329 7607 19363
rect 7757 19329 7791 19363
rect 7849 19329 7883 19363
rect 10609 19329 10643 19363
rect 10793 19329 10827 19363
rect 12173 19329 12207 19363
rect 12725 19329 12759 19363
rect 17601 19329 17635 19363
rect 24593 19329 24627 19363
rect 27169 19329 27203 19363
rect 27261 19329 27295 19363
rect 27353 19329 27387 19363
rect 27537 19329 27571 19363
rect 28089 19329 28123 19363
rect 30205 19329 30239 19363
rect 32781 19329 32815 19363
rect 33057 19329 33091 19363
rect 35909 19329 35943 19363
rect 36093 19329 36127 19363
rect 36185 19329 36219 19363
rect 36277 19329 36311 19363
rect 36553 19329 36587 19363
rect 36737 19329 36771 19363
rect 36829 19329 36863 19363
rect 36921 19329 36955 19363
rect 37565 19329 37599 19363
rect 37713 19329 37747 19363
rect 37841 19329 37875 19363
rect 38030 19329 38064 19363
rect 39497 19329 39531 19363
rect 39681 19329 39715 19363
rect 39773 19329 39807 19363
rect 39865 19329 39899 19363
rect 40325 19329 40359 19363
rect 40417 19329 40451 19363
rect 40693 19329 40727 19363
rect 40877 19329 40911 19363
rect 41061 19329 41095 19363
rect 41153 19329 41187 19363
rect 41269 19329 41303 19363
rect 43085 19329 43119 19363
rect 43729 19329 43763 19363
rect 44189 19329 44223 19363
rect 44557 19329 44591 19363
rect 47777 19329 47811 19363
rect 48079 19329 48113 19363
rect 50997 19329 51031 19363
rect 9873 19261 9907 19295
rect 19625 19261 19659 19295
rect 24869 19261 24903 19295
rect 28365 19261 28399 19295
rect 29837 19261 29871 19295
rect 30481 19261 30515 19295
rect 31953 19261 31987 19295
rect 33241 19261 33275 19295
rect 37381 19261 37415 19295
rect 38485 19261 38519 19295
rect 43821 19261 43855 19295
rect 44649 19261 44683 19295
rect 48237 19261 48271 19295
rect 18981 19193 19015 19227
rect 26985 19193 27019 19227
rect 7389 19125 7423 19159
rect 10517 19125 10551 19159
rect 10793 19125 10827 19159
rect 19073 19125 19107 19159
rect 26341 19125 26375 19159
rect 32137 19125 32171 19159
rect 32873 19125 32907 19159
rect 36461 19125 36495 19159
rect 38209 19125 38243 19159
rect 40141 19125 40175 19159
rect 42441 19125 42475 19159
rect 42993 19125 43027 19159
rect 44833 19125 44867 19159
rect 51181 19125 51215 19159
rect 8769 18921 8803 18955
rect 15926 18921 15960 18955
rect 18061 18921 18095 18955
rect 28365 18921 28399 18955
rect 29837 18921 29871 18955
rect 31125 18921 31159 18955
rect 31585 18921 31619 18955
rect 37289 18921 37323 18955
rect 38209 18921 38243 18955
rect 38577 18921 38611 18955
rect 40141 18921 40175 18955
rect 40417 18921 40451 18955
rect 41061 18921 41095 18955
rect 52009 18921 52043 18955
rect 19533 18853 19567 18887
rect 36829 18853 36863 18887
rect 38025 18853 38059 18887
rect 38669 18853 38703 18887
rect 39865 18853 39899 18887
rect 48605 18853 48639 18887
rect 52193 18853 52227 18887
rect 54493 18853 54527 18887
rect 7021 18785 7055 18819
rect 15669 18785 15703 18819
rect 18521 18785 18555 18819
rect 18613 18785 18647 18819
rect 19257 18785 19291 18819
rect 29009 18785 29043 18819
rect 34345 18785 34379 18819
rect 38209 18785 38243 18819
rect 40141 18785 40175 18819
rect 50261 18785 50295 18819
rect 54309 18785 54343 18819
rect 9413 18717 9447 18751
rect 10057 18717 10091 18751
rect 10241 18717 10275 18751
rect 18429 18717 18463 18751
rect 23305 18717 23339 18751
rect 28490 18717 28524 18751
rect 28917 18717 28951 18751
rect 29561 18717 29595 18751
rect 31309 18717 31343 18751
rect 31401 18717 31435 18751
rect 31677 18717 31711 18751
rect 32137 18717 32171 18751
rect 32413 18717 32447 18751
rect 32505 18717 32539 18751
rect 33241 18717 33275 18751
rect 33425 18717 33459 18751
rect 33517 18717 33551 18751
rect 33633 18717 33667 18751
rect 34069 18717 34103 18751
rect 34161 18717 34195 18751
rect 34437 18717 34471 18751
rect 34897 18717 34931 18751
rect 35449 18717 35483 18751
rect 36185 18717 36219 18751
rect 36278 18717 36312 18751
rect 36461 18717 36495 18751
rect 36553 18717 36587 18751
rect 36691 18717 36725 18751
rect 37381 18717 37415 18751
rect 37474 18717 37508 18751
rect 37657 18717 37691 18751
rect 37846 18717 37880 18751
rect 38117 18717 38151 18751
rect 38393 18717 38427 18751
rect 38853 18717 38887 18751
rect 39001 18717 39035 18751
rect 39129 18717 39163 18751
rect 39359 18717 39393 18751
rect 39589 18717 39623 18751
rect 40233 18717 40267 18751
rect 41245 18717 41279 18751
rect 43545 18717 43579 18751
rect 43821 18717 43855 18751
rect 48421 18717 48455 18751
rect 48697 18717 48731 18751
rect 49341 18717 49375 18751
rect 49985 18717 50019 18751
rect 54401 18717 54435 18751
rect 54677 18717 54711 18751
rect 7297 18649 7331 18683
rect 28273 18649 28307 18683
rect 29193 18649 29227 18683
rect 32321 18649 32355 18683
rect 37013 18649 37047 18683
rect 37749 18649 37783 18683
rect 39221 18649 39255 18683
rect 40877 18649 40911 18683
rect 43269 18649 43303 18683
rect 50537 18649 50571 18683
rect 54033 18649 54067 18683
rect 9965 18581 9999 18615
rect 10149 18581 10183 18615
rect 17417 18581 17451 18615
rect 19717 18581 19751 18615
rect 22661 18581 22695 18615
rect 28549 18581 28583 18615
rect 29285 18581 29319 18615
rect 29653 18581 29687 18615
rect 32689 18581 32723 18615
rect 33793 18581 33827 18615
rect 33885 18581 33919 18615
rect 39497 18581 39531 18615
rect 42533 18581 42567 18615
rect 43177 18581 43211 18615
rect 48237 18581 48271 18615
rect 52561 18581 52595 18615
rect 54861 18581 54895 18615
rect 20453 18377 20487 18411
rect 21649 18377 21683 18411
rect 23857 18377 23891 18411
rect 25053 18377 25087 18411
rect 25789 18377 25823 18411
rect 26065 18377 26099 18411
rect 28365 18377 28399 18411
rect 28917 18377 28951 18411
rect 36277 18377 36311 18411
rect 36553 18377 36587 18411
rect 36829 18377 36863 18411
rect 37473 18377 37507 18411
rect 40509 18377 40543 18411
rect 42625 18377 42659 18411
rect 49801 18377 49835 18411
rect 50997 18377 51031 18411
rect 54217 18377 54251 18411
rect 56609 18377 56643 18411
rect 22385 18309 22419 18343
rect 28457 18309 28491 18343
rect 29285 18309 29319 18343
rect 33885 18309 33919 18343
rect 36001 18309 36035 18343
rect 37657 18309 37691 18343
rect 38117 18309 38151 18343
rect 48329 18309 48363 18343
rect 50629 18309 50663 18343
rect 56149 18309 56183 18343
rect 9689 18241 9723 18275
rect 9873 18241 9907 18275
rect 18827 18241 18861 18275
rect 18981 18241 19015 18275
rect 20085 18241 20119 18275
rect 20269 18241 20303 18275
rect 20637 18241 20671 18275
rect 21281 18241 21315 18275
rect 24317 18241 24351 18275
rect 24501 18241 24535 18275
rect 25237 18241 25271 18275
rect 25513 18241 25547 18275
rect 25697 18241 25731 18275
rect 25973 18241 26007 18275
rect 26433 18241 26467 18275
rect 28089 18241 28123 18275
rect 28181 18241 28215 18275
rect 28273 18241 28307 18275
rect 28549 18241 28583 18275
rect 28641 18241 28675 18275
rect 29101 18241 29135 18275
rect 30665 18241 30699 18275
rect 32321 18241 32355 18275
rect 32413 18241 32447 18275
rect 32689 18241 32723 18275
rect 35725 18241 35759 18275
rect 35909 18241 35943 18275
rect 36093 18241 36127 18275
rect 36645 18241 36679 18275
rect 37289 18241 37323 18275
rect 42441 18241 42475 18275
rect 45293 18241 45327 18275
rect 48053 18241 48087 18275
rect 50261 18241 50295 18275
rect 50354 18241 50388 18275
rect 50537 18241 50571 18275
rect 50767 18241 50801 18275
rect 51181 18241 51215 18275
rect 52469 18241 52503 18275
rect 53021 18241 53055 18275
rect 54033 18241 54067 18275
rect 56425 18241 56459 18275
rect 14289 18173 14323 18207
rect 21373 18173 21407 18207
rect 22109 18173 22143 18207
rect 24409 18173 24443 18207
rect 26249 18173 26283 18207
rect 26341 18173 26375 18207
rect 26525 18173 26559 18207
rect 29469 18173 29503 18207
rect 33609 18173 33643 18207
rect 39773 18173 39807 18207
rect 41981 18173 42015 18207
rect 42257 18173 42291 18207
rect 42809 18173 42843 18207
rect 43085 18173 43119 18207
rect 45569 18173 45603 18207
rect 51457 18173 51491 18207
rect 51825 18173 51859 18207
rect 53665 18173 53699 18207
rect 53757 18173 53791 18207
rect 53849 18173 53883 18207
rect 18613 18105 18647 18139
rect 25329 18105 25363 18139
rect 25421 18105 25455 18139
rect 25973 18105 26007 18139
rect 35633 18105 35667 18139
rect 37105 18105 37139 18139
rect 50905 18105 50939 18139
rect 9689 18037 9723 18071
rect 13645 18037 13679 18071
rect 20177 18037 20211 18071
rect 27905 18037 27939 18071
rect 30481 18037 30515 18071
rect 30757 18037 30791 18071
rect 32137 18037 32171 18071
rect 32597 18037 32631 18071
rect 35357 18037 35391 18071
rect 37841 18037 37875 18071
rect 39221 18037 39255 18071
rect 44557 18037 44591 18071
rect 47041 18037 47075 18071
rect 51365 18037 51399 18071
rect 54677 18037 54711 18071
rect 27077 17833 27111 17867
rect 30113 17833 30147 17867
rect 30573 17833 30607 17867
rect 32873 17833 32907 17867
rect 33517 17833 33551 17867
rect 33793 17833 33827 17867
rect 43637 17833 43671 17867
rect 45845 17833 45879 17867
rect 48421 17833 48455 17867
rect 51733 17833 51767 17867
rect 53389 17833 53423 17867
rect 54585 17833 54619 17867
rect 16221 17765 16255 17799
rect 19349 17765 19383 17799
rect 20545 17765 20579 17799
rect 20637 17765 20671 17799
rect 21465 17765 21499 17799
rect 25697 17765 25731 17799
rect 36461 17765 36495 17799
rect 46305 17765 46339 17799
rect 10701 17697 10735 17731
rect 13277 17697 13311 17731
rect 13461 17697 13495 17731
rect 18245 17697 18279 17731
rect 18705 17697 18739 17731
rect 20729 17697 20763 17731
rect 26985 17697 27019 17731
rect 31125 17697 31159 17731
rect 31401 17697 31435 17731
rect 41337 17697 41371 17731
rect 42441 17697 42475 17731
rect 42901 17697 42935 17731
rect 44741 17697 44775 17731
rect 45753 17697 45787 17731
rect 47409 17697 47443 17731
rect 10425 17629 10459 17663
rect 14473 17629 14507 17663
rect 16865 17629 16899 17663
rect 17509 17629 17543 17663
rect 18521 17629 18555 17663
rect 20177 17629 20211 17663
rect 21649 17629 21683 17663
rect 25972 17629 26006 17663
rect 26065 17629 26099 17663
rect 27261 17629 27295 17663
rect 27353 17629 27387 17663
rect 27537 17629 27571 17663
rect 27629 17629 27663 17663
rect 27813 17629 27847 17663
rect 27997 17629 28031 17663
rect 28089 17629 28123 17663
rect 28273 17629 28307 17663
rect 28365 17629 28399 17663
rect 29653 17629 29687 17663
rect 29929 17629 29963 17663
rect 33333 17629 33367 17663
rect 34897 17629 34931 17663
rect 34989 17629 35023 17663
rect 35265 17629 35299 17663
rect 36645 17629 36679 17663
rect 36829 17629 36863 17663
rect 37013 17629 37047 17663
rect 37105 17629 37139 17663
rect 38945 17629 38979 17663
rect 39221 17629 39255 17663
rect 39865 17629 39899 17663
rect 40013 17629 40047 17663
rect 40233 17629 40267 17663
rect 40330 17629 40364 17663
rect 41705 17629 41739 17663
rect 42257 17629 42291 17663
rect 42349 17629 42383 17663
rect 42625 17629 42659 17663
rect 42717 17629 42751 17663
rect 42993 17629 43027 17663
rect 43177 17629 43211 17663
rect 43361 17629 43395 17663
rect 46029 17629 46063 17663
rect 46121 17629 46155 17663
rect 46397 17629 46431 17663
rect 46765 17629 46799 17663
rect 47777 17629 47811 17663
rect 47870 17629 47904 17663
rect 48145 17629 48179 17663
rect 48242 17629 48276 17663
rect 51365 17629 51399 17663
rect 51549 17629 51583 17663
rect 52745 17629 52779 17663
rect 52838 17629 52872 17663
rect 53113 17629 53147 17663
rect 53210 17629 53244 17663
rect 53941 17629 53975 17663
rect 54034 17629 54068 17663
rect 54406 17629 54440 17663
rect 13185 17561 13219 17595
rect 14749 17561 14783 17595
rect 21833 17561 21867 17595
rect 30665 17561 30699 17595
rect 33057 17561 33091 17595
rect 35081 17561 35115 17595
rect 36737 17561 36771 17595
rect 38209 17561 38243 17595
rect 40141 17561 40175 17595
rect 40601 17561 40635 17595
rect 43269 17561 43303 17595
rect 48053 17561 48087 17595
rect 53021 17561 53055 17595
rect 54217 17561 54251 17595
rect 54309 17561 54343 17595
rect 12173 17493 12207 17527
rect 12817 17493 12851 17527
rect 16313 17493 16347 17527
rect 21005 17493 21039 17527
rect 29745 17493 29779 17527
rect 30205 17493 30239 17527
rect 33149 17493 33183 17527
rect 34713 17493 34747 17527
rect 35449 17493 35483 17527
rect 37289 17493 37323 17527
rect 37473 17493 37507 17527
rect 40509 17493 40543 17527
rect 43545 17493 43579 17527
rect 44189 17493 44223 17527
rect 47593 17493 47627 17527
rect 15117 17289 15151 17323
rect 15485 17289 15519 17323
rect 15577 17289 15611 17323
rect 23673 17289 23707 17323
rect 30665 17289 30699 17323
rect 31033 17289 31067 17323
rect 31493 17289 31527 17323
rect 32229 17289 32263 17323
rect 43177 17289 43211 17323
rect 46305 17289 46339 17323
rect 50077 17289 50111 17323
rect 52377 17289 52411 17323
rect 9781 17221 9815 17255
rect 30205 17221 30239 17255
rect 32689 17221 32723 17255
rect 42533 17221 42567 17255
rect 44925 17221 44959 17255
rect 45937 17221 45971 17255
rect 46029 17221 46063 17255
rect 54125 17221 54159 17255
rect 9505 17153 9539 17187
rect 12173 17153 12207 17187
rect 14197 17153 14231 17187
rect 16129 17153 16163 17187
rect 18889 17153 18923 17187
rect 23121 17153 23155 17187
rect 23305 17153 23339 17187
rect 23581 17153 23615 17187
rect 23765 17153 23799 17187
rect 27813 17153 27847 17187
rect 28089 17153 28123 17187
rect 28273 17153 28307 17187
rect 28549 17153 28583 17187
rect 29285 17153 29319 17187
rect 29469 17153 29503 17187
rect 30021 17153 30055 17187
rect 30297 17153 30331 17187
rect 30481 17153 30515 17187
rect 30757 17153 30791 17187
rect 31309 17153 31343 17187
rect 31953 17153 31987 17187
rect 32597 17153 32631 17187
rect 32781 17153 32815 17187
rect 32965 17153 32999 17187
rect 33149 17153 33183 17187
rect 33609 17153 33643 17187
rect 34437 17153 34471 17187
rect 34529 17153 34563 17187
rect 34805 17153 34839 17187
rect 36645 17153 36679 17187
rect 36737 17153 36771 17187
rect 37013 17153 37047 17187
rect 38025 17153 38059 17187
rect 38301 17153 38335 17187
rect 38577 17153 38611 17187
rect 41061 17153 41095 17187
rect 41337 17153 41371 17187
rect 43085 17153 43119 17187
rect 43361 17153 43395 17187
rect 43453 17153 43487 17187
rect 43729 17153 43763 17187
rect 45201 17153 45235 17187
rect 45293 17153 45327 17187
rect 45569 17153 45603 17187
rect 45753 17153 45787 17187
rect 46121 17153 46155 17187
rect 46397 17153 46431 17187
rect 48329 17153 48363 17187
rect 52193 17153 52227 17187
rect 53849 17153 53883 17187
rect 53942 17153 53976 17187
rect 54217 17153 54251 17187
rect 54355 17153 54389 17187
rect 78045 17153 78079 17187
rect 12449 17085 12483 17119
rect 13921 17085 13955 17119
rect 14289 17085 14323 17119
rect 15669 17085 15703 17119
rect 16221 17085 16255 17119
rect 17049 17085 17083 17119
rect 17325 17085 17359 17119
rect 18797 17085 18831 17119
rect 19441 17085 19475 17119
rect 20729 17085 20763 17119
rect 27721 17085 27755 17119
rect 29745 17085 29779 17119
rect 31033 17085 31067 17119
rect 33425 17085 33459 17119
rect 34713 17085 34747 17119
rect 38485 17085 38519 17119
rect 38853 17085 38887 17119
rect 40325 17085 40359 17119
rect 41153 17085 41187 17119
rect 45017 17085 45051 17119
rect 50537 17085 50571 17119
rect 20177 17017 20211 17051
rect 20545 17017 20579 17051
rect 23397 17017 23431 17051
rect 29101 17017 29135 17051
rect 41705 17017 41739 17051
rect 49893 17017 49927 17051
rect 78229 17017 78263 17051
rect 11253 16949 11287 16983
rect 14473 16949 14507 16983
rect 16405 16949 16439 16983
rect 20637 16949 20671 16983
rect 20821 16949 20855 16983
rect 29653 16949 29687 16983
rect 29837 16949 29871 16983
rect 30849 16949 30883 16983
rect 31217 16949 31251 16983
rect 31769 16949 31803 16983
rect 32413 16949 32447 16983
rect 33793 16949 33827 16983
rect 33977 16949 34011 16983
rect 34253 16949 34287 16983
rect 36461 16949 36495 16983
rect 36921 16949 36955 16983
rect 38117 16949 38151 16983
rect 41521 16949 41555 16983
rect 42257 16949 42291 16983
rect 43637 16949 43671 16983
rect 45477 16949 45511 16983
rect 48605 16949 48639 16983
rect 53757 16949 53791 16983
rect 54493 16949 54527 16983
rect 77861 16949 77895 16983
rect 12817 16745 12851 16779
rect 20453 16745 20487 16779
rect 25421 16745 25455 16779
rect 25697 16745 25731 16779
rect 28273 16745 28307 16779
rect 38025 16745 38059 16779
rect 38393 16745 38427 16779
rect 42809 16745 42843 16779
rect 45845 16745 45879 16779
rect 46029 16745 46063 16779
rect 46305 16745 46339 16779
rect 50813 16745 50847 16779
rect 55597 16745 55631 16779
rect 11713 16677 11747 16711
rect 20545 16677 20579 16711
rect 22937 16677 22971 16711
rect 25789 16677 25823 16711
rect 26249 16677 26283 16711
rect 27813 16677 27847 16711
rect 44833 16677 44867 16711
rect 46765 16677 46799 16711
rect 12633 16609 12667 16643
rect 18337 16609 18371 16643
rect 18981 16609 19015 16643
rect 20637 16609 20671 16643
rect 25881 16609 25915 16643
rect 28273 16609 28307 16643
rect 36461 16609 36495 16643
rect 41061 16609 41095 16643
rect 41337 16609 41371 16643
rect 43085 16609 43119 16643
rect 43361 16609 43395 16643
rect 45293 16609 45327 16643
rect 46857 16609 46891 16643
rect 47133 16609 47167 16643
rect 52009 16609 52043 16643
rect 52285 16609 52319 16643
rect 56517 16609 56551 16643
rect 10609 16541 10643 16575
rect 12541 16541 12575 16575
rect 18061 16541 18095 16575
rect 18889 16541 18923 16575
rect 20085 16541 20119 16575
rect 22753 16541 22787 16575
rect 22937 16541 22971 16575
rect 23029 16541 23063 16575
rect 23213 16541 23247 16575
rect 23489 16541 23523 16575
rect 23673 16541 23707 16575
rect 23949 16541 23983 16575
rect 24133 16541 24167 16575
rect 26157 16541 26191 16575
rect 26433 16541 26467 16575
rect 26801 16541 26835 16575
rect 27629 16541 27663 16575
rect 28365 16541 28399 16575
rect 31585 16541 31619 16575
rect 36185 16541 36219 16575
rect 38531 16541 38565 16575
rect 38761 16541 38795 16575
rect 38944 16541 38978 16575
rect 39037 16541 39071 16575
rect 46213 16541 46247 16575
rect 46489 16541 46523 16575
rect 46581 16541 46615 16575
rect 48881 16541 48915 16575
rect 49249 16541 49283 16575
rect 49525 16541 49559 16575
rect 49893 16541 49927 16575
rect 50169 16541 50203 16575
rect 50317 16541 50351 16575
rect 50537 16541 50571 16575
rect 50675 16541 50709 16575
rect 51089 16541 51123 16575
rect 51457 16541 51491 16575
rect 54401 16541 54435 16575
rect 54769 16541 54803 16575
rect 54953 16541 54987 16575
rect 55045 16541 55079 16575
rect 55781 16541 55815 16575
rect 55965 16541 55999 16575
rect 56057 16541 56091 16575
rect 56149 16541 56183 16575
rect 11437 16473 11471 16507
rect 18153 16473 18187 16507
rect 26525 16473 26559 16507
rect 26617 16473 26651 16507
rect 27445 16473 27479 16507
rect 28089 16473 28123 16507
rect 31861 16473 31895 16507
rect 38669 16473 38703 16507
rect 48973 16473 49007 16507
rect 49065 16473 49099 16507
rect 49617 16473 49651 16507
rect 49709 16473 49743 16507
rect 50445 16473 50479 16507
rect 51181 16473 51215 16507
rect 51273 16473 51307 16507
rect 56425 16473 56459 16507
rect 56762 16473 56796 16507
rect 17693 16405 17727 16439
rect 18521 16405 18555 16439
rect 20913 16405 20947 16439
rect 23305 16405 23339 16439
rect 23765 16405 23799 16439
rect 24041 16405 24075 16439
rect 26065 16405 26099 16439
rect 28549 16405 28583 16439
rect 33333 16405 33367 16439
rect 33517 16405 33551 16439
rect 37933 16405 37967 16439
rect 48605 16405 48639 16439
rect 48697 16405 48731 16439
rect 49341 16405 49375 16439
rect 50905 16405 50939 16439
rect 51549 16405 51583 16439
rect 53757 16405 53791 16439
rect 53849 16405 53883 16439
rect 54585 16405 54619 16439
rect 57897 16405 57931 16439
rect 13277 16201 13311 16235
rect 17049 16201 17083 16235
rect 17509 16201 17543 16235
rect 20821 16201 20855 16235
rect 24593 16201 24627 16235
rect 24777 16201 24811 16235
rect 26065 16201 26099 16235
rect 27997 16201 28031 16235
rect 32137 16201 32171 16235
rect 35633 16201 35667 16235
rect 44741 16201 44775 16235
rect 44925 16201 44959 16235
rect 46213 16201 46247 16235
rect 47317 16201 47351 16235
rect 47593 16201 47627 16235
rect 48789 16201 48823 16235
rect 52561 16201 52595 16235
rect 52745 16201 52779 16235
rect 57069 16201 57103 16235
rect 57989 16201 58023 16235
rect 17233 16133 17267 16167
rect 27445 16133 27479 16167
rect 34161 16133 34195 16167
rect 45385 16133 45419 16167
rect 46765 16133 46799 16167
rect 49065 16133 49099 16167
rect 49893 16133 49927 16167
rect 50721 16133 50755 16167
rect 52193 16133 52227 16167
rect 53389 16133 53423 16167
rect 54677 16133 54711 16167
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 8585 16065 8619 16099
rect 11529 16065 11563 16099
rect 17141 16065 17175 16099
rect 18061 16065 18095 16099
rect 20361 16065 20395 16099
rect 20545 16065 20579 16099
rect 20729 16065 20763 16099
rect 21097 16065 21131 16099
rect 23213 16065 23247 16099
rect 23397 16065 23431 16099
rect 23489 16065 23523 16099
rect 23673 16065 23707 16099
rect 24041 16065 24075 16099
rect 24652 16065 24686 16099
rect 25605 16065 25639 16099
rect 25789 16065 25823 16099
rect 25881 16065 25915 16099
rect 27261 16065 27295 16099
rect 27997 16065 28031 16099
rect 28181 16065 28215 16099
rect 28457 16065 28491 16099
rect 32321 16065 32355 16099
rect 32413 16065 32447 16099
rect 32689 16065 32723 16099
rect 33885 16065 33919 16099
rect 45109 16065 45143 16099
rect 45257 16065 45291 16099
rect 45477 16065 45511 16099
rect 45574 16065 45608 16099
rect 45845 16065 45879 16099
rect 46029 16065 46063 16099
rect 46305 16065 46339 16099
rect 46673 16065 46707 16099
rect 46857 16065 46891 16099
rect 47041 16065 47075 16099
rect 48237 16065 48271 16099
rect 48329 16065 48363 16099
rect 48605 16065 48639 16099
rect 49525 16065 49559 16099
rect 49801 16065 49835 16099
rect 50169 16065 50203 16099
rect 50465 16065 50499 16099
rect 50629 16065 50663 16099
rect 50859 16065 50893 16099
rect 51079 16065 51113 16099
rect 51181 16065 51215 16099
rect 51365 16065 51399 16099
rect 51457 16065 51491 16099
rect 51733 16065 51767 16099
rect 51917 16065 51951 16099
rect 52010 16065 52044 16099
rect 52285 16065 52319 16099
rect 52423 16065 52457 16099
rect 52929 16065 52963 16099
rect 53113 16065 53147 16099
rect 53205 16065 53239 16099
rect 57713 16065 57747 16099
rect 8861 15997 8895 16031
rect 11805 15997 11839 16031
rect 13645 15997 13679 16031
rect 13921 15997 13955 16031
rect 15393 15997 15427 16031
rect 16037 15997 16071 16031
rect 20913 15997 20947 16031
rect 24133 15997 24167 16031
rect 24225 15997 24259 16031
rect 32597 15997 32631 16031
rect 48421 15997 48455 16031
rect 50077 15997 50111 16031
rect 54125 15997 54159 16031
rect 54401 15997 54435 16031
rect 56149 15997 56183 16031
rect 1593 15929 1627 15963
rect 16865 15929 16899 15963
rect 23949 15929 23983 15963
rect 35817 15929 35851 15963
rect 45753 15929 45787 15963
rect 50353 15929 50387 15963
rect 50997 15929 51031 15963
rect 10333 15861 10367 15895
rect 15485 15861 15519 15895
rect 17417 15861 17451 15895
rect 20545 15861 20579 15895
rect 21097 15861 21131 15895
rect 23397 15861 23431 15895
rect 25881 15861 25915 15895
rect 27077 15861 27111 15895
rect 28641 15861 28675 15895
rect 36001 15861 36035 15895
rect 46489 15861 46523 15895
rect 47133 15861 47167 15895
rect 48605 15861 48639 15895
rect 49249 15861 49283 15895
rect 49985 15861 50019 15895
rect 51641 15861 51675 15895
rect 8309 15657 8343 15691
rect 11805 15657 11839 15691
rect 14289 15657 14323 15691
rect 16129 15657 16163 15691
rect 19717 15657 19751 15691
rect 20545 15657 20579 15691
rect 25237 15657 25271 15691
rect 25697 15657 25731 15691
rect 27905 15657 27939 15691
rect 29653 15657 29687 15691
rect 31493 15657 31527 15691
rect 34345 15657 34379 15691
rect 49893 15657 49927 15691
rect 50721 15657 50755 15691
rect 53297 15657 53331 15691
rect 19625 15589 19659 15623
rect 20085 15589 20119 15623
rect 28641 15589 28675 15623
rect 56149 15589 56183 15623
rect 12449 15521 12483 15555
rect 13369 15521 13403 15555
rect 14749 15521 14783 15555
rect 14933 15521 14967 15555
rect 15761 15521 15795 15555
rect 19809 15521 19843 15555
rect 20453 15521 20487 15555
rect 20545 15521 20579 15555
rect 21281 15521 21315 15555
rect 25329 15521 25363 15555
rect 35449 15521 35483 15555
rect 38117 15521 38151 15555
rect 38577 15521 38611 15555
rect 39865 15521 39899 15555
rect 46581 15521 46615 15555
rect 55781 15521 55815 15555
rect 1409 15453 1443 15487
rect 1685 15453 1719 15487
rect 8125 15453 8159 15487
rect 12173 15453 12207 15487
rect 14657 15453 14691 15487
rect 15853 15453 15887 15487
rect 19257 15453 19291 15487
rect 20361 15453 20395 15487
rect 20913 15453 20947 15487
rect 21097 15453 21131 15487
rect 21373 15453 21407 15487
rect 21649 15453 21683 15487
rect 22753 15453 22787 15487
rect 22845 15453 22879 15487
rect 23029 15453 23063 15487
rect 23213 15453 23247 15487
rect 25237 15453 25271 15487
rect 25513 15453 25547 15487
rect 26065 15453 26099 15487
rect 26433 15453 26467 15487
rect 26801 15453 26835 15487
rect 27261 15453 27295 15487
rect 27721 15453 27755 15487
rect 28365 15453 28399 15487
rect 28825 15453 28859 15487
rect 29009 15453 29043 15487
rect 29101 15453 29135 15487
rect 29193 15453 29227 15487
rect 29745 15453 29779 15487
rect 33517 15453 33551 15487
rect 33885 15453 33919 15487
rect 34069 15453 34103 15487
rect 34161 15453 34195 15487
rect 34713 15453 34747 15487
rect 35265 15453 35299 15487
rect 35633 15453 35667 15487
rect 35817 15453 35851 15487
rect 35909 15453 35943 15487
rect 36553 15453 36587 15487
rect 37105 15453 37139 15487
rect 37933 15453 37967 15487
rect 38209 15453 38243 15487
rect 38853 15453 38887 15487
rect 39405 15453 39439 15487
rect 41889 15453 41923 15487
rect 44281 15453 44315 15487
rect 49709 15453 49743 15487
rect 50169 15453 50203 15487
rect 50353 15453 50387 15487
rect 50445 15453 50479 15487
rect 50537 15453 50571 15487
rect 54309 15453 54343 15487
rect 54585 15453 54619 15487
rect 54677 15453 54711 15487
rect 55505 15453 55539 15487
rect 55597 15453 55631 15487
rect 55873 15453 55907 15487
rect 55965 15453 55999 15487
rect 20729 15385 20763 15419
rect 28457 15385 28491 15419
rect 28641 15385 28675 15419
rect 30021 15385 30055 15419
rect 32689 15385 32723 15419
rect 36001 15385 36035 15419
rect 36369 15385 36403 15419
rect 37381 15385 37415 15419
rect 37565 15385 37599 15419
rect 38393 15385 38427 15419
rect 38761 15385 38795 15419
rect 40141 15385 40175 15419
rect 42165 15385 42199 15419
rect 45661 15385 45695 15419
rect 45753 15385 45787 15419
rect 54493 15385 54527 15419
rect 1593 15317 1627 15351
rect 12265 15317 12299 15351
rect 12817 15317 12851 15351
rect 22661 15317 22695 15351
rect 23121 15317 23155 15351
rect 29377 15317 29411 15351
rect 33701 15317 33735 15351
rect 37749 15317 37783 15351
rect 41613 15317 41647 15351
rect 43637 15317 43671 15351
rect 43729 15317 43763 15351
rect 46765 15317 46799 15351
rect 50905 15317 50939 15351
rect 54861 15317 54895 15351
rect 55321 15317 55355 15351
rect 17233 15113 17267 15147
rect 25697 15113 25731 15147
rect 26341 15113 26375 15147
rect 29009 15113 29043 15147
rect 40233 15113 40267 15147
rect 42441 15113 42475 15147
rect 43361 15113 43395 15147
rect 47685 15113 47719 15147
rect 56609 15113 56643 15147
rect 19533 15045 19567 15079
rect 20545 15045 20579 15079
rect 24133 15045 24167 15079
rect 27353 15045 27387 15079
rect 27445 15045 27479 15079
rect 35541 15045 35575 15079
rect 37841 15045 37875 15079
rect 43637 15045 43671 15079
rect 55137 15045 55171 15079
rect 7573 14977 7607 15011
rect 7757 14977 7791 15011
rect 7941 14977 7975 15011
rect 8217 14977 8251 15011
rect 8769 14977 8803 15011
rect 9505 14977 9539 15011
rect 13001 14977 13035 15011
rect 16865 14977 16899 15011
rect 18613 14977 18647 15011
rect 22477 14977 22511 15011
rect 22661 14977 22695 15011
rect 22937 14977 22971 15011
rect 23121 14977 23155 15011
rect 23213 14977 23247 15011
rect 23397 14977 23431 15011
rect 23949 14977 23983 15011
rect 25329 14977 25363 15011
rect 25513 14977 25547 15011
rect 26249 14977 26283 15011
rect 26427 14977 26461 15011
rect 27077 14977 27111 15011
rect 27170 14977 27204 15011
rect 27583 14977 27617 15011
rect 28641 14977 28675 15011
rect 28917 14977 28951 15011
rect 29101 14977 29135 15011
rect 33241 14977 33275 15011
rect 35265 14977 35299 15011
rect 37289 14977 37323 15011
rect 37565 14977 37599 15011
rect 39497 14977 39531 15011
rect 39645 14977 39679 15011
rect 39773 14977 39807 15011
rect 39865 14977 39899 15011
rect 39962 14977 39996 15011
rect 40417 14977 40451 15011
rect 41061 14977 41095 15011
rect 41797 14977 41831 15011
rect 41981 14977 42015 15011
rect 42625 14977 42659 15011
rect 44281 14977 44315 15011
rect 46489 14977 46523 15011
rect 46857 14977 46891 15011
rect 48053 14977 48087 15011
rect 48145 14977 48179 15011
rect 48237 14977 48271 15011
rect 48421 14977 48455 15011
rect 49341 14977 49375 15011
rect 50537 14977 50571 15011
rect 50997 14977 51031 15011
rect 54861 14977 54895 15011
rect 8309 14909 8343 14943
rect 9781 14909 9815 14943
rect 11253 14909 11287 14943
rect 13093 14909 13127 14943
rect 16957 14909 16991 14943
rect 19165 14909 19199 14943
rect 19625 14909 19659 14943
rect 20177 14909 20211 14943
rect 32321 14909 32355 14943
rect 32597 14909 32631 14943
rect 33517 14909 33551 14943
rect 40693 14909 40727 14943
rect 41245 14909 41279 14943
rect 42901 14909 42935 14943
rect 44557 14909 44591 14943
rect 45109 14909 45143 14943
rect 45661 14909 45695 14943
rect 8953 14841 8987 14875
rect 20085 14841 20119 14875
rect 24317 14841 24351 14875
rect 28549 14841 28583 14875
rect 35081 14841 35115 14875
rect 40141 14841 40175 14875
rect 40601 14841 40635 14875
rect 42809 14841 42843 14875
rect 43913 14841 43947 14875
rect 13277 14773 13311 14807
rect 18981 14773 19015 14807
rect 19073 14773 19107 14807
rect 19993 14773 20027 14807
rect 22661 14773 22695 14807
rect 23121 14773 23155 14807
rect 23397 14773 23431 14807
rect 25329 14773 25363 14807
rect 27721 14773 27755 14807
rect 28733 14773 28767 14807
rect 34989 14773 35023 14807
rect 37013 14773 37047 14807
rect 39313 14773 39347 14807
rect 42165 14773 42199 14807
rect 44097 14773 44131 14807
rect 44465 14773 44499 14807
rect 46673 14773 46707 14807
rect 47869 14773 47903 14807
rect 49065 14773 49099 14807
rect 50261 14773 50295 14807
rect 50629 14773 50663 14807
rect 50905 14773 50939 14807
rect 54217 14773 54251 14807
rect 1593 14569 1627 14603
rect 14657 14569 14691 14603
rect 19625 14569 19659 14603
rect 19717 14569 19751 14603
rect 20085 14569 20119 14603
rect 22937 14569 22971 14603
rect 23213 14569 23247 14603
rect 28181 14569 28215 14603
rect 34161 14569 34195 14603
rect 35541 14569 35575 14603
rect 37289 14569 37323 14603
rect 42073 14569 42107 14603
rect 42993 14569 43027 14603
rect 44005 14569 44039 14603
rect 47501 14569 47535 14603
rect 53573 14569 53607 14603
rect 14105 14501 14139 14535
rect 27997 14501 28031 14535
rect 34805 14501 34839 14535
rect 44465 14501 44499 14535
rect 48329 14501 48363 14535
rect 12633 14433 12667 14467
rect 13461 14433 13495 14467
rect 14933 14433 14967 14467
rect 16681 14433 16715 14467
rect 17325 14433 17359 14467
rect 19809 14433 19843 14467
rect 20545 14433 20579 14467
rect 23029 14433 23063 14467
rect 23305 14433 23339 14467
rect 31309 14433 31343 14467
rect 37105 14433 37139 14467
rect 45753 14433 45787 14467
rect 49985 14433 50019 14467
rect 1409 14365 1443 14399
rect 1685 14365 1719 14399
rect 7665 14365 7699 14399
rect 12357 14365 12391 14399
rect 14289 14365 14323 14399
rect 14381 14365 14415 14399
rect 19257 14365 19291 14399
rect 20453 14365 20487 14399
rect 22753 14365 22787 14399
rect 23213 14365 23247 14399
rect 23673 14365 23707 14399
rect 27353 14365 27387 14399
rect 27446 14365 27480 14399
rect 27818 14365 27852 14399
rect 30297 14365 30331 14399
rect 30481 14365 30515 14399
rect 33149 14365 33183 14399
rect 33425 14365 33459 14399
rect 34989 14365 35023 14399
rect 35720 14365 35754 14399
rect 36092 14365 36126 14399
rect 36185 14365 36219 14399
rect 36277 14365 36311 14399
rect 36461 14365 36495 14399
rect 36645 14365 36679 14399
rect 37468 14365 37502 14399
rect 37657 14365 37691 14399
rect 37840 14365 37874 14399
rect 37933 14365 37967 14399
rect 41429 14365 41463 14399
rect 41522 14365 41556 14399
rect 41797 14365 41831 14399
rect 41935 14365 41969 14399
rect 42441 14365 42475 14399
rect 42533 14365 42567 14399
rect 42809 14365 42843 14399
rect 43361 14365 43395 14399
rect 43454 14365 43488 14399
rect 43729 14365 43763 14399
rect 43867 14365 43901 14399
rect 47685 14365 47719 14399
rect 47833 14365 47867 14399
rect 48150 14365 48184 14399
rect 48605 14365 48639 14399
rect 48789 14365 48823 14399
rect 48881 14365 48915 14399
rect 49341 14365 49375 14399
rect 50353 14365 50387 14399
rect 50445 14365 50479 14399
rect 50721 14365 50755 14399
rect 51096 14365 51130 14399
rect 51182 14365 51216 14399
rect 51457 14365 51491 14399
rect 51573 14365 51607 14399
rect 51825 14365 51859 14399
rect 54217 14365 54251 14399
rect 54580 14365 54614 14399
rect 54769 14365 54803 14399
rect 54952 14365 54986 14399
rect 55045 14365 55079 14399
rect 15209 14297 15243 14331
rect 17601 14297 17635 14331
rect 27629 14297 27663 14331
rect 27721 14297 27755 14331
rect 31585 14297 31619 14331
rect 35817 14297 35851 14331
rect 35909 14297 35943 14331
rect 36553 14297 36587 14331
rect 37565 14297 37599 14331
rect 41705 14297 41739 14331
rect 42625 14297 42659 14331
rect 43637 14297 43671 14331
rect 44189 14297 44223 14331
rect 44649 14297 44683 14331
rect 45017 14297 45051 14331
rect 45201 14297 45235 14331
rect 46029 14297 46063 14331
rect 47961 14297 47995 14331
rect 48053 14297 48087 14331
rect 50537 14297 50571 14331
rect 51365 14297 51399 14331
rect 52101 14297 52135 14331
rect 53665 14297 53699 14331
rect 54677 14297 54711 14331
rect 7849 14229 7883 14263
rect 11989 14229 12023 14263
rect 12449 14229 12483 14263
rect 12909 14229 12943 14263
rect 14473 14229 14507 14263
rect 16773 14229 16807 14263
rect 17693 14229 17727 14263
rect 18153 14229 18187 14263
rect 20821 14229 20855 14263
rect 22569 14229 22603 14263
rect 23581 14229 23615 14263
rect 23857 14229 23891 14263
rect 30113 14229 30147 14263
rect 33057 14229 33091 14263
rect 36829 14229 36863 14263
rect 36921 14229 36955 14263
rect 42257 14229 42291 14263
rect 43085 14229 43119 14263
rect 48421 14229 48455 14263
rect 50169 14229 50203 14263
rect 51733 14229 51767 14263
rect 54401 14229 54435 14263
rect 1593 14025 1627 14059
rect 13277 14025 13311 14059
rect 15761 14025 15795 14059
rect 16221 14025 16255 14059
rect 21465 14025 21499 14059
rect 22201 14025 22235 14059
rect 25789 14025 25823 14059
rect 28365 14025 28399 14059
rect 31493 14025 31527 14059
rect 32229 14025 32263 14059
rect 33149 14025 33183 14059
rect 46397 14025 46431 14059
rect 47133 14025 47167 14059
rect 47593 14025 47627 14059
rect 8217 13957 8251 13991
rect 11805 13957 11839 13991
rect 18429 13957 18463 13991
rect 24041 13957 24075 13991
rect 24685 13957 24719 13991
rect 25237 13957 25271 13991
rect 26341 13957 26375 13991
rect 27537 13957 27571 13991
rect 27905 13957 27939 13991
rect 32505 13957 32539 13991
rect 36277 13957 36311 13991
rect 36369 13957 36403 13991
rect 40877 13957 40911 13991
rect 44097 13957 44131 13991
rect 48145 13957 48179 13991
rect 1409 13889 1443 13923
rect 1685 13889 1719 13923
rect 11529 13889 11563 13923
rect 16129 13889 16163 13923
rect 17785 13889 17819 13923
rect 17969 13889 18003 13923
rect 18245 13889 18279 13923
rect 18521 13889 18555 13923
rect 21557 13889 21591 13923
rect 22385 13889 22419 13923
rect 22569 13889 22603 13923
rect 22661 13889 22695 13923
rect 22753 13889 22787 13923
rect 22937 13889 22971 13923
rect 23213 13889 23247 13923
rect 23673 13889 23707 13923
rect 23821 13889 23855 13923
rect 23949 13889 23983 13923
rect 24138 13889 24172 13923
rect 24409 13889 24443 13923
rect 24502 13889 24536 13923
rect 24777 13889 24811 13923
rect 24874 13889 24908 13923
rect 25145 13889 25179 13923
rect 25513 13889 25547 13923
rect 25605 13889 25639 13923
rect 26065 13889 26099 13923
rect 26157 13889 26191 13923
rect 27353 13889 27387 13923
rect 27445 13889 27479 13923
rect 27721 13889 27755 13923
rect 27813 13889 27847 13923
rect 28089 13889 28123 13923
rect 28181 13889 28215 13923
rect 31677 13889 31711 13923
rect 32408 13889 32442 13923
rect 32597 13889 32631 13923
rect 32780 13889 32814 13923
rect 32873 13889 32907 13923
rect 33931 13889 33965 13923
rect 34069 13889 34103 13923
rect 34161 13889 34195 13923
rect 34344 13889 34378 13923
rect 34437 13889 34471 13923
rect 36093 13889 36127 13923
rect 36461 13889 36495 13923
rect 36829 13889 36863 13923
rect 40601 13889 40635 13923
rect 40785 13889 40819 13923
rect 46581 13889 46615 13923
rect 46673 13889 46707 13923
rect 46949 13889 46983 13923
rect 49893 13889 49927 13923
rect 52009 13889 52043 13923
rect 52193 13889 52227 13923
rect 52469 13889 52503 13923
rect 53665 13889 53699 13923
rect 7941 13821 7975 13855
rect 9689 13821 9723 13855
rect 16405 13821 16439 13855
rect 23397 13821 23431 13855
rect 25973 13821 26007 13855
rect 29561 13821 29595 13855
rect 29837 13821 29871 13855
rect 31953 13821 31987 13855
rect 36921 13821 36955 13855
rect 40509 13821 40543 13855
rect 43821 13821 43855 13855
rect 47869 13821 47903 13855
rect 49617 13821 49651 13855
rect 50169 13821 50203 13855
rect 51641 13821 51675 13855
rect 24317 13753 24351 13787
rect 25053 13753 25087 13787
rect 25881 13753 25915 13787
rect 31309 13753 31343 13787
rect 40325 13753 40359 13787
rect 18153 13685 18187 13719
rect 18521 13685 18555 13719
rect 27169 13685 27203 13719
rect 27905 13685 27939 13719
rect 31861 13685 31895 13719
rect 33057 13685 33091 13719
rect 33793 13685 33827 13719
rect 36645 13685 36679 13719
rect 40049 13685 40083 13719
rect 40417 13685 40451 13719
rect 45569 13685 45603 13719
rect 46857 13685 46891 13719
rect 52377 13685 52411 13719
rect 53928 13685 53962 13719
rect 55413 13685 55447 13719
rect 18613 13481 18647 13515
rect 21557 13481 21591 13515
rect 21741 13481 21775 13515
rect 23213 13481 23247 13515
rect 27445 13481 27479 13515
rect 29193 13481 29227 13515
rect 29929 13481 29963 13515
rect 32505 13481 32539 13515
rect 37105 13481 37139 13515
rect 38945 13481 38979 13515
rect 39405 13481 39439 13515
rect 40417 13481 40451 13515
rect 40509 13481 40543 13515
rect 41521 13481 41555 13515
rect 43177 13481 43211 13515
rect 50169 13481 50203 13515
rect 53849 13481 53883 13515
rect 37197 13413 37231 13447
rect 37565 13413 37599 13447
rect 38761 13413 38795 13447
rect 39515 13413 39549 13447
rect 40785 13413 40819 13447
rect 43545 13413 43579 13447
rect 50629 13413 50663 13447
rect 54217 13413 54251 13447
rect 9045 13345 9079 13379
rect 19901 13345 19935 13379
rect 26617 13345 26651 13379
rect 26709 13345 26743 13379
rect 26801 13345 26835 13379
rect 26893 13345 26927 13379
rect 30205 13345 30239 13379
rect 30297 13345 30331 13379
rect 35265 13345 35299 13379
rect 37473 13345 37507 13379
rect 39313 13345 39347 13379
rect 40969 13345 41003 13379
rect 41337 13345 41371 13379
rect 54309 13345 54343 13379
rect 8585 13277 8619 13311
rect 17233 13277 17267 13311
rect 17325 13277 17359 13311
rect 17693 13277 17727 13311
rect 18061 13277 18095 13311
rect 19349 13277 19383 13311
rect 19717 13277 19751 13311
rect 23397 13277 23431 13311
rect 23581 13277 23615 13311
rect 23765 13277 23799 13311
rect 27353 13277 27387 13311
rect 28089 13277 28123 13311
rect 28273 13277 28307 13311
rect 28457 13277 28491 13311
rect 28733 13277 28767 13311
rect 29101 13277 29135 13311
rect 30113 13277 30147 13311
rect 30389 13277 30423 13311
rect 35081 13277 35115 13311
rect 35357 13277 35391 13311
rect 35817 13277 35851 13311
rect 36369 13277 36403 13311
rect 36737 13277 36771 13311
rect 37013 13277 37047 13311
rect 38117 13277 38151 13311
rect 38210 13277 38244 13311
rect 38393 13277 38427 13311
rect 38582 13277 38616 13311
rect 39129 13277 39163 13311
rect 39681 13277 39715 13311
rect 39865 13277 39899 13311
rect 40049 13277 40083 13311
rect 40233 13277 40267 13311
rect 41153 13277 41187 13311
rect 42993 13277 43027 13311
rect 43269 13277 43303 13311
rect 43913 13277 43947 13311
rect 44465 13277 44499 13311
rect 45017 13277 45051 13311
rect 45110 13277 45144 13311
rect 45293 13277 45327 13311
rect 45482 13277 45516 13311
rect 50353 13277 50387 13311
rect 50445 13277 50479 13311
rect 50721 13277 50755 13311
rect 54033 13277 54067 13311
rect 9321 13209 9355 13243
rect 16957 13209 16991 13243
rect 18429 13209 18463 13243
rect 18629 13209 18663 13243
rect 21373 13209 21407 13243
rect 23489 13209 23523 13243
rect 27997 13209 28031 13243
rect 28917 13209 28951 13243
rect 32413 13209 32447 13243
rect 38485 13209 38519 13243
rect 40141 13209 40175 13243
rect 43729 13209 43763 13243
rect 45385 13209 45419 13243
rect 8769 13141 8803 13175
rect 10793 13141 10827 13175
rect 18797 13141 18831 13175
rect 19441 13141 19475 13175
rect 21578 13141 21612 13175
rect 23949 13141 23983 13175
rect 26433 13141 26467 13175
rect 32137 13141 32171 13175
rect 34897 13141 34931 13175
rect 36829 13141 36863 13175
rect 39129 13141 39163 13175
rect 42809 13141 42843 13175
rect 44649 13141 44683 13175
rect 45661 13141 45695 13175
rect 13829 12937 13863 12971
rect 15025 12937 15059 12971
rect 22201 12937 22235 12971
rect 22477 12937 22511 12971
rect 33241 12937 33275 12971
rect 36277 12937 36311 12971
rect 37105 12937 37139 12971
rect 37841 12937 37875 12971
rect 38853 12937 38887 12971
rect 19625 12869 19659 12903
rect 22109 12869 22143 12903
rect 31033 12869 31067 12903
rect 31249 12869 31283 12903
rect 31861 12869 31895 12903
rect 32413 12869 32447 12903
rect 34713 12869 34747 12903
rect 37473 12869 37507 12903
rect 37565 12869 37599 12903
rect 38025 12869 38059 12903
rect 42993 12869 43027 12903
rect 45017 12869 45051 12903
rect 13921 12801 13955 12835
rect 14289 12801 14323 12835
rect 15393 12801 15427 12835
rect 17141 12801 17175 12835
rect 18061 12801 18095 12835
rect 18337 12801 18371 12835
rect 18613 12801 18647 12835
rect 18797 12801 18831 12835
rect 18889 12801 18923 12835
rect 19073 12801 19107 12835
rect 19349 12801 19383 12835
rect 19809 12801 19843 12835
rect 19901 12801 19935 12835
rect 20085 12801 20119 12835
rect 20821 12801 20855 12835
rect 22318 12801 22352 12835
rect 25421 12801 25455 12835
rect 25513 12801 25547 12835
rect 25697 12801 25731 12835
rect 25789 12801 25823 12835
rect 31677 12801 31711 12835
rect 31953 12801 31987 12835
rect 33333 12801 33367 12835
rect 33609 12801 33643 12835
rect 36645 12801 36679 12835
rect 36921 12801 36955 12835
rect 37289 12801 37323 12835
rect 37657 12801 37691 12835
rect 38209 12801 38243 12835
rect 40601 12801 40635 12835
rect 42717 12801 42751 12835
rect 44649 12801 44683 12835
rect 45109 12801 45143 12835
rect 50813 12801 50847 12835
rect 51181 12801 51215 12835
rect 14105 12733 14139 12767
rect 14933 12733 14967 12767
rect 15301 12733 15335 12767
rect 17877 12733 17911 12767
rect 19533 12733 19567 12767
rect 21833 12733 21867 12767
rect 33057 12733 33091 12767
rect 34437 12733 34471 12767
rect 36737 12733 36771 12767
rect 40785 12733 40819 12767
rect 40877 12733 40911 12767
rect 41337 12733 41371 12767
rect 41981 12733 42015 12767
rect 44465 12733 44499 12767
rect 45385 12733 45419 12767
rect 18521 12665 18555 12699
rect 20177 12665 20211 12699
rect 31401 12665 31435 12699
rect 13461 12597 13495 12631
rect 17693 12597 17727 12631
rect 20913 12597 20947 12631
rect 25237 12597 25271 12631
rect 31217 12597 31251 12631
rect 31493 12597 31527 12631
rect 36185 12597 36219 12631
rect 40417 12597 40451 12631
rect 46857 12597 46891 12631
rect 50997 12597 51031 12631
rect 14197 12393 14231 12427
rect 17003 12393 17037 12427
rect 19809 12393 19843 12427
rect 23673 12393 23707 12427
rect 24501 12393 24535 12427
rect 25697 12393 25731 12427
rect 32873 12393 32907 12427
rect 35633 12393 35667 12427
rect 42165 12393 42199 12427
rect 42901 12393 42935 12427
rect 44465 12393 44499 12427
rect 45293 12393 45327 12427
rect 45661 12393 45695 12427
rect 37473 12325 37507 12359
rect 15209 12257 15243 12291
rect 17877 12257 17911 12291
rect 25053 12257 25087 12291
rect 25973 12257 26007 12291
rect 27261 12257 27295 12291
rect 27353 12257 27387 12291
rect 27537 12257 27571 12291
rect 31401 12257 31435 12291
rect 40693 12257 40727 12291
rect 46949 12257 46983 12291
rect 50353 12257 50387 12291
rect 52469 12257 52503 12291
rect 14473 12189 14507 12223
rect 15577 12189 15611 12223
rect 18153 12189 18187 12223
rect 18337 12189 18371 12223
rect 19717 12189 19751 12223
rect 19901 12189 19935 12223
rect 21189 12189 21223 12223
rect 23489 12189 23523 12223
rect 23765 12189 23799 12223
rect 24133 12189 24167 12223
rect 24409 12189 24443 12223
rect 24593 12189 24627 12223
rect 25881 12189 25915 12223
rect 26157 12189 26191 12223
rect 26249 12189 26283 12223
rect 27445 12189 27479 12223
rect 27721 12189 27755 12223
rect 27905 12189 27939 12223
rect 27997 12189 28031 12223
rect 28089 12189 28123 12223
rect 28457 12189 28491 12223
rect 28549 12189 28583 12223
rect 28733 12189 28767 12223
rect 28825 12189 28859 12223
rect 31125 12189 31159 12223
rect 33057 12189 33091 12223
rect 33150 12189 33184 12223
rect 33333 12189 33367 12223
rect 33425 12189 33459 12223
rect 33522 12189 33556 12223
rect 33977 12189 34011 12223
rect 34161 12189 34195 12223
rect 34253 12189 34287 12223
rect 34989 12189 35023 12223
rect 35082 12189 35116 12223
rect 35265 12189 35299 12223
rect 35495 12189 35529 12223
rect 37289 12189 37323 12223
rect 37749 12189 37783 12223
rect 37842 12189 37876 12223
rect 38117 12189 38151 12223
rect 38214 12189 38248 12223
rect 40417 12189 40451 12223
rect 42257 12189 42291 12223
rect 42350 12189 42384 12223
rect 42625 12189 42659 12223
rect 42722 12189 42756 12223
rect 45477 12189 45511 12223
rect 45753 12189 45787 12223
rect 46397 12189 46431 12223
rect 47133 12189 47167 12223
rect 55413 12189 55447 12223
rect 55597 12189 55631 12223
rect 55965 12189 55999 12223
rect 56149 12189 56183 12223
rect 17141 12121 17175 12155
rect 18429 12121 18463 12155
rect 25329 12121 25363 12155
rect 26433 12121 26467 12155
rect 28365 12121 28399 12155
rect 33793 12121 33827 12155
rect 35357 12121 35391 12155
rect 38025 12121 38059 12155
rect 42533 12121 42567 12155
rect 47409 12121 47443 12155
rect 50629 12121 50663 12155
rect 52745 12121 52779 12155
rect 18245 12053 18279 12087
rect 21097 12053 21131 12087
rect 23305 12053 23339 12087
rect 23949 12053 23983 12087
rect 25237 12053 25271 12087
rect 27077 12053 27111 12087
rect 29009 12053 29043 12087
rect 29193 12053 29227 12087
rect 33701 12053 33735 12087
rect 38393 12053 38427 12087
rect 48881 12053 48915 12087
rect 52101 12053 52135 12087
rect 54217 12053 54251 12087
rect 56241 12053 56275 12087
rect 14473 11849 14507 11883
rect 17049 11849 17083 11883
rect 22937 11849 22971 11883
rect 34345 11849 34379 11883
rect 40417 11849 40451 11883
rect 47685 11849 47719 11883
rect 48329 11849 48363 11883
rect 49709 11849 49743 11883
rect 50721 11849 50755 11883
rect 13001 11781 13035 11815
rect 17325 11781 17359 11815
rect 17417 11781 17451 11815
rect 17555 11781 17589 11815
rect 26065 11781 26099 11815
rect 33977 11781 34011 11815
rect 48697 11781 48731 11815
rect 49433 11781 49467 11815
rect 49801 11781 49835 11815
rect 12725 11713 12759 11747
rect 17233 11713 17267 11747
rect 17693 11713 17727 11747
rect 22661 11713 22695 11747
rect 22845 11713 22879 11747
rect 23213 11713 23247 11747
rect 23305 11713 23339 11747
rect 23673 11713 23707 11747
rect 23949 11713 23983 11747
rect 24317 11713 24351 11747
rect 24501 11713 24535 11747
rect 25237 11713 25271 11747
rect 25421 11713 25455 11747
rect 25605 11713 25639 11747
rect 27445 11713 27479 11747
rect 27537 11713 27571 11747
rect 27629 11713 27663 11747
rect 27721 11713 27755 11747
rect 28181 11713 28215 11747
rect 29469 11713 29503 11747
rect 34253 11713 34287 11747
rect 36640 11713 36674 11747
rect 36737 11713 36771 11747
rect 36829 11713 36863 11747
rect 36957 11713 36991 11747
rect 37105 11713 37139 11747
rect 37841 11713 37875 11747
rect 38393 11713 38427 11747
rect 39773 11713 39807 11747
rect 39866 11713 39900 11747
rect 40049 11713 40083 11747
rect 40138 11713 40172 11747
rect 40238 11713 40272 11747
rect 47869 11713 47903 11747
rect 47961 11713 47995 11747
rect 48237 11713 48271 11747
rect 48513 11713 48547 11747
rect 48605 11713 48639 11747
rect 48881 11713 48915 11747
rect 49157 11713 49191 11747
rect 49341 11713 49375 11747
rect 49525 11713 49559 11747
rect 50077 11713 50111 11747
rect 50905 11713 50939 11747
rect 50997 11713 51031 11747
rect 51273 11713 51307 11747
rect 51733 11713 51767 11747
rect 52285 11713 52319 11747
rect 53021 11713 53055 11747
rect 54217 11713 54251 11747
rect 22753 11645 22787 11679
rect 24225 11645 24259 11679
rect 24409 11645 24443 11679
rect 25881 11645 25915 11679
rect 25973 11645 26007 11679
rect 27905 11645 27939 11679
rect 29745 11645 29779 11679
rect 36277 11645 36311 11679
rect 37289 11645 37323 11679
rect 38669 11645 38703 11679
rect 39037 11645 39071 11679
rect 39589 11645 39623 11679
rect 48973 11645 49007 11679
rect 49893 11645 49927 11679
rect 52745 11645 52779 11679
rect 54493 11645 54527 11679
rect 17877 11509 17911 11543
rect 23397 11509 23431 11543
rect 23489 11509 23523 11543
rect 23765 11509 23799 11543
rect 24133 11509 24167 11543
rect 26433 11509 26467 11543
rect 27261 11509 27295 11543
rect 31217 11509 31251 11543
rect 32505 11509 32539 11543
rect 36461 11509 36495 11543
rect 38209 11509 38243 11543
rect 38577 11509 38611 11543
rect 48145 11509 48179 11543
rect 49801 11509 49835 11543
rect 50261 11509 50295 11543
rect 51181 11509 51215 11543
rect 52469 11509 52503 11543
rect 55965 11509 55999 11543
rect 18889 11305 18923 11339
rect 23305 11305 23339 11339
rect 23489 11305 23523 11339
rect 26801 11305 26835 11339
rect 27813 11305 27847 11339
rect 29745 11305 29779 11339
rect 42257 11305 42291 11339
rect 44005 11305 44039 11339
rect 45661 11305 45695 11339
rect 48329 11305 48363 11339
rect 49065 11305 49099 11339
rect 51365 11305 51399 11339
rect 54493 11305 54527 11339
rect 54953 11305 54987 11339
rect 22385 11237 22419 11271
rect 37473 11237 37507 11271
rect 39681 11237 39715 11271
rect 52561 11237 52595 11271
rect 17141 11169 17175 11203
rect 17417 11169 17451 11203
rect 20637 11169 20671 11203
rect 25513 11169 25547 11203
rect 27905 11169 27939 11203
rect 30297 11169 30331 11203
rect 35725 11169 35759 11203
rect 37933 11169 37967 11203
rect 38209 11169 38243 11203
rect 53113 11169 53147 11203
rect 54217 11169 54251 11203
rect 22477 11101 22511 11135
rect 25789 11101 25823 11135
rect 26341 11101 26375 11135
rect 26433 11101 26467 11135
rect 26617 11101 26651 11135
rect 27813 11101 27847 11135
rect 30113 11101 30147 11135
rect 30665 11101 30699 11135
rect 42073 11101 42107 11135
rect 42349 11101 42383 11135
rect 42993 11101 43027 11135
rect 43545 11101 43579 11135
rect 43913 11101 43947 11135
rect 44189 11101 44223 11135
rect 44281 11101 44315 11135
rect 48605 11101 48639 11135
rect 51549 11101 51583 11135
rect 51641 11101 51675 11135
rect 52009 11101 52043 11135
rect 52285 11101 52319 11135
rect 52377 11101 52411 11135
rect 52653 11101 52687 11135
rect 52837 11101 52871 11135
rect 52929 11101 52963 11135
rect 53205 11101 53239 11135
rect 53665 11101 53699 11135
rect 54677 11101 54711 11135
rect 54769 11101 54803 11135
rect 55045 11101 55079 11135
rect 19073 11033 19107 11067
rect 20913 11033 20947 11067
rect 23121 11033 23155 11067
rect 23321 11033 23355 11067
rect 28273 11033 28307 11067
rect 28457 11033 28491 11067
rect 30205 11033 30239 11067
rect 36001 11033 36035 11067
rect 44557 11033 44591 11067
rect 45385 11033 45419 11067
rect 48789 11033 48823 11067
rect 52193 11033 52227 11067
rect 26249 10965 26283 10999
rect 28181 10965 28215 10999
rect 28641 10965 28675 10999
rect 41889 10965 41923 10999
rect 42441 10965 42475 10999
rect 44465 10965 44499 10999
rect 45845 10965 45879 10999
rect 19625 10761 19659 10795
rect 19717 10761 19751 10795
rect 32781 10761 32815 10795
rect 36277 10761 36311 10795
rect 39497 10761 39531 10795
rect 42073 10761 42107 10795
rect 43913 10761 43947 10795
rect 45753 10761 45787 10795
rect 49341 10761 49375 10795
rect 50261 10761 50295 10795
rect 54769 10761 54803 10795
rect 32505 10693 32539 10727
rect 41705 10693 41739 10727
rect 44281 10693 44315 10727
rect 46213 10693 46247 10727
rect 46305 10693 46339 10727
rect 50813 10693 50847 10727
rect 51825 10693 51859 10727
rect 54401 10693 54435 10727
rect 17877 10625 17911 10659
rect 26157 10625 26191 10659
rect 26341 10625 26375 10659
rect 26617 10625 26651 10659
rect 28641 10625 28675 10659
rect 28825 10625 28859 10659
rect 29561 10625 29595 10659
rect 32965 10625 32999 10659
rect 33149 10625 33183 10659
rect 33241 10625 33275 10659
rect 33333 10625 33367 10659
rect 36461 10625 36495 10659
rect 36645 10625 36679 10659
rect 36737 10625 36771 10659
rect 37841 10625 37875 10659
rect 38853 10625 38887 10659
rect 41429 10625 41463 10659
rect 41577 10625 41611 10659
rect 41797 10625 41831 10659
rect 41935 10625 41969 10659
rect 42717 10625 42751 10659
rect 43361 10625 43395 10659
rect 43545 10625 43579 10659
rect 43637 10625 43671 10659
rect 43729 10625 43763 10659
rect 46116 10625 46150 10659
rect 46488 10625 46522 10659
rect 46581 10625 46615 10659
rect 47593 10625 47627 10659
rect 49985 10625 50019 10659
rect 51089 10625 51123 10659
rect 54217 10625 54251 10659
rect 54493 10625 54527 10659
rect 54585 10625 54619 10659
rect 18153 10557 18187 10591
rect 21189 10557 21223 10591
rect 21465 10557 21499 10591
rect 28733 10557 28767 10591
rect 28917 10557 28951 10591
rect 29377 10557 29411 10591
rect 29745 10557 29779 10591
rect 33609 10557 33643 10591
rect 33885 10557 33919 10591
rect 35357 10557 35391 10591
rect 38577 10557 38611 10591
rect 42165 10557 42199 10591
rect 42441 10557 42475 10591
rect 44005 10557 44039 10591
rect 47869 10557 47903 10591
rect 45937 10489 45971 10523
rect 46673 10489 46707 10523
rect 21649 10421 21683 10455
rect 26801 10421 26835 10455
rect 28457 10421 28491 10455
rect 32413 10421 32447 10455
rect 33517 10421 33551 10455
rect 49433 10421 49467 10455
rect 50353 10421 50387 10455
rect 50997 10421 51031 10455
rect 54861 10421 54895 10455
rect 25421 10217 25455 10251
rect 32781 10217 32815 10251
rect 32965 10217 32999 10251
rect 33885 10217 33919 10251
rect 39681 10217 39715 10251
rect 43545 10217 43579 10251
rect 47961 10217 47995 10251
rect 48421 10217 48455 10251
rect 48605 10217 48639 10251
rect 50169 10217 50203 10251
rect 39497 10149 39531 10183
rect 49893 10149 49927 10183
rect 26341 10081 26375 10115
rect 32689 10081 32723 10115
rect 35265 10081 35299 10115
rect 39957 10081 39991 10115
rect 41797 10081 41831 10115
rect 45293 10081 45327 10115
rect 47041 10081 47075 10115
rect 52653 10081 52687 10115
rect 55321 10081 55355 10115
rect 57069 10081 57103 10115
rect 25605 10013 25639 10047
rect 26617 10013 26651 10047
rect 26801 10013 26835 10047
rect 26985 10013 27019 10047
rect 30941 10013 30975 10047
rect 33517 10013 33551 10047
rect 34529 10013 34563 10047
rect 38848 10013 38882 10047
rect 39037 10013 39071 10047
rect 39220 10013 39254 10047
rect 39313 10013 39347 10047
rect 43821 10013 43855 10047
rect 44097 10013 44131 10047
rect 47685 10013 47719 10047
rect 48145 10013 48179 10047
rect 48237 10013 48271 10047
rect 48513 10013 48547 10047
rect 48789 10013 48823 10047
rect 48881 10013 48915 10047
rect 49157 10013 49191 10047
rect 49249 10013 49283 10047
rect 49525 10013 49559 10047
rect 49617 10013 49651 10047
rect 50353 10013 50387 10047
rect 50446 10013 50480 10047
rect 50629 10013 50663 10047
rect 50721 10013 50755 10047
rect 50818 10013 50852 10047
rect 51268 10013 51302 10047
rect 51457 10013 51491 10047
rect 51585 10013 51619 10047
rect 51733 10013 51767 10047
rect 51917 10013 51951 10047
rect 52010 10013 52044 10047
rect 52382 10013 52416 10047
rect 55045 10013 55079 10047
rect 26893 9945 26927 9979
rect 31217 9945 31251 9979
rect 38945 9945 38979 9979
rect 40233 9945 40267 9979
rect 42073 9945 42107 9979
rect 44005 9945 44039 9979
rect 45569 9945 45603 9979
rect 48973 9945 49007 9979
rect 49433 9945 49467 9979
rect 51365 9945 51399 9979
rect 52193 9945 52227 9979
rect 52285 9945 52319 9979
rect 52929 9945 52963 9979
rect 54493 9945 54527 9979
rect 55597 9945 55631 9979
rect 19717 9877 19751 9911
rect 27169 9877 27203 9911
rect 34713 9877 34747 9911
rect 38669 9877 38703 9911
rect 41705 9877 41739 9911
rect 47133 9877 47167 9911
rect 49801 9877 49835 9911
rect 50997 9877 51031 9911
rect 51089 9877 51123 9911
rect 52561 9877 52595 9911
rect 54401 9877 54435 9911
rect 57161 9877 57195 9911
rect 27353 9673 27387 9707
rect 31401 9673 31435 9707
rect 40785 9673 40819 9707
rect 45661 9673 45695 9707
rect 49801 9673 49835 9707
rect 50169 9673 50203 9707
rect 51365 9673 51399 9707
rect 51917 9673 51951 9707
rect 52837 9673 52871 9707
rect 55689 9673 55723 9707
rect 28365 9605 28399 9639
rect 35725 9605 35759 9639
rect 40601 9605 40635 9639
rect 42717 9605 42751 9639
rect 43913 9605 43947 9639
rect 48973 9605 49007 9639
rect 50445 9605 50479 9639
rect 50537 9605 50571 9639
rect 50997 9605 51031 9639
rect 51089 9605 51123 9639
rect 51641 9605 51675 9639
rect 28089 9537 28123 9571
rect 31585 9537 31619 9571
rect 31677 9537 31711 9571
rect 31953 9537 31987 9571
rect 32689 9537 32723 9571
rect 33977 9537 34011 9571
rect 34069 9537 34103 9571
rect 34345 9537 34379 9571
rect 34989 9537 35023 9571
rect 35173 9537 35207 9571
rect 35265 9537 35299 9571
rect 35357 9537 35391 9571
rect 37657 9537 37691 9571
rect 40509 9537 40543 9571
rect 40969 9537 41003 9571
rect 41061 9537 41095 9571
rect 41337 9537 41371 9571
rect 41521 9537 41555 9571
rect 42625 9537 42659 9571
rect 42809 9537 42843 9571
rect 42993 9537 43027 9571
rect 43264 9537 43298 9571
rect 43361 9537 43395 9571
rect 43453 9537 43487 9571
rect 43581 9537 43615 9571
rect 43729 9537 43763 9571
rect 45845 9537 45879 9571
rect 45937 9537 45971 9571
rect 46213 9537 46247 9571
rect 48881 9537 48915 9571
rect 49065 9537 49099 9571
rect 49249 9537 49283 9571
rect 49341 9537 49375 9571
rect 50353 9537 50387 9571
rect 50721 9537 50755 9571
rect 50813 9537 50847 9571
rect 51181 9537 51215 9571
rect 51457 9537 51491 9571
rect 53021 9537 53055 9571
rect 53297 9537 53331 9571
rect 54493 9537 54527 9571
rect 54677 9537 54711 9571
rect 54769 9537 54803 9571
rect 54861 9537 54895 9571
rect 55183 9537 55217 9571
rect 55413 9537 55447 9571
rect 55505 9537 55539 9571
rect 56609 9537 56643 9571
rect 27997 9469 28031 9503
rect 29929 9469 29963 9503
rect 33333 9469 33367 9503
rect 37933 9469 37967 9503
rect 40049 9469 40083 9503
rect 42165 9469 42199 9503
rect 33793 9401 33827 9435
rect 42441 9401 42475 9435
rect 49525 9401 49559 9435
rect 56057 9401 56091 9435
rect 29837 9333 29871 9367
rect 31861 9333 31895 9367
rect 34253 9333 34287 9367
rect 35541 9333 35575 9367
rect 35909 9333 35943 9367
rect 39405 9333 39439 9367
rect 39497 9333 39531 9367
rect 40325 9333 40359 9367
rect 41245 9333 41279 9367
rect 43085 9333 43119 9367
rect 46121 9333 46155 9367
rect 48697 9333 48731 9367
rect 49893 9333 49927 9367
rect 53205 9333 53239 9367
rect 55045 9333 55079 9367
rect 55229 9333 55263 9367
rect 28273 9129 28307 9163
rect 31861 9129 31895 9163
rect 34529 9129 34563 9163
rect 38209 9129 38243 9163
rect 42901 9129 42935 9163
rect 49249 9129 49283 9163
rect 49709 9129 49743 9163
rect 50629 9129 50663 9163
rect 51273 9129 51307 9163
rect 37289 9061 37323 9095
rect 38669 9061 38703 9095
rect 43637 9061 43671 9095
rect 50445 9061 50479 9095
rect 26525 8993 26559 9027
rect 26801 8993 26835 9027
rect 32781 8993 32815 9027
rect 35265 8993 35299 9027
rect 37381 8993 37415 9027
rect 43453 8993 43487 9027
rect 49801 8993 49835 9027
rect 51365 8993 51399 9027
rect 30757 8925 30791 8959
rect 31125 8925 31159 8959
rect 31309 8925 31343 8959
rect 31493 8925 31527 8959
rect 31677 8925 31711 8959
rect 32045 8925 32079 8959
rect 32193 8925 32227 8959
rect 32410 8925 32444 8959
rect 32549 8925 32583 8959
rect 35909 8925 35943 8959
rect 36002 8925 36036 8959
rect 36277 8925 36311 8959
rect 36374 8925 36408 8959
rect 36645 8925 36679 8959
rect 36738 8925 36772 8959
rect 37110 8925 37144 8959
rect 37565 8925 37599 8959
rect 38393 8925 38427 8959
rect 38485 8925 38519 8959
rect 38761 8925 38795 8959
rect 41981 8925 42015 8959
rect 42073 8925 42107 8959
rect 43959 8925 43993 8959
rect 44097 8925 44131 8959
rect 44372 8925 44406 8959
rect 44465 8925 44499 8959
rect 50813 8925 50847 8959
rect 51181 8925 51215 8959
rect 51273 8925 51307 8959
rect 51549 8925 51583 8959
rect 31585 8857 31619 8891
rect 32321 8857 32355 8891
rect 33057 8857 33091 8891
rect 36185 8857 36219 8891
rect 36921 8857 36955 8891
rect 37013 8857 37047 8891
rect 44189 8857 44223 8891
rect 45385 8857 45419 8891
rect 50905 8857 50939 8891
rect 50997 8857 51031 8891
rect 28365 8789 28399 8823
rect 30941 8789 30975 8823
rect 32689 8789 32723 8823
rect 34713 8789 34747 8823
rect 36553 8789 36587 8823
rect 41337 8789 41371 8823
rect 42257 8789 42291 8823
rect 43821 8789 43855 8823
rect 50169 8789 50203 8823
rect 51733 8789 51767 8823
rect 31585 8585 31619 8619
rect 32873 8585 32907 8619
rect 36461 8585 36495 8619
rect 38761 8585 38795 8619
rect 43453 8585 43487 8619
rect 45477 8585 45511 8619
rect 45661 8585 45695 8619
rect 49525 8585 49559 8619
rect 50997 8585 51031 8619
rect 51181 8585 51215 8619
rect 31217 8517 31251 8551
rect 36737 8517 36771 8551
rect 37105 8517 37139 8551
rect 37289 8517 37323 8551
rect 38393 8517 38427 8551
rect 41245 8517 41279 8551
rect 41337 8517 41371 8551
rect 43913 8517 43947 8551
rect 44281 8517 44315 8551
rect 45017 8517 45051 8551
rect 50629 8517 50663 8551
rect 50721 8517 50755 8551
rect 51549 8517 51583 8551
rect 28917 8449 28951 8483
rect 31028 8449 31062 8483
rect 31125 8449 31159 8483
rect 31400 8449 31434 8483
rect 31493 8449 31527 8483
rect 33057 8449 33091 8483
rect 33333 8449 33367 8483
rect 35081 8449 35115 8483
rect 35174 8449 35208 8483
rect 35357 8449 35391 8483
rect 35449 8449 35483 8483
rect 35587 8449 35621 8483
rect 35817 8449 35851 8483
rect 35910 8449 35944 8483
rect 36093 8449 36127 8483
rect 36185 8449 36219 8483
rect 36282 8449 36316 8483
rect 37473 8449 37507 8483
rect 37565 8449 37599 8483
rect 38209 8449 38243 8483
rect 38485 8449 38519 8483
rect 38577 8449 38611 8483
rect 40601 8449 40635 8483
rect 41148 8449 41182 8483
rect 41520 8449 41554 8483
rect 41613 8449 41647 8483
rect 42441 8449 42475 8483
rect 42625 8449 42659 8483
rect 42718 8449 42752 8483
rect 42901 8449 42935 8483
rect 42993 8449 43027 8483
rect 43090 8449 43124 8483
rect 43637 8449 43671 8483
rect 44005 8449 44039 8483
rect 44189 8449 44223 8483
rect 44373 8449 44407 8483
rect 44649 8449 44683 8483
rect 44742 8449 44776 8483
rect 44925 8449 44959 8483
rect 45114 8449 45148 8483
rect 48789 8449 48823 8483
rect 48881 8449 48915 8483
rect 49157 8449 49191 8483
rect 49617 8449 49651 8483
rect 50353 8449 50387 8483
rect 50501 8449 50535 8483
rect 50818 8449 50852 8483
rect 51273 8449 51307 8483
rect 51366 8449 51400 8483
rect 51641 8449 51675 8483
rect 51738 8449 51772 8483
rect 53481 8449 53515 8483
rect 54953 8449 54987 8483
rect 78045 8449 78079 8483
rect 29193 8381 29227 8415
rect 33241 8381 33275 8415
rect 40785 8381 40819 8415
rect 40877 8381 40911 8415
rect 43729 8381 43763 8415
rect 47133 8381 47167 8415
rect 47409 8381 47443 8415
rect 49065 8381 49099 8415
rect 50261 8381 50295 8415
rect 53757 8381 53791 8415
rect 54401 8381 54435 8415
rect 30665 8313 30699 8347
rect 35725 8313 35759 8347
rect 36829 8313 36863 8347
rect 37749 8313 37783 8347
rect 40969 8313 41003 8347
rect 43269 8313 43303 8347
rect 52009 8313 52043 8347
rect 53021 8313 53055 8347
rect 53665 8313 53699 8347
rect 78229 8313 78263 8347
rect 30849 8245 30883 8279
rect 37289 8245 37323 8279
rect 40417 8245 40451 8279
rect 43637 8245 43671 8279
rect 44557 8245 44591 8279
rect 45293 8245 45327 8279
rect 48605 8245 48639 8279
rect 51917 8245 51951 8279
rect 53297 8245 53331 8279
rect 30205 8041 30239 8075
rect 35449 8041 35483 8075
rect 35633 8041 35667 8075
rect 41613 8041 41647 8075
rect 42625 8041 42659 8075
rect 42809 8041 42843 8075
rect 43361 8041 43395 8075
rect 44557 8041 44591 8075
rect 45937 8041 45971 8075
rect 47317 8041 47351 8075
rect 49985 8041 50019 8075
rect 52929 8041 52963 8075
rect 54861 8041 54895 8075
rect 78045 8041 78079 8075
rect 36093 7973 36127 8007
rect 36553 7973 36587 8007
rect 45017 7973 45051 8007
rect 55045 7973 55079 8007
rect 77769 7973 77803 8007
rect 31401 7905 31435 7939
rect 35909 7905 35943 7939
rect 37657 7905 37691 7939
rect 38485 7905 38519 7939
rect 39865 7905 39899 7939
rect 40141 7905 40175 7939
rect 42901 7905 42935 7939
rect 46029 7905 46063 7939
rect 46857 7905 46891 7939
rect 48237 7905 48271 7939
rect 48513 7905 48547 7939
rect 50261 7905 50295 7939
rect 51181 7905 51215 7939
rect 53113 7905 53147 7939
rect 30389 7837 30423 7871
rect 30573 7837 30607 7871
rect 30665 7837 30699 7871
rect 30757 7837 30791 7871
rect 31677 7837 31711 7871
rect 31769 7837 31803 7871
rect 32045 7837 32079 7871
rect 34897 7837 34931 7871
rect 35265 7837 35299 7871
rect 38301 7837 38335 7871
rect 38393 7837 38427 7871
rect 38669 7837 38703 7871
rect 38761 7837 38795 7871
rect 39221 7837 39255 7871
rect 39313 7837 39347 7871
rect 42073 7837 42107 7871
rect 42257 7837 42291 7871
rect 42441 7837 42475 7871
rect 45385 7837 45419 7871
rect 45661 7837 45695 7871
rect 45753 7837 45787 7871
rect 46673 7837 46707 7871
rect 46765 7837 46799 7871
rect 47041 7837 47075 7871
rect 47133 7837 47167 7871
rect 47593 7837 47627 7871
rect 47685 7837 47719 7871
rect 55505 7837 55539 7871
rect 55689 7837 55723 7871
rect 55873 7837 55907 7871
rect 77585 7837 77619 7871
rect 77861 7837 77895 7871
rect 78229 7837 78263 7871
rect 31861 7769 31895 7803
rect 35081 7769 35115 7803
rect 35173 7769 35207 7803
rect 39037 7769 39071 7803
rect 42349 7769 42383 7803
rect 45569 7769 45603 7803
rect 47409 7769 47443 7803
rect 51457 7769 51491 7803
rect 53389 7769 53423 7803
rect 55597 7769 55631 7803
rect 31493 7701 31527 7735
rect 36277 7701 36311 7735
rect 38945 7701 38979 7735
rect 50353 7701 50387 7735
rect 55321 7701 55355 7735
rect 77309 7701 77343 7735
rect 77401 7701 77435 7735
rect 78413 7701 78447 7735
rect 31769 7497 31803 7531
rect 37289 7497 37323 7531
rect 43269 7497 43303 7531
rect 44005 7497 44039 7531
rect 51549 7497 51583 7531
rect 53481 7497 53515 7531
rect 42717 7429 42751 7463
rect 49985 7429 50019 7463
rect 50077 7429 50111 7463
rect 54953 7429 54987 7463
rect 55321 7429 55355 7463
rect 30941 7361 30975 7395
rect 31033 7361 31067 7395
rect 31309 7361 31343 7395
rect 32137 7361 32171 7395
rect 32781 7361 32815 7395
rect 33701 7361 33735 7395
rect 33885 7361 33919 7395
rect 39037 7361 39071 7395
rect 42441 7361 42475 7395
rect 42625 7361 42659 7395
rect 42809 7361 42843 7395
rect 43453 7361 43487 7395
rect 43637 7361 43671 7395
rect 43729 7361 43763 7395
rect 43821 7361 43855 7395
rect 44189 7361 44223 7395
rect 49893 7361 49927 7395
rect 50261 7361 50295 7395
rect 51733 7361 51767 7395
rect 53297 7361 53331 7395
rect 53660 7361 53694 7395
rect 53757 7361 53791 7395
rect 53849 7361 53883 7395
rect 53977 7361 54011 7395
rect 54125 7361 54159 7395
rect 54401 7361 54435 7395
rect 54677 7361 54711 7395
rect 54769 7361 54803 7395
rect 77769 7361 77803 7395
rect 78045 7361 78079 7395
rect 31217 7293 31251 7327
rect 32965 7293 32999 7327
rect 33517 7293 33551 7327
rect 33609 7293 33643 7327
rect 38761 7293 38795 7327
rect 52009 7293 52043 7327
rect 52745 7293 52779 7327
rect 55045 7293 55079 7327
rect 56793 7293 56827 7327
rect 77953 7225 77987 7259
rect 30757 7157 30791 7191
rect 34069 7157 34103 7191
rect 42993 7157 43027 7191
rect 49709 7157 49743 7191
rect 51917 7157 51951 7191
rect 54493 7157 54527 7191
rect 56885 7157 56919 7191
rect 77677 7157 77711 7191
rect 78229 7157 78263 7191
rect 30100 6953 30134 6987
rect 32229 6953 32263 6987
rect 34081 6953 34115 6987
rect 46213 6953 46247 6987
rect 47225 6953 47259 6987
rect 53297 6953 53331 6987
rect 41061 6885 41095 6919
rect 29837 6817 29871 6851
rect 31585 6817 31619 6851
rect 32505 6817 32539 6851
rect 35449 6817 35483 6851
rect 41981 6817 42015 6851
rect 42533 6817 42567 6851
rect 44741 6817 44775 6851
rect 45017 6817 45051 6851
rect 49801 6817 49835 6851
rect 31677 6749 31711 6783
rect 32045 6749 32079 6783
rect 34345 6749 34379 6783
rect 35265 6749 35299 6783
rect 35541 6749 35575 6783
rect 36093 6749 36127 6783
rect 36645 6749 36679 6783
rect 37013 6749 37047 6783
rect 37381 6749 37415 6783
rect 38296 6749 38330 6783
rect 38485 6749 38519 6783
rect 38668 6749 38702 6783
rect 38761 6749 38795 6783
rect 40509 6749 40543 6783
rect 40877 6749 40911 6783
rect 41245 6749 41279 6783
rect 41797 6749 41831 6783
rect 41889 6749 41923 6783
rect 42165 6749 42199 6783
rect 42257 6749 42291 6783
rect 42993 6749 43027 6783
rect 46397 6749 46431 6783
rect 46490 6749 46524 6783
rect 46862 6749 46896 6783
rect 47133 6749 47167 6783
rect 47409 6749 47443 6783
rect 49525 6749 49559 6783
rect 49617 6749 49651 6783
rect 49893 6749 49927 6783
rect 77769 6749 77803 6783
rect 77861 6749 77895 6783
rect 37105 6681 37139 6715
rect 37197 6681 37231 6715
rect 37565 6681 37599 6715
rect 38393 6681 38427 6715
rect 40693 6681 40727 6715
rect 40785 6681 40819 6715
rect 43269 6681 43303 6715
rect 46673 6681 46707 6715
rect 46765 6681 46799 6715
rect 31861 6613 31895 6647
rect 32597 6613 32631 6647
rect 35081 6613 35115 6647
rect 36829 6613 36863 6647
rect 37657 6613 37691 6647
rect 38117 6613 38151 6647
rect 42441 6613 42475 6647
rect 47041 6613 47075 6647
rect 47593 6613 47627 6647
rect 49341 6613 49375 6647
rect 78045 6613 78079 6647
rect 30113 6409 30147 6443
rect 33701 6409 33735 6443
rect 36553 6409 36587 6443
rect 40141 6409 40175 6443
rect 42809 6409 42843 6443
rect 42993 6409 43027 6443
rect 44281 6409 44315 6443
rect 45109 6409 45143 6443
rect 47593 6409 47627 6443
rect 51181 6409 51215 6443
rect 54953 6409 54987 6443
rect 30297 6341 30331 6375
rect 31585 6341 31619 6375
rect 31677 6341 31711 6375
rect 33425 6341 33459 6375
rect 35081 6341 35115 6375
rect 41613 6341 41647 6375
rect 44741 6341 44775 6375
rect 44833 6341 44867 6375
rect 45201 6341 45235 6375
rect 49065 6341 49099 6375
rect 49709 6341 49743 6375
rect 31493 6273 31527 6307
rect 31861 6273 31895 6307
rect 33057 6273 33091 6307
rect 33205 6273 33239 6307
rect 33333 6273 33367 6307
rect 33522 6273 33556 6307
rect 34805 6273 34839 6307
rect 38485 6273 38519 6307
rect 43177 6273 43211 6307
rect 43269 6273 43303 6307
rect 43545 6273 43579 6307
rect 44465 6273 44499 6307
rect 44613 6273 44647 6307
rect 44971 6273 45005 6307
rect 46489 6273 46523 6307
rect 53757 6273 53791 6307
rect 53849 6273 53883 6307
rect 53941 6273 53975 6307
rect 54125 6273 54159 6307
rect 54769 6273 54803 6307
rect 78045 6273 78079 6307
rect 31033 6205 31067 6239
rect 38761 6205 38795 6239
rect 39221 6205 39255 6239
rect 39773 6205 39807 6239
rect 41889 6205 41923 6239
rect 45937 6205 45971 6239
rect 46213 6205 46247 6239
rect 49341 6205 49375 6239
rect 49433 6205 49467 6239
rect 53389 6205 53423 6239
rect 38669 6137 38703 6171
rect 78229 6137 78263 6171
rect 31309 6069 31343 6103
rect 38301 6069 38335 6103
rect 43453 6069 43487 6103
rect 46305 6069 46339 6103
rect 46673 6069 46707 6103
rect 52837 6069 52871 6103
rect 53573 6069 53607 6103
rect 54217 6069 54251 6103
rect 55229 6069 55263 6103
rect 32229 5865 32263 5899
rect 35357 5865 35391 5899
rect 39589 5865 39623 5899
rect 45017 5865 45051 5899
rect 49893 5865 49927 5899
rect 53297 5865 53331 5899
rect 32137 5797 32171 5831
rect 78045 5797 78079 5831
rect 30389 5729 30423 5763
rect 37841 5729 37875 5763
rect 38117 5729 38151 5763
rect 46489 5729 46523 5763
rect 46765 5729 46799 5763
rect 55137 5729 55171 5763
rect 33655 5661 33689 5695
rect 33793 5661 33827 5695
rect 34068 5661 34102 5695
rect 34161 5661 34195 5695
rect 34713 5661 34747 5695
rect 34806 5661 34840 5695
rect 35178 5661 35212 5695
rect 36645 5661 36679 5695
rect 36793 5661 36827 5695
rect 36921 5661 36955 5695
rect 37151 5661 37185 5695
rect 41608 5661 41642 5695
rect 41705 5661 41739 5695
rect 41797 5661 41831 5695
rect 41925 5661 41959 5695
rect 42073 5661 42107 5695
rect 49709 5661 49743 5695
rect 50348 5661 50382 5695
rect 50445 5661 50479 5695
rect 50720 5661 50754 5695
rect 50813 5661 50847 5695
rect 50925 5661 50959 5695
rect 51181 5661 51215 5695
rect 51273 5661 51307 5695
rect 51549 5661 51583 5695
rect 53389 5661 53423 5695
rect 77861 5661 77895 5695
rect 78229 5661 78263 5695
rect 30665 5593 30699 5627
rect 33885 5593 33919 5627
rect 34989 5593 35023 5627
rect 35081 5593 35115 5627
rect 37013 5593 37047 5627
rect 50537 5593 50571 5627
rect 51089 5593 51123 5627
rect 51825 5593 51859 5627
rect 53665 5593 53699 5627
rect 55413 5593 55447 5627
rect 55873 5593 55907 5627
rect 33517 5525 33551 5559
rect 37289 5525 37323 5559
rect 41429 5525 41463 5559
rect 49341 5525 49375 5559
rect 49525 5525 49559 5559
rect 50169 5525 50203 5559
rect 51457 5525 51491 5559
rect 55505 5525 55539 5559
rect 56149 5525 56183 5559
rect 77677 5525 77711 5559
rect 78413 5525 78447 5559
rect 30941 5321 30975 5355
rect 36829 5321 36863 5355
rect 43545 5321 43579 5355
rect 44005 5321 44039 5355
rect 53113 5321 53147 5355
rect 34989 5253 35023 5287
rect 42901 5253 42935 5287
rect 42993 5253 43027 5287
rect 53297 5253 53331 5287
rect 31125 5185 31159 5219
rect 31217 5185 31251 5219
rect 31493 5185 31527 5219
rect 33149 5185 33183 5219
rect 33333 5185 33367 5219
rect 34345 5185 34379 5219
rect 34713 5185 34747 5219
rect 34897 5185 34931 5219
rect 35081 5185 35115 5219
rect 36277 5185 36311 5219
rect 36369 5185 36403 5219
rect 36461 5185 36495 5219
rect 36645 5185 36679 5219
rect 37013 5185 37047 5219
rect 37473 5185 37507 5219
rect 38853 5185 38887 5219
rect 42763 5185 42797 5219
rect 43121 5185 43155 5219
rect 43269 5185 43303 5219
rect 43453 5185 43487 5219
rect 44097 5185 44131 5219
rect 49709 5185 49743 5219
rect 50721 5185 50755 5219
rect 51917 5185 51951 5219
rect 52009 5185 52043 5219
rect 52285 5185 52319 5219
rect 54677 5185 54711 5219
rect 55137 5185 55171 5219
rect 78045 5185 78079 5219
rect 78321 5185 78355 5219
rect 31401 5117 31435 5151
rect 33425 5117 33459 5151
rect 33701 5117 33735 5151
rect 37749 5117 37783 5151
rect 38301 5117 38335 5151
rect 49893 5117 49927 5151
rect 49985 5117 50019 5151
rect 50077 5117 50111 5151
rect 51733 5117 51767 5151
rect 54125 5117 54159 5151
rect 36001 5049 36035 5083
rect 54861 5049 54895 5083
rect 32965 4981 32999 5015
rect 35265 4981 35299 5015
rect 36093 4981 36127 5015
rect 37289 4981 37323 5015
rect 37657 4981 37691 5015
rect 42625 4981 42659 5015
rect 49525 4981 49559 5015
rect 52193 4981 52227 5015
rect 78137 4981 78171 5015
rect 29929 4777 29963 4811
rect 44557 4777 44591 4811
rect 47409 4777 47443 4811
rect 51653 4777 51687 4811
rect 53389 4777 53423 4811
rect 33793 4709 33827 4743
rect 38669 4709 38703 4743
rect 41613 4709 41647 4743
rect 47225 4709 47259 4743
rect 53849 4709 53883 4743
rect 32045 4641 32079 4675
rect 32321 4641 32355 4675
rect 35725 4641 35759 4675
rect 37197 4641 37231 4675
rect 41705 4641 41739 4675
rect 42257 4641 42291 4675
rect 50169 4641 50203 4675
rect 51917 4641 51951 4675
rect 30021 4573 30055 4607
rect 30205 4573 30239 4607
rect 35449 4573 35483 4607
rect 35541 4573 35575 4607
rect 35817 4573 35851 4607
rect 36921 4573 36955 4607
rect 39865 4573 39899 4607
rect 42809 4573 42843 4607
rect 45017 4573 45051 4607
rect 45201 4573 45235 4607
rect 45385 4573 45419 4607
rect 46673 4573 46707 4607
rect 47041 4573 47075 4607
rect 47317 4573 47351 4607
rect 47593 4573 47627 4607
rect 47685 4573 47719 4607
rect 53573 4573 53607 4607
rect 53665 4573 53699 4607
rect 53941 4573 53975 4607
rect 78229 4573 78263 4607
rect 78505 4573 78539 4607
rect 35909 4505 35943 4539
rect 36645 4505 36679 4539
rect 40141 4505 40175 4539
rect 43085 4505 43119 4539
rect 45293 4505 45327 4539
rect 46857 4505 46891 4539
rect 46949 4505 46983 4539
rect 30113 4437 30147 4471
rect 35265 4437 35299 4471
rect 45569 4437 45603 4471
rect 47869 4437 47903 4471
rect 78321 4437 78355 4471
rect 36921 4233 36955 4267
rect 40509 4233 40543 4267
rect 43361 4233 43395 4267
rect 47593 4233 47627 4267
rect 41981 4165 42015 4199
rect 31493 4097 31527 4131
rect 36093 4097 36127 4131
rect 36369 4097 36403 4131
rect 36461 4097 36495 4131
rect 36737 4097 36771 4131
rect 37289 4097 37323 4131
rect 40693 4097 40727 4131
rect 41245 4097 41279 4131
rect 41337 4097 41371 4131
rect 41613 4097 41647 4131
rect 41889 4097 41923 4131
rect 42073 4097 42107 4131
rect 42257 4097 42291 4131
rect 43177 4097 43211 4131
rect 43545 4097 43579 4131
rect 44741 4097 44775 4131
rect 45293 4097 45327 4131
rect 45385 4097 45419 4131
rect 45661 4097 45695 4131
rect 58449 4097 58483 4131
rect 58633 4097 58667 4131
rect 34345 4029 34379 4063
rect 35817 4029 35851 4063
rect 37841 4029 37875 4063
rect 40969 4029 41003 4063
rect 42625 4029 42659 4063
rect 43821 4029 43855 4063
rect 44097 4029 44131 4063
rect 49065 4029 49099 4063
rect 49341 4029 49375 4063
rect 36645 3961 36679 3995
rect 40877 3961 40911 3995
rect 41705 3961 41739 3995
rect 43729 3961 43763 3995
rect 45569 3961 45603 3995
rect 58265 3961 58299 3995
rect 31677 3893 31711 3927
rect 31953 3893 31987 3927
rect 36185 3893 36219 3927
rect 41061 3893 41095 3927
rect 41521 3893 41555 3927
rect 45109 3893 45143 3927
rect 56425 3893 56459 3927
rect 30021 3689 30055 3723
rect 46765 3689 46799 3723
rect 50353 3689 50387 3723
rect 50997 3689 51031 3723
rect 57161 3689 57195 3723
rect 59369 3689 59403 3723
rect 72617 3689 72651 3723
rect 32321 3621 32355 3655
rect 32597 3621 32631 3655
rect 38669 3621 38703 3655
rect 42901 3621 42935 3655
rect 44649 3621 44683 3655
rect 56149 3621 56183 3655
rect 58909 3621 58943 3655
rect 30205 3553 30239 3587
rect 30481 3553 30515 3587
rect 41153 3553 41187 3587
rect 45017 3553 45051 3587
rect 45293 3553 45327 3587
rect 59093 3553 59127 3587
rect 72525 3553 72559 3587
rect 32137 3485 32171 3519
rect 44281 3485 44315 3519
rect 50629 3485 50663 3519
rect 51273 3485 51307 3519
rect 55321 3485 55355 3519
rect 56333 3485 56367 3519
rect 56517 3485 56551 3519
rect 56609 3485 56643 3519
rect 57529 3485 57563 3519
rect 57621 3485 57655 3519
rect 58173 3485 58207 3519
rect 58541 3485 58575 3519
rect 59001 3485 59035 3519
rect 72341 3485 72375 3519
rect 72709 3485 72743 3519
rect 72985 3485 73019 3519
rect 38945 3417 38979 3451
rect 41429 3417 41463 3451
rect 43637 3417 43671 3451
rect 43821 3417 43855 3451
rect 44465 3417 44499 3451
rect 51181 3417 51215 3451
rect 55965 3417 55999 3451
rect 58633 3417 58667 3451
rect 59553 3417 59587 3451
rect 72617 3417 72651 3451
rect 31953 3349 31987 3383
rect 50813 3349 50847 3383
rect 50981 3349 51015 3383
rect 56793 3349 56827 3383
rect 56977 3349 57011 3383
rect 57161 3349 57195 3383
rect 58357 3349 58391 3383
rect 58725 3349 58759 3383
rect 72157 3349 72191 3383
rect 72893 3349 72927 3383
rect 78045 3349 78079 3383
rect 78505 3349 78539 3383
rect 31861 3145 31895 3179
rect 45109 3145 45143 3179
rect 54309 3145 54343 3179
rect 57897 3145 57931 3179
rect 58265 3145 58299 3179
rect 59369 3145 59403 3179
rect 66177 3145 66211 3179
rect 68385 3145 68419 3179
rect 68937 3145 68971 3179
rect 72525 3145 72559 3179
rect 72617 3145 72651 3179
rect 73537 3145 73571 3179
rect 78137 3145 78171 3179
rect 45017 3077 45051 3111
rect 50822 3077 50856 3111
rect 53665 3077 53699 3111
rect 53849 3077 53883 3111
rect 54033 3077 54067 3111
rect 55781 3077 55815 3111
rect 59921 3077 59955 3111
rect 66637 3077 66671 3111
rect 69121 3077 69155 3111
rect 71053 3077 71087 3111
rect 72065 3077 72099 3111
rect 73445 3077 73479 3111
rect 74273 3077 74307 3111
rect 74365 3077 74399 3111
rect 32321 3009 32355 3043
rect 35357 3009 35391 3043
rect 37933 3009 37967 3043
rect 38200 3009 38234 3043
rect 39405 3009 39439 3043
rect 39957 3009 39991 3043
rect 40213 3009 40247 3043
rect 44566 3009 44600 3043
rect 44833 3009 44867 3043
rect 45569 3009 45603 3043
rect 46213 3009 46247 3043
rect 46857 3009 46891 3043
rect 47593 3009 47627 3043
rect 48789 3009 48823 3043
rect 49433 3009 49467 3043
rect 51089 3009 51123 3043
rect 51365 3009 51399 3043
rect 51457 3009 51491 3043
rect 56149 3009 56183 3043
rect 56425 3009 56459 3043
rect 56701 3009 56735 3043
rect 57713 3009 57747 3043
rect 58725 3009 58759 3043
rect 59001 3009 59035 3043
rect 59553 3009 59587 3043
rect 59829 3009 59863 3043
rect 60197 3009 60231 3043
rect 61577 3009 61611 3043
rect 61945 3009 61979 3043
rect 62221 3009 62255 3043
rect 62589 3009 62623 3043
rect 63049 3009 63083 3043
rect 63417 3009 63451 3043
rect 63509 3009 63543 3043
rect 63877 3009 63911 3043
rect 64153 3009 64187 3043
rect 64521 3009 64555 3043
rect 66361 3009 66395 3043
rect 68201 3009 68235 3043
rect 68753 3009 68787 3043
rect 70961 3009 70995 3043
rect 71145 3009 71179 3043
rect 72341 3009 72375 3043
rect 72801 3009 72835 3043
rect 73077 3009 73111 3043
rect 74089 3009 74123 3043
rect 74181 3009 74215 3043
rect 76205 3009 76239 3043
rect 76389 3009 76423 3043
rect 77677 3009 77711 3043
rect 77853 3009 77887 3043
rect 78321 3009 78355 3043
rect 35633 2941 35667 2975
rect 37105 2941 37139 2975
rect 42073 2941 42107 2975
rect 56057 2941 56091 2975
rect 56241 2941 56275 2975
rect 58357 2941 58391 2975
rect 58449 2941 58483 2975
rect 58817 2941 58851 2975
rect 59737 2941 59771 2975
rect 60013 2941 60047 2975
rect 66545 2941 66579 2975
rect 72249 2941 72283 2975
rect 72985 2941 73019 2975
rect 74549 2941 74583 2975
rect 39313 2873 39347 2907
rect 41337 2873 41371 2907
rect 49617 2873 49651 2907
rect 59185 2873 59219 2907
rect 60381 2873 60415 2907
rect 32505 2805 32539 2839
rect 39589 2805 39623 2839
rect 41429 2805 41463 2839
rect 43361 2805 43395 2839
rect 43453 2805 43487 2839
rect 45753 2805 45787 2839
rect 46397 2805 46431 2839
rect 47041 2805 47075 2839
rect 47777 2805 47811 2839
rect 48973 2805 49007 2839
rect 49709 2805 49743 2839
rect 51181 2805 51215 2839
rect 51641 2805 51675 2839
rect 53481 2805 53515 2839
rect 54125 2805 54159 2839
rect 56609 2805 56643 2839
rect 57437 2805 57471 2839
rect 58725 2805 58759 2839
rect 59553 2805 59587 2839
rect 59921 2805 59955 2839
rect 61761 2805 61795 2839
rect 62405 2805 62439 2839
rect 63233 2805 63267 2839
rect 63693 2805 63727 2839
rect 64337 2805 64371 2839
rect 65993 2805 66027 2839
rect 66637 2805 66671 2839
rect 68569 2805 68603 2839
rect 72341 2805 72375 2839
rect 73077 2805 73111 2839
rect 76573 2805 76607 2839
rect 78045 2805 78079 2839
rect 38669 2601 38703 2635
rect 39957 2601 39991 2635
rect 43729 2601 43763 2635
rect 50537 2601 50571 2635
rect 54125 2601 54159 2635
rect 54585 2601 54619 2635
rect 58449 2601 58483 2635
rect 60013 2601 60047 2635
rect 66637 2601 66671 2635
rect 69673 2601 69707 2635
rect 70317 2601 70351 2635
rect 71605 2601 71639 2635
rect 72249 2601 72283 2635
rect 72433 2601 72467 2635
rect 73537 2601 73571 2635
rect 74181 2601 74215 2635
rect 75469 2601 75503 2635
rect 76113 2601 76147 2635
rect 77401 2601 77435 2635
rect 77769 2601 77803 2635
rect 44649 2533 44683 2567
rect 50813 2533 50847 2567
rect 53113 2533 53147 2567
rect 54401 2533 54435 2567
rect 55413 2533 55447 2567
rect 58081 2533 58115 2567
rect 60657 2533 60691 2567
rect 61301 2533 61335 2567
rect 67281 2533 67315 2567
rect 67925 2533 67959 2567
rect 69213 2533 69247 2567
rect 74825 2533 74859 2567
rect 39497 2465 39531 2499
rect 44373 2465 44407 2499
rect 46857 2465 46891 2499
rect 54677 2465 54711 2499
rect 55689 2465 55723 2499
rect 72617 2465 72651 2499
rect 32965 2397 32999 2431
rect 38025 2397 38059 2431
rect 38209 2397 38243 2431
rect 38301 2397 38335 2431
rect 38393 2397 38427 2431
rect 38945 2397 38979 2431
rect 40141 2397 40175 2431
rect 40417 2397 40451 2431
rect 40601 2397 40635 2431
rect 42901 2397 42935 2431
rect 43085 2397 43119 2431
rect 43269 2397 43303 2431
rect 43361 2397 43395 2431
rect 43453 2397 43487 2431
rect 43821 2397 43855 2431
rect 44833 2397 44867 2431
rect 45017 2397 45051 2431
rect 45385 2397 45419 2431
rect 45661 2397 45695 2431
rect 45845 2397 45879 2431
rect 46213 2397 46247 2431
rect 46489 2397 46523 2431
rect 47133 2397 47167 2431
rect 47777 2397 47811 2431
rect 48697 2397 48731 2431
rect 49065 2397 49099 2431
rect 49709 2397 49743 2431
rect 50353 2397 50387 2431
rect 50629 2397 50663 2431
rect 51273 2397 51307 2431
rect 51641 2397 51675 2431
rect 52285 2397 52319 2431
rect 52929 2397 52963 2431
rect 53573 2397 53607 2431
rect 53941 2397 53975 2431
rect 54217 2397 54251 2431
rect 54585 2397 54619 2431
rect 54861 2397 54895 2431
rect 55321 2397 55355 2431
rect 57529 2397 57563 2431
rect 57897 2397 57931 2431
rect 58265 2397 58299 2431
rect 58541 2397 58575 2431
rect 58909 2397 58943 2431
rect 59553 2397 59587 2431
rect 60197 2397 60231 2431
rect 60841 2397 60875 2431
rect 61485 2397 61519 2431
rect 61945 2397 61979 2431
rect 62589 2397 62623 2431
rect 63233 2397 63267 2431
rect 63877 2397 63911 2431
rect 64521 2397 64555 2431
rect 65165 2397 65199 2431
rect 65809 2397 65843 2431
rect 66453 2397 66487 2431
rect 67097 2397 67131 2431
rect 67741 2397 67775 2431
rect 68661 2397 68695 2431
rect 69029 2397 69063 2431
rect 69857 2397 69891 2431
rect 70501 2397 70535 2431
rect 70961 2397 70995 2431
rect 71789 2397 71823 2431
rect 71973 2397 72007 2431
rect 72433 2397 72467 2431
rect 72709 2397 72743 2431
rect 72893 2397 72927 2431
rect 73721 2397 73755 2431
rect 74365 2397 74399 2431
rect 75009 2397 75043 2431
rect 75653 2397 75687 2431
rect 76297 2397 76331 2431
rect 76757 2397 76791 2431
rect 77585 2397 77619 2431
rect 77953 2397 77987 2431
rect 78045 2397 78079 2431
rect 38853 2329 38887 2363
rect 40785 2329 40819 2363
rect 49525 2329 49559 2363
rect 50169 2329 50203 2363
rect 51365 2329 51399 2363
rect 53389 2329 53423 2363
rect 55965 2329 55999 2363
rect 59001 2329 59035 2363
rect 73353 2329 73387 2363
rect 73813 2329 73847 2363
rect 33149 2261 33183 2295
rect 42717 2261 42751 2295
rect 45201 2261 45235 2295
rect 45569 2261 45603 2295
rect 46029 2261 46063 2295
rect 46397 2261 46431 2295
rect 46673 2261 46707 2295
rect 47317 2261 47351 2295
rect 47961 2261 47995 2295
rect 48513 2261 48547 2295
rect 49249 2261 49283 2295
rect 49893 2261 49927 2295
rect 51089 2261 51123 2295
rect 51825 2261 51859 2295
rect 52193 2261 52227 2295
rect 52469 2261 52503 2295
rect 52837 2261 52871 2295
rect 53757 2261 53791 2295
rect 55045 2261 55079 2295
rect 57437 2261 57471 2295
rect 57713 2261 57747 2295
rect 58725 2261 58759 2295
rect 59277 2261 59311 2295
rect 59369 2261 59403 2295
rect 59921 2261 59955 2295
rect 60565 2261 60599 2295
rect 61209 2261 61243 2295
rect 62129 2261 62163 2295
rect 62773 2261 62807 2295
rect 63417 2261 63451 2295
rect 64061 2261 64095 2295
rect 64705 2261 64739 2295
rect 65073 2261 65107 2295
rect 65349 2261 65383 2295
rect 65717 2261 65751 2295
rect 65993 2261 66027 2295
rect 66269 2261 66303 2295
rect 67005 2261 67039 2295
rect 67649 2261 67683 2295
rect 68477 2261 68511 2295
rect 68937 2261 68971 2295
rect 69581 2261 69615 2295
rect 70225 2261 70259 2295
rect 70869 2261 70903 2295
rect 71145 2261 71179 2295
rect 71513 2261 71547 2295
rect 72157 2261 72191 2295
rect 73077 2261 73111 2295
rect 74089 2261 74123 2295
rect 74733 2261 74767 2295
rect 75377 2261 75411 2295
rect 76021 2261 76055 2295
rect 76941 2261 76975 2295
rect 77309 2261 77343 2295
rect 78229 2261 78263 2295
<< metal1 >>
rect 1104 37562 78844 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 78844 37562
rect 1104 37488 78844 37510
rect 38654 37408 38660 37460
rect 38712 37448 38718 37460
rect 38841 37451 38899 37457
rect 38841 37448 38853 37451
rect 38712 37420 38853 37448
rect 38712 37408 38718 37420
rect 38841 37417 38853 37420
rect 38887 37417 38899 37451
rect 38841 37411 38899 37417
rect 45094 37408 45100 37460
rect 45152 37448 45158 37460
rect 45557 37451 45615 37457
rect 45557 37448 45569 37451
rect 45152 37420 45569 37448
rect 45152 37408 45158 37420
rect 45557 37417 45569 37420
rect 45603 37417 45615 37451
rect 45557 37411 45615 37417
rect 46382 37408 46388 37460
rect 46440 37448 46446 37460
rect 46661 37451 46719 37457
rect 46661 37448 46673 37451
rect 46440 37420 46673 37448
rect 46440 37408 46446 37420
rect 46661 37417 46673 37420
rect 46707 37417 46719 37451
rect 46661 37411 46719 37417
rect 43806 37340 43812 37392
rect 43864 37380 43870 37392
rect 44177 37383 44235 37389
rect 44177 37380 44189 37383
rect 43864 37352 44189 37380
rect 43864 37340 43870 37352
rect 44177 37349 44189 37352
rect 44223 37349 44235 37383
rect 44177 37343 44235 37349
rect 36262 37204 36268 37256
rect 36320 37204 36326 37256
rect 40494 37204 40500 37256
rect 40552 37204 40558 37256
rect 40773 37247 40831 37253
rect 40773 37213 40785 37247
rect 40819 37244 40831 37247
rect 40862 37244 40868 37256
rect 40819 37216 40868 37244
rect 40819 37213 40831 37216
rect 40773 37207 40831 37213
rect 40862 37204 40868 37216
rect 40920 37204 40926 37256
rect 39117 37179 39175 37185
rect 39117 37145 39129 37179
rect 39163 37176 39175 37179
rect 39390 37176 39396 37188
rect 39163 37148 39396 37176
rect 39163 37145 39175 37148
rect 39117 37139 39175 37145
rect 39390 37136 39396 37148
rect 39448 37136 39454 37188
rect 43898 37136 43904 37188
rect 43956 37176 43962 37188
rect 43993 37179 44051 37185
rect 43993 37176 44005 37179
rect 43956 37148 44005 37176
rect 43956 37136 43962 37148
rect 43993 37145 44005 37148
rect 44039 37145 44051 37179
rect 43993 37139 44051 37145
rect 44358 37136 44364 37188
rect 44416 37176 44422 37188
rect 45281 37179 45339 37185
rect 45281 37176 45293 37179
rect 44416 37148 45293 37176
rect 44416 37136 44422 37148
rect 45281 37145 45293 37148
rect 45327 37145 45339 37179
rect 45281 37139 45339 37145
rect 46106 37136 46112 37188
rect 46164 37176 46170 37188
rect 46569 37179 46627 37185
rect 46569 37176 46581 37179
rect 46164 37148 46581 37176
rect 46164 37136 46170 37148
rect 46569 37145 46581 37148
rect 46615 37145 46627 37179
rect 46569 37139 46627 37145
rect 35434 37068 35440 37120
rect 35492 37108 35498 37120
rect 35713 37111 35771 37117
rect 35713 37108 35725 37111
rect 35492 37080 35725 37108
rect 35492 37068 35498 37080
rect 35713 37077 35725 37080
rect 35759 37077 35771 37111
rect 35713 37071 35771 37077
rect 1104 37018 78844 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 66314 37018
rect 66366 36966 66378 37018
rect 66430 36966 66442 37018
rect 66494 36966 66506 37018
rect 66558 36966 66570 37018
rect 66622 36966 78844 37018
rect 1104 36944 78844 36966
rect 35621 36907 35679 36913
rect 35621 36873 35633 36907
rect 35667 36904 35679 36907
rect 36262 36904 36268 36916
rect 35667 36876 36268 36904
rect 35667 36873 35679 36876
rect 35621 36867 35679 36873
rect 36262 36864 36268 36876
rect 36320 36864 36326 36916
rect 39942 36864 39948 36916
rect 40000 36904 40006 36916
rect 40313 36907 40371 36913
rect 40313 36904 40325 36907
rect 40000 36876 40325 36904
rect 40000 36864 40006 36876
rect 40313 36873 40325 36876
rect 40359 36873 40371 36907
rect 40313 36867 40371 36873
rect 40586 36864 40592 36916
rect 40644 36904 40650 36916
rect 40681 36907 40739 36913
rect 40681 36904 40693 36907
rect 40644 36876 40693 36904
rect 40644 36864 40650 36876
rect 40681 36873 40693 36876
rect 40727 36873 40739 36907
rect 40681 36867 40739 36873
rect 41141 36907 41199 36913
rect 41141 36873 41153 36907
rect 41187 36904 41199 36907
rect 41230 36904 41236 36916
rect 41187 36876 41236 36904
rect 41187 36873 41199 36876
rect 41141 36867 41199 36873
rect 41230 36864 41236 36876
rect 41288 36864 41294 36916
rect 41785 36907 41843 36913
rect 41785 36873 41797 36907
rect 41831 36904 41843 36907
rect 41874 36904 41880 36916
rect 41831 36876 41880 36904
rect 41831 36873 41843 36876
rect 41785 36867 41843 36873
rect 41874 36864 41880 36876
rect 41932 36864 41938 36916
rect 42518 36864 42524 36916
rect 42576 36904 42582 36916
rect 42613 36907 42671 36913
rect 42613 36904 42625 36907
rect 42576 36876 42625 36904
rect 42576 36864 42582 36876
rect 42613 36873 42625 36876
rect 42659 36873 42671 36907
rect 42613 36867 42671 36873
rect 42889 36907 42947 36913
rect 42889 36873 42901 36907
rect 42935 36904 42947 36907
rect 43162 36904 43168 36916
rect 42935 36876 43168 36904
rect 42935 36873 42947 36876
rect 42889 36867 42947 36873
rect 43162 36864 43168 36876
rect 43220 36864 43226 36916
rect 44450 36864 44456 36916
rect 44508 36904 44514 36916
rect 45189 36907 45247 36913
rect 45189 36904 45201 36907
rect 44508 36876 45201 36904
rect 44508 36864 44514 36876
rect 45189 36873 45201 36876
rect 45235 36873 45247 36907
rect 45189 36867 45247 36873
rect 45649 36907 45707 36913
rect 45649 36873 45661 36907
rect 45695 36904 45707 36907
rect 45738 36904 45744 36916
rect 45695 36876 45744 36904
rect 45695 36873 45707 36876
rect 45649 36867 45707 36873
rect 45738 36864 45744 36876
rect 45796 36864 45802 36916
rect 46106 36864 46112 36916
rect 46164 36864 46170 36916
rect 46937 36907 46995 36913
rect 46937 36873 46949 36907
rect 46983 36904 46995 36907
rect 47026 36904 47032 36916
rect 46983 36876 47032 36904
rect 46983 36873 46995 36876
rect 46937 36867 46995 36873
rect 47026 36864 47032 36876
rect 47084 36864 47090 36916
rect 47670 36864 47676 36916
rect 47728 36864 47734 36916
rect 48225 36907 48283 36913
rect 48225 36873 48237 36907
rect 48271 36904 48283 36907
rect 48314 36904 48320 36916
rect 48271 36876 48320 36904
rect 48271 36873 48283 36876
rect 48225 36867 48283 36873
rect 48314 36864 48320 36876
rect 48372 36864 48378 36916
rect 48958 36864 48964 36916
rect 49016 36864 49022 36916
rect 49421 36907 49479 36913
rect 49421 36873 49433 36907
rect 49467 36904 49479 36907
rect 49602 36904 49608 36916
rect 49467 36876 49608 36904
rect 49467 36873 49479 36876
rect 49421 36867 49479 36873
rect 49602 36864 49608 36876
rect 49660 36864 49666 36916
rect 50157 36907 50215 36913
rect 50157 36873 50169 36907
rect 50203 36904 50215 36907
rect 50246 36904 50252 36916
rect 50203 36876 50252 36904
rect 50203 36873 50215 36876
rect 50157 36867 50215 36873
rect 50246 36864 50252 36876
rect 50304 36864 50310 36916
rect 50801 36907 50859 36913
rect 50801 36873 50813 36907
rect 50847 36904 50859 36907
rect 50890 36904 50896 36916
rect 50847 36876 50896 36904
rect 50847 36873 50859 36876
rect 50801 36867 50859 36873
rect 50890 36864 50896 36876
rect 50948 36864 50954 36916
rect 51445 36907 51503 36913
rect 51445 36873 51457 36907
rect 51491 36904 51503 36907
rect 51534 36904 51540 36916
rect 51491 36876 51540 36904
rect 51491 36873 51503 36876
rect 51445 36867 51503 36873
rect 51534 36864 51540 36876
rect 51592 36864 51598 36916
rect 52089 36907 52147 36913
rect 52089 36873 52101 36907
rect 52135 36904 52147 36907
rect 52178 36904 52184 36916
rect 52135 36876 52184 36904
rect 52135 36873 52147 36876
rect 52089 36867 52147 36873
rect 52178 36864 52184 36876
rect 52236 36864 52242 36916
rect 52822 36864 52828 36916
rect 52880 36864 52886 36916
rect 53466 36864 53472 36916
rect 53524 36864 53530 36916
rect 53929 36907 53987 36913
rect 53929 36873 53941 36907
rect 53975 36904 53987 36907
rect 54110 36904 54116 36916
rect 53975 36876 54116 36904
rect 53975 36873 53987 36876
rect 53929 36867 53987 36873
rect 54110 36864 54116 36876
rect 54168 36864 54174 36916
rect 54573 36907 54631 36913
rect 54573 36873 54585 36907
rect 54619 36904 54631 36907
rect 54754 36904 54760 36916
rect 54619 36876 54760 36904
rect 54619 36873 54631 36876
rect 54573 36867 54631 36873
rect 54754 36864 54760 36876
rect 54812 36864 54818 36916
rect 55217 36907 55275 36913
rect 55217 36873 55229 36907
rect 55263 36904 55275 36907
rect 55398 36904 55404 36916
rect 55263 36876 55404 36904
rect 55263 36873 55275 36876
rect 55217 36867 55275 36873
rect 55398 36864 55404 36876
rect 55456 36864 55462 36916
rect 55861 36907 55919 36913
rect 55861 36873 55873 36907
rect 55907 36904 55919 36907
rect 56042 36904 56048 36916
rect 55907 36876 56048 36904
rect 55907 36873 55919 36876
rect 55861 36867 55919 36873
rect 56042 36864 56048 36876
rect 56100 36864 56106 36916
rect 56597 36907 56655 36913
rect 56597 36873 56609 36907
rect 56643 36904 56655 36907
rect 56686 36904 56692 36916
rect 56643 36876 56692 36904
rect 56643 36873 56655 36876
rect 56597 36867 56655 36873
rect 56686 36864 56692 36876
rect 56744 36864 56750 36916
rect 57241 36907 57299 36913
rect 57241 36873 57253 36907
rect 57287 36904 57299 36907
rect 57330 36904 57336 36916
rect 57287 36876 57336 36904
rect 57287 36873 57299 36876
rect 57241 36867 57299 36873
rect 57330 36864 57336 36876
rect 57388 36864 57394 36916
rect 57974 36864 57980 36916
rect 58032 36864 58038 36916
rect 58529 36907 58587 36913
rect 58529 36873 58541 36907
rect 58575 36904 58587 36907
rect 58618 36904 58624 36916
rect 58575 36876 58624 36904
rect 58575 36873 58587 36876
rect 58529 36867 58587 36873
rect 58618 36864 58624 36876
rect 58676 36864 58682 36916
rect 59173 36907 59231 36913
rect 59173 36873 59185 36907
rect 59219 36904 59231 36907
rect 59262 36904 59268 36916
rect 59219 36876 59268 36904
rect 59219 36873 59231 36876
rect 59173 36867 59231 36873
rect 59262 36864 59268 36876
rect 59320 36864 59326 36916
rect 59906 36864 59912 36916
rect 59964 36864 59970 36916
rect 60461 36907 60519 36913
rect 60461 36873 60473 36907
rect 60507 36904 60519 36907
rect 60550 36904 60556 36916
rect 60507 36876 60556 36904
rect 60507 36873 60519 36876
rect 60461 36867 60519 36873
rect 60550 36864 60556 36876
rect 60608 36864 60614 36916
rect 61194 36864 61200 36916
rect 61252 36864 61258 36916
rect 61657 36907 61715 36913
rect 61657 36873 61669 36907
rect 61703 36904 61715 36907
rect 61838 36904 61844 36916
rect 61703 36876 61844 36904
rect 61703 36873 61715 36876
rect 61657 36867 61715 36873
rect 61838 36864 61844 36876
rect 61896 36864 61902 36916
rect 62393 36907 62451 36913
rect 62393 36873 62405 36907
rect 62439 36904 62451 36907
rect 62482 36904 62488 36916
rect 62439 36876 62488 36904
rect 62439 36873 62451 36876
rect 62393 36867 62451 36873
rect 62482 36864 62488 36876
rect 62540 36864 62546 36916
rect 63126 36864 63132 36916
rect 63184 36904 63190 36916
rect 63221 36907 63279 36913
rect 63221 36904 63233 36907
rect 63184 36876 63233 36904
rect 63184 36864 63190 36876
rect 63221 36873 63233 36876
rect 63267 36873 63279 36907
rect 63221 36867 63279 36873
rect 63681 36907 63739 36913
rect 63681 36873 63693 36907
rect 63727 36904 63739 36907
rect 63770 36904 63776 36916
rect 63727 36876 63776 36904
rect 63727 36873 63739 36876
rect 63681 36867 63739 36873
rect 63770 36864 63776 36876
rect 63828 36864 63834 36916
rect 64325 36907 64383 36913
rect 64325 36873 64337 36907
rect 64371 36904 64383 36907
rect 64414 36904 64420 36916
rect 64371 36876 64420 36904
rect 64371 36873 64383 36876
rect 64325 36867 64383 36873
rect 64414 36864 64420 36876
rect 64472 36864 64478 36916
rect 64969 36907 65027 36913
rect 64969 36873 64981 36907
rect 65015 36904 65027 36907
rect 65058 36904 65064 36916
rect 65015 36876 65064 36904
rect 65015 36873 65027 36876
rect 64969 36867 65027 36873
rect 65058 36864 65064 36876
rect 65116 36864 65122 36916
rect 65518 36864 65524 36916
rect 65576 36904 65582 36916
rect 65613 36907 65671 36913
rect 65613 36904 65625 36907
rect 65576 36876 65625 36904
rect 65576 36864 65582 36876
rect 65613 36873 65625 36876
rect 65659 36873 65671 36907
rect 65613 36867 65671 36873
rect 66254 36864 66260 36916
rect 66312 36864 66318 36916
rect 66901 36907 66959 36913
rect 66901 36873 66913 36907
rect 66947 36904 66959 36907
rect 66990 36904 66996 36916
rect 66947 36876 66996 36904
rect 66947 36873 66959 36876
rect 66901 36867 66959 36873
rect 66990 36864 66996 36876
rect 67048 36864 67054 36916
rect 67545 36907 67603 36913
rect 67545 36873 67557 36907
rect 67591 36904 67603 36907
rect 67634 36904 67640 36916
rect 67591 36876 67640 36904
rect 67591 36873 67603 36876
rect 67545 36867 67603 36873
rect 67634 36864 67640 36876
rect 67692 36864 67698 36916
rect 68278 36864 68284 36916
rect 68336 36904 68342 36916
rect 68373 36907 68431 36913
rect 68373 36904 68385 36907
rect 68336 36876 68385 36904
rect 68336 36864 68342 36876
rect 68373 36873 68385 36876
rect 68419 36873 68431 36907
rect 68373 36867 68431 36873
rect 68833 36907 68891 36913
rect 68833 36873 68845 36907
rect 68879 36904 68891 36907
rect 68922 36904 68928 36916
rect 68879 36876 68928 36904
rect 68879 36873 68891 36876
rect 68833 36867 68891 36873
rect 68922 36864 68928 36876
rect 68980 36864 68986 36916
rect 69477 36907 69535 36913
rect 69477 36873 69489 36907
rect 69523 36904 69535 36907
rect 69566 36904 69572 36916
rect 69523 36876 69572 36904
rect 69523 36873 69535 36876
rect 69477 36867 69535 36873
rect 69566 36864 69572 36876
rect 69624 36864 69630 36916
rect 70121 36907 70179 36913
rect 70121 36873 70133 36907
rect 70167 36904 70179 36907
rect 70210 36904 70216 36916
rect 70167 36876 70216 36904
rect 70167 36873 70179 36876
rect 70121 36867 70179 36873
rect 70210 36864 70216 36876
rect 70268 36864 70274 36916
rect 70765 36907 70823 36913
rect 70765 36873 70777 36907
rect 70811 36904 70823 36907
rect 70854 36904 70860 36916
rect 70811 36876 70860 36904
rect 70811 36873 70823 36876
rect 70765 36867 70823 36873
rect 70854 36864 70860 36876
rect 70912 36864 70918 36916
rect 71409 36907 71467 36913
rect 71409 36873 71421 36907
rect 71455 36904 71467 36907
rect 71498 36904 71504 36916
rect 71455 36876 71504 36904
rect 71455 36873 71467 36876
rect 71409 36867 71467 36873
rect 71498 36864 71504 36876
rect 71556 36864 71562 36916
rect 72053 36907 72111 36913
rect 72053 36873 72065 36907
rect 72099 36904 72111 36907
rect 72142 36904 72148 36916
rect 72099 36876 72148 36904
rect 72099 36873 72111 36876
rect 72053 36867 72111 36873
rect 72142 36864 72148 36876
rect 72200 36864 72206 36916
rect 72513 36907 72571 36913
rect 72513 36873 72525 36907
rect 72559 36904 72571 36907
rect 72786 36904 72792 36916
rect 72559 36876 72792 36904
rect 72559 36873 72571 36876
rect 72513 36867 72571 36873
rect 72786 36864 72792 36876
rect 72844 36864 72850 36916
rect 72881 36907 72939 36913
rect 72881 36873 72893 36907
rect 72927 36904 72939 36907
rect 73430 36904 73436 36916
rect 72927 36876 73436 36904
rect 72927 36873 72939 36876
rect 72881 36867 72939 36873
rect 73430 36864 73436 36876
rect 73488 36864 73494 36916
rect 35374 36808 36308 36836
rect 32861 36771 32919 36777
rect 32861 36737 32873 36771
rect 32907 36768 32919 36771
rect 33137 36771 33195 36777
rect 33137 36768 33149 36771
rect 32907 36740 33149 36768
rect 32907 36737 32919 36740
rect 32861 36731 32919 36737
rect 33137 36737 33149 36740
rect 33183 36737 33195 36771
rect 33137 36731 33195 36737
rect 35434 36728 35440 36780
rect 35492 36768 35498 36780
rect 35713 36771 35771 36777
rect 35713 36768 35725 36771
rect 35492 36740 35725 36768
rect 35492 36728 35498 36740
rect 35713 36737 35725 36740
rect 35759 36737 35771 36771
rect 35713 36731 35771 36737
rect 35897 36771 35955 36777
rect 35897 36737 35909 36771
rect 35943 36737 35955 36771
rect 36280 36768 36308 36808
rect 36354 36796 36360 36848
rect 36412 36836 36418 36848
rect 36693 36839 36751 36845
rect 36693 36836 36705 36839
rect 36412 36808 36705 36836
rect 36412 36796 36418 36808
rect 36693 36805 36705 36808
rect 36739 36805 36751 36839
rect 36693 36799 36751 36805
rect 36814 36796 36820 36848
rect 36872 36836 36878 36848
rect 36909 36839 36967 36845
rect 36909 36836 36921 36839
rect 36872 36808 36921 36836
rect 36872 36796 36878 36808
rect 36909 36805 36921 36808
rect 36955 36805 36967 36839
rect 40402 36836 40408 36848
rect 39698 36808 40408 36836
rect 36909 36799 36967 36805
rect 40402 36796 40408 36808
rect 40460 36796 40466 36848
rect 44910 36836 44916 36848
rect 44666 36808 44916 36836
rect 44910 36796 44916 36808
rect 44968 36836 44974 36848
rect 45373 36839 45431 36845
rect 45373 36836 45385 36839
rect 44968 36808 45385 36836
rect 44968 36796 44974 36808
rect 45373 36805 45385 36808
rect 45419 36805 45431 36839
rect 45373 36799 45431 36805
rect 37458 36768 37464 36780
rect 36280 36740 37464 36768
rect 35897 36731 35955 36737
rect 2041 36703 2099 36709
rect 2041 36669 2053 36703
rect 2087 36700 2099 36703
rect 2130 36700 2136 36712
rect 2087 36672 2136 36700
rect 2087 36669 2099 36672
rect 2041 36663 2099 36669
rect 2130 36660 2136 36672
rect 2188 36660 2194 36712
rect 32214 36660 32220 36712
rect 32272 36660 32278 36712
rect 33226 36660 33232 36712
rect 33284 36660 33290 36712
rect 33870 36660 33876 36712
rect 33928 36660 33934 36712
rect 34146 36660 34152 36712
rect 34204 36660 34210 36712
rect 35912 36632 35940 36731
rect 37458 36728 37464 36740
rect 37516 36728 37522 36780
rect 40494 36728 40500 36780
rect 40552 36728 40558 36780
rect 40862 36728 40868 36780
rect 40920 36728 40926 36780
rect 41325 36771 41383 36777
rect 41325 36737 41337 36771
rect 41371 36768 41383 36771
rect 41417 36771 41475 36777
rect 41417 36768 41429 36771
rect 41371 36740 41429 36768
rect 41371 36737 41383 36740
rect 41325 36731 41383 36737
rect 41417 36737 41429 36740
rect 41463 36737 41475 36771
rect 41417 36731 41475 36737
rect 41969 36771 42027 36777
rect 41969 36737 41981 36771
rect 42015 36768 42027 36771
rect 42061 36771 42119 36777
rect 42061 36768 42073 36771
rect 42015 36740 42073 36768
rect 42015 36737 42027 36740
rect 41969 36731 42027 36737
rect 42061 36737 42073 36740
rect 42107 36737 42119 36771
rect 42061 36731 42119 36737
rect 42429 36771 42487 36777
rect 42429 36737 42441 36771
rect 42475 36768 42487 36771
rect 42518 36768 42524 36780
rect 42475 36740 42524 36768
rect 42475 36737 42487 36740
rect 42429 36731 42487 36737
rect 42518 36728 42524 36740
rect 42576 36728 42582 36780
rect 43070 36728 43076 36780
rect 43128 36728 43134 36780
rect 45002 36728 45008 36780
rect 45060 36728 45066 36780
rect 45833 36771 45891 36777
rect 45833 36737 45845 36771
rect 45879 36737 45891 36771
rect 45833 36731 45891 36737
rect 36170 36660 36176 36712
rect 36228 36700 36234 36712
rect 38197 36703 38255 36709
rect 38197 36700 38209 36703
rect 36228 36672 38209 36700
rect 36228 36660 36234 36672
rect 38197 36669 38209 36672
rect 38243 36669 38255 36703
rect 38197 36663 38255 36669
rect 38470 36660 38476 36712
rect 38528 36660 38534 36712
rect 42242 36660 42248 36712
rect 42300 36700 42306 36712
rect 43165 36703 43223 36709
rect 43165 36700 43177 36703
rect 42300 36672 43177 36700
rect 42300 36660 42306 36672
rect 43165 36669 43177 36672
rect 43211 36669 43223 36703
rect 43165 36663 43223 36669
rect 43441 36703 43499 36709
rect 43441 36669 43453 36703
rect 43487 36700 43499 36703
rect 43530 36700 43536 36712
rect 43487 36672 43536 36700
rect 43487 36669 43499 36672
rect 43441 36663 43499 36669
rect 43530 36660 43536 36672
rect 43588 36660 43594 36712
rect 45848 36700 45876 36731
rect 45922 36728 45928 36780
rect 45980 36728 45986 36780
rect 47121 36771 47179 36777
rect 47121 36737 47133 36771
rect 47167 36768 47179 36771
rect 47213 36771 47271 36777
rect 47213 36768 47225 36771
rect 47167 36740 47225 36768
rect 47167 36737 47179 36740
rect 47121 36731 47179 36737
rect 47213 36737 47225 36740
rect 47259 36737 47271 36771
rect 47213 36731 47271 36737
rect 47762 36728 47768 36780
rect 47820 36768 47826 36780
rect 47857 36771 47915 36777
rect 47857 36768 47869 36771
rect 47820 36740 47869 36768
rect 47820 36728 47826 36740
rect 47857 36737 47869 36740
rect 47903 36737 47915 36771
rect 47857 36731 47915 36737
rect 48409 36771 48467 36777
rect 48409 36737 48421 36771
rect 48455 36768 48467 36771
rect 48501 36771 48559 36777
rect 48501 36768 48513 36771
rect 48455 36740 48513 36768
rect 48455 36737 48467 36740
rect 48409 36731 48467 36737
rect 48501 36737 48513 36740
rect 48547 36737 48559 36771
rect 48501 36731 48559 36737
rect 48774 36728 48780 36780
rect 48832 36728 48838 36780
rect 49605 36771 49663 36777
rect 49605 36737 49617 36771
rect 49651 36768 49663 36771
rect 49697 36771 49755 36777
rect 49697 36768 49709 36771
rect 49651 36740 49709 36768
rect 49651 36737 49663 36740
rect 49605 36731 49663 36737
rect 49697 36737 49709 36740
rect 49743 36737 49755 36771
rect 49697 36731 49755 36737
rect 50341 36771 50399 36777
rect 50341 36737 50353 36771
rect 50387 36768 50399 36771
rect 50433 36771 50491 36777
rect 50433 36768 50445 36771
rect 50387 36740 50445 36768
rect 50387 36737 50399 36740
rect 50341 36731 50399 36737
rect 50433 36737 50445 36740
rect 50479 36737 50491 36771
rect 50433 36731 50491 36737
rect 50985 36771 51043 36777
rect 50985 36737 50997 36771
rect 51031 36768 51043 36771
rect 51077 36771 51135 36777
rect 51077 36768 51089 36771
rect 51031 36740 51089 36768
rect 51031 36737 51043 36740
rect 50985 36731 51043 36737
rect 51077 36737 51089 36740
rect 51123 36737 51135 36771
rect 51077 36731 51135 36737
rect 51629 36771 51687 36777
rect 51629 36737 51641 36771
rect 51675 36768 51687 36771
rect 51721 36771 51779 36777
rect 51721 36768 51733 36771
rect 51675 36740 51733 36768
rect 51675 36737 51687 36740
rect 51629 36731 51687 36737
rect 51721 36737 51733 36740
rect 51767 36737 51779 36771
rect 51721 36731 51779 36737
rect 52273 36771 52331 36777
rect 52273 36737 52285 36771
rect 52319 36768 52331 36771
rect 52365 36771 52423 36777
rect 52365 36768 52377 36771
rect 52319 36740 52377 36768
rect 52319 36737 52331 36740
rect 52273 36731 52331 36737
rect 52365 36737 52377 36740
rect 52411 36737 52423 36771
rect 52365 36731 52423 36737
rect 52914 36728 52920 36780
rect 52972 36768 52978 36780
rect 53009 36771 53067 36777
rect 53009 36768 53021 36771
rect 52972 36740 53021 36768
rect 52972 36728 52978 36740
rect 53009 36737 53021 36740
rect 53055 36737 53067 36771
rect 53009 36731 53067 36737
rect 53282 36728 53288 36780
rect 53340 36728 53346 36780
rect 54113 36771 54171 36777
rect 54113 36737 54125 36771
rect 54159 36768 54171 36771
rect 54205 36771 54263 36777
rect 54205 36768 54217 36771
rect 54159 36740 54217 36768
rect 54159 36737 54171 36740
rect 54113 36731 54171 36737
rect 54205 36737 54217 36740
rect 54251 36737 54263 36771
rect 54205 36731 54263 36737
rect 54757 36771 54815 36777
rect 54757 36737 54769 36771
rect 54803 36768 54815 36771
rect 54849 36771 54907 36777
rect 54849 36768 54861 36771
rect 54803 36740 54861 36768
rect 54803 36737 54815 36740
rect 54757 36731 54815 36737
rect 54849 36737 54861 36740
rect 54895 36737 54907 36771
rect 54849 36731 54907 36737
rect 55401 36771 55459 36777
rect 55401 36737 55413 36771
rect 55447 36768 55459 36771
rect 55493 36771 55551 36777
rect 55493 36768 55505 36771
rect 55447 36740 55505 36768
rect 55447 36737 55459 36740
rect 55401 36731 55459 36737
rect 55493 36737 55505 36740
rect 55539 36737 55551 36771
rect 55493 36731 55551 36737
rect 56045 36771 56103 36777
rect 56045 36737 56057 36771
rect 56091 36768 56103 36771
rect 56137 36771 56195 36777
rect 56137 36768 56149 36771
rect 56091 36740 56149 36768
rect 56091 36737 56103 36740
rect 56045 36731 56103 36737
rect 56137 36737 56149 36740
rect 56183 36737 56195 36771
rect 56137 36731 56195 36737
rect 56781 36771 56839 36777
rect 56781 36737 56793 36771
rect 56827 36768 56839 36771
rect 56873 36771 56931 36777
rect 56873 36768 56885 36771
rect 56827 36740 56885 36768
rect 56827 36737 56839 36740
rect 56781 36731 56839 36737
rect 56873 36737 56885 36740
rect 56919 36737 56931 36771
rect 56873 36731 56931 36737
rect 57425 36771 57483 36777
rect 57425 36737 57437 36771
rect 57471 36768 57483 36771
rect 57517 36771 57575 36777
rect 57517 36768 57529 36771
rect 57471 36740 57529 36768
rect 57471 36737 57483 36740
rect 57425 36731 57483 36737
rect 57517 36737 57529 36740
rect 57563 36737 57575 36771
rect 57517 36731 57575 36737
rect 58066 36728 58072 36780
rect 58124 36768 58130 36780
rect 58161 36771 58219 36777
rect 58161 36768 58173 36771
rect 58124 36740 58173 36768
rect 58124 36728 58130 36740
rect 58161 36737 58173 36740
rect 58207 36737 58219 36771
rect 58161 36731 58219 36737
rect 58713 36771 58771 36777
rect 58713 36737 58725 36771
rect 58759 36768 58771 36771
rect 58805 36771 58863 36777
rect 58805 36768 58817 36771
rect 58759 36740 58817 36768
rect 58759 36737 58771 36740
rect 58713 36731 58771 36737
rect 58805 36737 58817 36740
rect 58851 36737 58863 36771
rect 58805 36731 58863 36737
rect 59357 36771 59415 36777
rect 59357 36737 59369 36771
rect 59403 36768 59415 36771
rect 59449 36771 59507 36777
rect 59449 36768 59461 36771
rect 59403 36740 59461 36768
rect 59403 36737 59415 36740
rect 59357 36731 59415 36737
rect 59449 36737 59461 36740
rect 59495 36737 59507 36771
rect 59449 36731 59507 36737
rect 60093 36771 60151 36777
rect 60093 36737 60105 36771
rect 60139 36737 60151 36771
rect 60093 36731 60151 36737
rect 46201 36703 46259 36709
rect 46201 36700 46213 36703
rect 45848 36672 46213 36700
rect 46201 36669 46213 36672
rect 46247 36669 46259 36703
rect 60108 36700 60136 36731
rect 60642 36728 60648 36780
rect 60700 36728 60706 36780
rect 61010 36728 61016 36780
rect 61068 36728 61074 36780
rect 61841 36771 61899 36777
rect 61841 36737 61853 36771
rect 61887 36768 61899 36771
rect 61933 36771 61991 36777
rect 61933 36768 61945 36771
rect 61887 36740 61945 36768
rect 61887 36737 61899 36740
rect 61841 36731 61899 36737
rect 61933 36737 61945 36740
rect 61979 36737 61991 36771
rect 61933 36731 61991 36737
rect 62577 36771 62635 36777
rect 62577 36737 62589 36771
rect 62623 36768 62635 36771
rect 62669 36771 62727 36777
rect 62669 36768 62681 36771
rect 62623 36740 62681 36768
rect 62623 36737 62635 36740
rect 62577 36731 62635 36737
rect 62669 36737 62681 36740
rect 62715 36737 62727 36771
rect 62669 36731 62727 36737
rect 63037 36771 63095 36777
rect 63037 36737 63049 36771
rect 63083 36768 63095 36771
rect 63126 36768 63132 36780
rect 63083 36740 63132 36768
rect 63083 36737 63095 36740
rect 63037 36731 63095 36737
rect 63126 36728 63132 36740
rect 63184 36728 63190 36780
rect 63865 36771 63923 36777
rect 63865 36737 63877 36771
rect 63911 36768 63923 36771
rect 63957 36771 64015 36777
rect 63957 36768 63969 36771
rect 63911 36740 63969 36768
rect 63911 36737 63923 36740
rect 63865 36731 63923 36737
rect 63957 36737 63969 36740
rect 64003 36737 64015 36771
rect 63957 36731 64015 36737
rect 64509 36771 64567 36777
rect 64509 36737 64521 36771
rect 64555 36768 64567 36771
rect 64601 36771 64659 36777
rect 64601 36768 64613 36771
rect 64555 36740 64613 36768
rect 64555 36737 64567 36740
rect 64509 36731 64567 36737
rect 64601 36737 64613 36740
rect 64647 36737 64659 36771
rect 64601 36731 64659 36737
rect 65153 36771 65211 36777
rect 65153 36737 65165 36771
rect 65199 36768 65211 36771
rect 65245 36771 65303 36777
rect 65245 36768 65257 36771
rect 65199 36740 65257 36768
rect 65199 36737 65211 36740
rect 65153 36731 65211 36737
rect 65245 36737 65257 36740
rect 65291 36737 65303 36771
rect 65245 36731 65303 36737
rect 65797 36771 65855 36777
rect 65797 36737 65809 36771
rect 65843 36768 65855 36771
rect 65889 36771 65947 36777
rect 65889 36768 65901 36771
rect 65843 36740 65901 36768
rect 65843 36737 65855 36740
rect 65797 36731 65855 36737
rect 65889 36737 65901 36740
rect 65935 36737 65947 36771
rect 65889 36731 65947 36737
rect 66441 36771 66499 36777
rect 66441 36737 66453 36771
rect 66487 36768 66499 36771
rect 66533 36771 66591 36777
rect 66533 36768 66545 36771
rect 66487 36740 66545 36768
rect 66487 36737 66499 36740
rect 66441 36731 66499 36737
rect 66533 36737 66545 36740
rect 66579 36737 66591 36771
rect 66533 36731 66591 36737
rect 67085 36771 67143 36777
rect 67085 36737 67097 36771
rect 67131 36768 67143 36771
rect 67177 36771 67235 36777
rect 67177 36768 67189 36771
rect 67131 36740 67189 36768
rect 67131 36737 67143 36740
rect 67085 36731 67143 36737
rect 67177 36737 67189 36740
rect 67223 36737 67235 36771
rect 67177 36731 67235 36737
rect 67729 36771 67787 36777
rect 67729 36737 67741 36771
rect 67775 36768 67787 36771
rect 67821 36771 67879 36777
rect 67821 36768 67833 36771
rect 67775 36740 67833 36768
rect 67775 36737 67787 36740
rect 67729 36731 67787 36737
rect 67821 36737 67833 36740
rect 67867 36737 67879 36771
rect 67821 36731 67879 36737
rect 68189 36771 68247 36777
rect 68189 36737 68201 36771
rect 68235 36768 68247 36771
rect 68278 36768 68284 36780
rect 68235 36740 68284 36768
rect 68235 36737 68247 36740
rect 68189 36731 68247 36737
rect 68278 36728 68284 36740
rect 68336 36728 68342 36780
rect 69017 36771 69075 36777
rect 69017 36737 69029 36771
rect 69063 36768 69075 36771
rect 69109 36771 69167 36777
rect 69109 36768 69121 36771
rect 69063 36740 69121 36768
rect 69063 36737 69075 36740
rect 69017 36731 69075 36737
rect 69109 36737 69121 36740
rect 69155 36737 69167 36771
rect 69109 36731 69167 36737
rect 69661 36771 69719 36777
rect 69661 36737 69673 36771
rect 69707 36768 69719 36771
rect 69753 36771 69811 36777
rect 69753 36768 69765 36771
rect 69707 36740 69765 36768
rect 69707 36737 69719 36740
rect 69661 36731 69719 36737
rect 69753 36737 69765 36740
rect 69799 36737 69811 36771
rect 69753 36731 69811 36737
rect 70305 36771 70363 36777
rect 70305 36737 70317 36771
rect 70351 36768 70363 36771
rect 70397 36771 70455 36777
rect 70397 36768 70409 36771
rect 70351 36740 70409 36768
rect 70351 36737 70363 36740
rect 70305 36731 70363 36737
rect 70397 36737 70409 36740
rect 70443 36737 70455 36771
rect 70397 36731 70455 36737
rect 70949 36771 71007 36777
rect 70949 36737 70961 36771
rect 70995 36768 71007 36771
rect 71041 36771 71099 36777
rect 71041 36768 71053 36771
rect 70995 36740 71053 36768
rect 70995 36737 71007 36740
rect 70949 36731 71007 36737
rect 71041 36737 71053 36740
rect 71087 36737 71099 36771
rect 71041 36731 71099 36737
rect 71593 36771 71651 36777
rect 71593 36737 71605 36771
rect 71639 36768 71651 36771
rect 71685 36771 71743 36777
rect 71685 36768 71697 36771
rect 71639 36740 71697 36768
rect 71639 36737 71651 36740
rect 71593 36731 71651 36737
rect 71685 36737 71697 36740
rect 71731 36737 71743 36771
rect 71685 36731 71743 36737
rect 72234 36728 72240 36780
rect 72292 36728 72298 36780
rect 72697 36771 72755 36777
rect 72697 36737 72709 36771
rect 72743 36737 72755 36771
rect 72697 36731 72755 36737
rect 73065 36771 73123 36777
rect 73065 36737 73077 36771
rect 73111 36768 73123 36771
rect 73617 36771 73675 36777
rect 73617 36768 73629 36771
rect 73111 36740 73629 36768
rect 73111 36737 73123 36740
rect 73065 36731 73123 36737
rect 73617 36737 73629 36740
rect 73663 36737 73675 36771
rect 73617 36731 73675 36737
rect 60737 36703 60795 36709
rect 60737 36700 60749 36703
rect 60108 36672 60749 36700
rect 46201 36663 46259 36669
rect 60737 36669 60749 36672
rect 60783 36669 60795 36703
rect 72712 36700 72740 36731
rect 73341 36703 73399 36709
rect 73341 36700 73353 36703
rect 72712 36672 73353 36700
rect 60737 36663 60795 36669
rect 73341 36669 73353 36672
rect 73387 36669 73399 36703
rect 73341 36663 73399 36669
rect 36078 36632 36084 36644
rect 35912 36604 36084 36632
rect 36078 36592 36084 36604
rect 36136 36632 36142 36644
rect 36541 36635 36599 36641
rect 36541 36632 36553 36635
rect 36136 36604 36553 36632
rect 36136 36592 36142 36604
rect 36541 36601 36553 36604
rect 36587 36601 36599 36635
rect 36541 36595 36599 36601
rect 33413 36567 33471 36573
rect 33413 36533 33425 36567
rect 33459 36564 33471 36567
rect 33502 36564 33508 36576
rect 33459 36536 33508 36564
rect 33459 36533 33471 36536
rect 33413 36527 33471 36533
rect 33502 36524 33508 36536
rect 33560 36524 33566 36576
rect 35710 36524 35716 36576
rect 35768 36564 35774 36576
rect 35897 36567 35955 36573
rect 35897 36564 35909 36567
rect 35768 36536 35909 36564
rect 35768 36524 35774 36536
rect 35897 36533 35909 36536
rect 35943 36533 35955 36567
rect 35897 36527 35955 36533
rect 36725 36567 36783 36573
rect 36725 36533 36737 36567
rect 36771 36564 36783 36567
rect 37274 36564 37280 36576
rect 36771 36536 37280 36564
rect 36771 36533 36783 36536
rect 36725 36527 36783 36533
rect 37274 36524 37280 36536
rect 37332 36524 37338 36576
rect 39482 36524 39488 36576
rect 39540 36564 39546 36576
rect 39945 36567 40003 36573
rect 39945 36564 39957 36567
rect 39540 36536 39957 36564
rect 39540 36524 39546 36536
rect 39945 36533 39957 36536
rect 39991 36533 40003 36567
rect 39945 36527 40003 36533
rect 44542 36524 44548 36576
rect 44600 36564 44606 36576
rect 44913 36567 44971 36573
rect 44913 36564 44925 36567
rect 44600 36536 44925 36564
rect 44600 36524 44606 36536
rect 44913 36533 44925 36536
rect 44959 36533 44971 36567
rect 44913 36527 44971 36533
rect 1104 36474 78844 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 78844 36474
rect 1104 36400 78844 36422
rect 1302 36320 1308 36372
rect 1360 36360 1366 36372
rect 2317 36363 2375 36369
rect 2317 36360 2329 36363
rect 1360 36332 2329 36360
rect 1360 36320 1366 36332
rect 2317 36329 2329 36332
rect 2363 36329 2375 36363
rect 2317 36323 2375 36329
rect 32033 36363 32091 36369
rect 32033 36329 32045 36363
rect 32079 36360 32091 36363
rect 32214 36360 32220 36372
rect 32079 36332 32220 36360
rect 32079 36329 32091 36332
rect 32033 36323 32091 36329
rect 32214 36320 32220 36332
rect 32272 36320 32278 36372
rect 34146 36320 34152 36372
rect 34204 36360 34210 36372
rect 34977 36363 35035 36369
rect 34977 36360 34989 36363
rect 34204 36332 34989 36360
rect 34204 36320 34210 36332
rect 34977 36329 34989 36332
rect 35023 36329 35035 36363
rect 34977 36323 35035 36329
rect 35621 36363 35679 36369
rect 35621 36329 35633 36363
rect 35667 36360 35679 36363
rect 35667 36332 37504 36360
rect 35667 36329 35679 36332
rect 35621 36323 35679 36329
rect 34698 36252 34704 36304
rect 34756 36292 34762 36304
rect 35636 36292 35664 36323
rect 34756 36264 35664 36292
rect 35897 36295 35955 36301
rect 34756 36252 34762 36264
rect 35897 36261 35909 36295
rect 35943 36292 35955 36295
rect 37476 36292 37504 36332
rect 38470 36320 38476 36372
rect 38528 36360 38534 36372
rect 38749 36363 38807 36369
rect 38749 36360 38761 36363
rect 38528 36332 38761 36360
rect 38528 36320 38534 36332
rect 38749 36329 38761 36332
rect 38795 36329 38807 36363
rect 38749 36323 38807 36329
rect 39206 36320 39212 36372
rect 39264 36360 39270 36372
rect 39669 36363 39727 36369
rect 39669 36360 39681 36363
rect 39264 36332 39681 36360
rect 39264 36320 39270 36332
rect 39669 36329 39681 36332
rect 39715 36329 39727 36363
rect 39669 36323 39727 36329
rect 42518 36320 42524 36372
rect 42576 36320 42582 36372
rect 43070 36320 43076 36372
rect 43128 36320 43134 36372
rect 43530 36320 43536 36372
rect 43588 36320 43594 36372
rect 43714 36320 43720 36372
rect 43772 36320 43778 36372
rect 44358 36320 44364 36372
rect 44416 36320 44422 36372
rect 44637 36363 44695 36369
rect 44637 36329 44649 36363
rect 44683 36360 44695 36363
rect 45002 36360 45008 36372
rect 44683 36332 45008 36360
rect 44683 36329 44695 36332
rect 44637 36323 44695 36329
rect 45002 36320 45008 36332
rect 45060 36320 45066 36372
rect 47762 36320 47768 36372
rect 47820 36320 47826 36372
rect 48774 36320 48780 36372
rect 48832 36320 48838 36372
rect 52914 36320 52920 36372
rect 52972 36320 52978 36372
rect 53282 36320 53288 36372
rect 53340 36320 53346 36372
rect 58066 36320 58072 36372
rect 58124 36320 58130 36372
rect 60642 36320 60648 36372
rect 60700 36320 60706 36372
rect 61010 36320 61016 36372
rect 61068 36320 61074 36372
rect 63126 36320 63132 36372
rect 63184 36320 63190 36372
rect 68278 36320 68284 36372
rect 68336 36320 68342 36372
rect 72234 36320 72240 36372
rect 72292 36320 72298 36372
rect 39022 36292 39028 36304
rect 35943 36264 36308 36292
rect 37476 36264 39028 36292
rect 35943 36261 35955 36264
rect 35897 36255 35955 36261
rect 2501 36227 2559 36233
rect 2501 36224 2513 36227
rect 2056 36196 2513 36224
rect 2056 36165 2084 36196
rect 2501 36193 2513 36196
rect 2547 36193 2559 36227
rect 2501 36187 2559 36193
rect 33502 36184 33508 36236
rect 33560 36184 33566 36236
rect 33781 36227 33839 36233
rect 33781 36193 33793 36227
rect 33827 36224 33839 36227
rect 33870 36224 33876 36236
rect 33827 36196 33876 36224
rect 33827 36193 33839 36196
rect 33781 36187 33839 36193
rect 33870 36184 33876 36196
rect 33928 36224 33934 36236
rect 36170 36224 36176 36236
rect 33928 36196 36176 36224
rect 33928 36184 33934 36196
rect 36170 36184 36176 36196
rect 36228 36184 36234 36236
rect 36280 36224 36308 36264
rect 39022 36252 39028 36264
rect 39080 36252 39086 36304
rect 36449 36227 36507 36233
rect 36449 36224 36461 36227
rect 36280 36196 36461 36224
rect 36449 36193 36461 36196
rect 36495 36193 36507 36227
rect 36449 36187 36507 36193
rect 38194 36184 38200 36236
rect 38252 36224 38258 36236
rect 38252 36196 39344 36224
rect 38252 36184 38258 36196
rect 2041 36159 2099 36165
rect 2041 36125 2053 36159
rect 2087 36125 2099 36159
rect 2041 36119 2099 36125
rect 2130 36116 2136 36168
rect 2188 36116 2194 36168
rect 34977 36159 35035 36165
rect 34977 36125 34989 36159
rect 35023 36125 35035 36159
rect 34977 36119 35035 36125
rect 34992 36088 35020 36119
rect 35158 36116 35164 36168
rect 35216 36116 35222 36168
rect 35897 36159 35955 36165
rect 35897 36125 35909 36159
rect 35943 36125 35955 36159
rect 35897 36119 35955 36125
rect 35710 36088 35716 36100
rect 33074 36060 34008 36088
rect 34992 36060 35716 36088
rect 934 35980 940 36032
rect 992 36020 998 36032
rect 33980 36029 34008 36060
rect 35710 36048 35716 36060
rect 35768 36048 35774 36100
rect 35912 36088 35940 36119
rect 36078 36116 36084 36168
rect 36136 36116 36142 36168
rect 38565 36159 38623 36165
rect 38565 36156 38577 36159
rect 37936 36128 38577 36156
rect 36722 36088 36728 36100
rect 35912 36060 36728 36088
rect 36722 36048 36728 36060
rect 36780 36048 36786 36100
rect 37458 36048 37464 36100
rect 37516 36048 37522 36100
rect 1857 36023 1915 36029
rect 1857 36020 1869 36023
rect 992 35992 1869 36020
rect 992 35980 998 35992
rect 1857 35989 1869 35992
rect 1903 35989 1915 36023
rect 1857 35983 1915 35989
rect 33965 36023 34023 36029
rect 33965 35989 33977 36023
rect 34011 36020 34023 36023
rect 34606 36020 34612 36032
rect 34011 35992 34612 36020
rect 34011 35989 34023 35992
rect 33965 35983 34023 35989
rect 34606 35980 34612 35992
rect 34664 35980 34670 36032
rect 36354 35980 36360 36032
rect 36412 36020 36418 36032
rect 37936 36029 37964 36128
rect 38565 36125 38577 36128
rect 38611 36125 38623 36159
rect 38565 36119 38623 36125
rect 38933 36159 38991 36165
rect 38933 36125 38945 36159
rect 38979 36156 38991 36159
rect 39022 36156 39028 36168
rect 38979 36128 39028 36156
rect 38979 36125 38991 36128
rect 38933 36119 38991 36125
rect 39022 36116 39028 36128
rect 39080 36116 39086 36168
rect 39206 36116 39212 36168
rect 39264 36116 39270 36168
rect 39316 36165 39344 36196
rect 42242 36184 42248 36236
rect 42300 36184 42306 36236
rect 45738 36184 45744 36236
rect 45796 36224 45802 36236
rect 46293 36227 46351 36233
rect 46293 36224 46305 36227
rect 45796 36196 46305 36224
rect 45796 36184 45802 36196
rect 46293 36193 46305 36196
rect 46339 36193 46351 36227
rect 46293 36187 46351 36193
rect 39301 36159 39359 36165
rect 39301 36125 39313 36159
rect 39347 36125 39359 36159
rect 39301 36119 39359 36125
rect 44082 36116 44088 36168
rect 44140 36116 44146 36168
rect 44177 36159 44235 36165
rect 44177 36125 44189 36159
rect 44223 36156 44235 36159
rect 44358 36156 44364 36168
rect 44223 36128 44364 36156
rect 44223 36125 44235 36128
rect 44177 36119 44235 36125
rect 44358 36116 44364 36128
rect 44416 36116 44422 36168
rect 46106 36116 46112 36168
rect 46164 36116 46170 36168
rect 46385 36159 46443 36165
rect 46385 36125 46397 36159
rect 46431 36156 46443 36159
rect 46474 36156 46480 36168
rect 46431 36128 46480 36156
rect 46431 36125 46443 36128
rect 46385 36119 46443 36125
rect 46474 36116 46480 36128
rect 46532 36116 46538 36168
rect 38378 36048 38384 36100
rect 38436 36088 38442 36100
rect 38436 36060 39252 36088
rect 38436 36048 38442 36060
rect 37921 36023 37979 36029
rect 37921 36020 37933 36023
rect 36412 35992 37933 36020
rect 36412 35980 36418 35992
rect 37921 35989 37933 35992
rect 37967 35989 37979 36023
rect 37921 35983 37979 35989
rect 38010 35980 38016 36032
rect 38068 35980 38074 36032
rect 39114 35980 39120 36032
rect 39172 35980 39178 36032
rect 39224 36020 39252 36060
rect 39482 36048 39488 36100
rect 39540 36048 39546 36100
rect 40402 36048 40408 36100
rect 40460 36088 40466 36100
rect 40460 36060 40802 36088
rect 40460 36048 40466 36060
rect 41966 36048 41972 36100
rect 42024 36048 42030 36100
rect 39500 36020 39528 36048
rect 39224 35992 39528 36020
rect 40497 36023 40555 36029
rect 40497 35989 40509 36023
rect 40543 36020 40555 36023
rect 40678 36020 40684 36032
rect 40543 35992 40684 36020
rect 40543 35989 40555 35992
rect 40497 35983 40555 35989
rect 40678 35980 40684 35992
rect 40736 35980 40742 36032
rect 43717 36023 43775 36029
rect 43717 35989 43729 36023
rect 43763 36020 43775 36023
rect 44266 36020 44272 36032
rect 43763 35992 44272 36020
rect 43763 35989 43775 35992
rect 43717 35983 43775 35989
rect 44266 35980 44272 35992
rect 44324 35980 44330 36032
rect 45922 35980 45928 36032
rect 45980 35980 45986 36032
rect 1104 35930 78844 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 66314 35930
rect 66366 35878 66378 35930
rect 66430 35878 66442 35930
rect 66494 35878 66506 35930
rect 66558 35878 66570 35930
rect 66622 35878 78844 35930
rect 1104 35856 78844 35878
rect 32674 35816 32680 35828
rect 32324 35788 32680 35816
rect 32324 35757 32352 35788
rect 32674 35776 32680 35788
rect 32732 35776 32738 35828
rect 32769 35819 32827 35825
rect 32769 35785 32781 35819
rect 32815 35816 32827 35819
rect 33226 35816 33232 35828
rect 32815 35788 33232 35816
rect 32815 35785 32827 35788
rect 32769 35779 32827 35785
rect 32309 35751 32367 35757
rect 32309 35717 32321 35751
rect 32355 35717 32367 35751
rect 32784 35748 32812 35779
rect 33226 35776 33232 35788
rect 33284 35776 33290 35828
rect 35158 35776 35164 35828
rect 35216 35816 35222 35828
rect 35342 35816 35348 35828
rect 35216 35788 35348 35816
rect 35216 35776 35222 35788
rect 35342 35776 35348 35788
rect 35400 35816 35406 35828
rect 36081 35819 36139 35825
rect 36081 35816 36093 35819
rect 35400 35788 36093 35816
rect 35400 35776 35406 35788
rect 36081 35785 36093 35788
rect 36127 35785 36139 35819
rect 36081 35779 36139 35785
rect 36262 35776 36268 35828
rect 36320 35816 36326 35828
rect 36357 35819 36415 35825
rect 36357 35816 36369 35819
rect 36320 35788 36369 35816
rect 36320 35776 36326 35788
rect 36357 35785 36369 35788
rect 36403 35785 36415 35819
rect 36814 35816 36820 35828
rect 36357 35779 36415 35785
rect 36648 35788 36820 35816
rect 36648 35757 36676 35788
rect 36814 35776 36820 35788
rect 36872 35816 36878 35828
rect 38381 35819 38439 35825
rect 36872 35788 38148 35816
rect 36872 35776 36878 35788
rect 32309 35711 32367 35717
rect 32692 35720 32812 35748
rect 36633 35751 36691 35757
rect 2041 35683 2099 35689
rect 2041 35649 2053 35683
rect 2087 35680 2099 35683
rect 2133 35683 2191 35689
rect 2133 35680 2145 35683
rect 2087 35652 2145 35680
rect 2087 35649 2099 35652
rect 2041 35643 2099 35649
rect 2133 35649 2145 35652
rect 2179 35649 2191 35683
rect 2133 35643 2191 35649
rect 31757 35683 31815 35689
rect 31757 35649 31769 35683
rect 31803 35680 31815 35683
rect 32125 35683 32183 35689
rect 32125 35680 32137 35683
rect 31803 35652 32137 35680
rect 31803 35649 31815 35652
rect 31757 35643 31815 35649
rect 32125 35649 32137 35652
rect 32171 35649 32183 35683
rect 32125 35643 32183 35649
rect 32398 35640 32404 35692
rect 32456 35680 32462 35692
rect 32493 35683 32551 35689
rect 32493 35680 32505 35683
rect 32456 35652 32505 35680
rect 32456 35640 32462 35652
rect 32493 35649 32505 35652
rect 32539 35680 32551 35683
rect 32585 35683 32643 35689
rect 32585 35680 32597 35683
rect 32539 35652 32597 35680
rect 32539 35649 32551 35652
rect 32493 35643 32551 35649
rect 32585 35649 32597 35652
rect 32631 35649 32643 35683
rect 32585 35643 32643 35649
rect 31941 35615 31999 35621
rect 31941 35581 31953 35615
rect 31987 35612 31999 35615
rect 32692 35612 32720 35720
rect 36633 35717 36645 35751
rect 36679 35717 36691 35751
rect 36633 35711 36691 35717
rect 37001 35751 37059 35757
rect 37001 35717 37013 35751
rect 37047 35748 37059 35751
rect 38010 35748 38016 35760
rect 37047 35720 38016 35748
rect 37047 35717 37059 35720
rect 37001 35711 37059 35717
rect 38010 35708 38016 35720
rect 38068 35708 38074 35760
rect 38120 35748 38148 35788
rect 38381 35785 38393 35819
rect 38427 35816 38439 35819
rect 39114 35816 39120 35828
rect 38427 35788 39120 35816
rect 38427 35785 38439 35788
rect 38381 35779 38439 35785
rect 39114 35776 39120 35788
rect 39172 35776 39178 35828
rect 40773 35819 40831 35825
rect 40773 35785 40785 35819
rect 40819 35816 40831 35819
rect 41525 35819 41583 35825
rect 41525 35816 41537 35819
rect 40819 35788 41537 35816
rect 40819 35785 40831 35788
rect 40773 35779 40831 35785
rect 41525 35785 41537 35788
rect 41571 35785 41583 35819
rect 41525 35779 41583 35785
rect 41693 35819 41751 35825
rect 41693 35785 41705 35819
rect 41739 35816 41751 35819
rect 41966 35816 41972 35828
rect 41739 35788 41972 35816
rect 41739 35785 41751 35788
rect 41693 35779 41751 35785
rect 41966 35776 41972 35788
rect 42024 35776 42030 35828
rect 44266 35776 44272 35828
rect 44324 35816 44330 35828
rect 44361 35819 44419 35825
rect 44361 35816 44373 35819
rect 44324 35788 44373 35816
rect 44324 35776 44330 35788
rect 44361 35785 44373 35788
rect 44407 35785 44419 35819
rect 44361 35779 44419 35785
rect 46474 35776 46480 35828
rect 46532 35816 46538 35828
rect 47305 35819 47363 35825
rect 47305 35816 47317 35819
rect 46532 35788 47317 35816
rect 46532 35776 46538 35788
rect 47305 35785 47317 35788
rect 47351 35785 47363 35819
rect 47305 35779 47363 35785
rect 41322 35748 41328 35760
rect 38120 35720 38424 35748
rect 38396 35692 38424 35720
rect 40604 35720 40908 35748
rect 41283 35720 41328 35748
rect 32766 35640 32772 35692
rect 32824 35640 32830 35692
rect 36265 35683 36323 35689
rect 36265 35649 36277 35683
rect 36311 35680 36323 35683
rect 36354 35680 36360 35692
rect 36311 35652 36360 35680
rect 36311 35649 36323 35652
rect 36265 35643 36323 35649
rect 36354 35640 36360 35652
rect 36412 35640 36418 35692
rect 36449 35683 36507 35689
rect 36449 35649 36461 35683
rect 36495 35680 36507 35683
rect 36725 35683 36783 35689
rect 36725 35680 36737 35683
rect 36495 35652 36737 35680
rect 36495 35649 36507 35652
rect 36449 35643 36507 35649
rect 36725 35649 36737 35652
rect 36771 35680 36783 35683
rect 37274 35680 37280 35692
rect 36771 35652 37280 35680
rect 36771 35649 36783 35652
rect 36725 35643 36783 35649
rect 37274 35640 37280 35652
rect 37332 35680 37338 35692
rect 38194 35680 38200 35692
rect 37332 35652 38200 35680
rect 37332 35640 37338 35652
rect 38194 35640 38200 35652
rect 38252 35640 38258 35692
rect 38378 35640 38384 35692
rect 38436 35640 38442 35692
rect 40604 35689 40632 35720
rect 40880 35692 40908 35720
rect 41322 35708 41328 35720
rect 41380 35748 41386 35760
rect 43714 35748 43720 35760
rect 41380 35720 43720 35748
rect 41380 35708 41386 35720
rect 43714 35708 43720 35720
rect 43772 35708 43778 35760
rect 45738 35748 45744 35760
rect 45526 35720 45744 35748
rect 40589 35683 40647 35689
rect 40589 35649 40601 35683
rect 40635 35649 40647 35683
rect 40589 35643 40647 35649
rect 40678 35640 40684 35692
rect 40736 35680 40742 35692
rect 40773 35683 40831 35689
rect 40773 35680 40785 35683
rect 40736 35652 40785 35680
rect 40736 35640 40742 35652
rect 40773 35649 40785 35652
rect 40819 35649 40831 35683
rect 40773 35643 40831 35649
rect 31987 35584 32720 35612
rect 40788 35612 40816 35643
rect 40862 35640 40868 35692
rect 40920 35640 40926 35692
rect 41049 35683 41107 35689
rect 41049 35649 41061 35683
rect 41095 35649 41107 35683
rect 41049 35643 41107 35649
rect 41064 35612 41092 35643
rect 44542 35640 44548 35692
rect 44600 35640 44606 35692
rect 44726 35640 44732 35692
rect 44784 35640 44790 35692
rect 44821 35683 44879 35689
rect 44821 35649 44833 35683
rect 44867 35680 44879 35683
rect 45526 35680 45554 35720
rect 45738 35708 45744 35720
rect 45796 35708 45802 35760
rect 45833 35751 45891 35757
rect 45833 35717 45845 35751
rect 45879 35748 45891 35751
rect 45922 35748 45928 35760
rect 45879 35720 45928 35748
rect 45879 35717 45891 35720
rect 45833 35711 45891 35717
rect 45922 35708 45928 35720
rect 45980 35708 45986 35760
rect 44867 35652 45554 35680
rect 46966 35652 47716 35680
rect 44867 35649 44879 35652
rect 44821 35643 44879 35649
rect 40788 35584 41092 35612
rect 31987 35581 31999 35584
rect 31941 35575 31999 35581
rect 42242 35572 42248 35624
rect 42300 35612 42306 35624
rect 45557 35615 45615 35621
rect 45557 35612 45569 35615
rect 42300 35584 45569 35612
rect 42300 35572 42306 35584
rect 45557 35581 45569 35584
rect 45603 35612 45615 35615
rect 45922 35612 45928 35624
rect 45603 35584 45928 35612
rect 45603 35581 45615 35584
rect 45557 35575 45615 35581
rect 45922 35572 45928 35584
rect 45980 35572 45986 35624
rect 36722 35504 36728 35556
rect 36780 35544 36786 35556
rect 37001 35547 37059 35553
rect 37001 35544 37013 35547
rect 36780 35516 37013 35544
rect 36780 35504 36786 35516
rect 37001 35513 37013 35516
rect 37047 35513 37059 35547
rect 37001 35507 37059 35513
rect 934 35436 940 35488
rect 992 35476 998 35488
rect 1857 35479 1915 35485
rect 1857 35476 1869 35479
rect 992 35448 1869 35476
rect 992 35436 998 35448
rect 1857 35445 1869 35448
rect 1903 35445 1915 35479
rect 1857 35439 1915 35445
rect 31478 35436 31484 35488
rect 31536 35476 31542 35488
rect 47688 35485 47716 35652
rect 31573 35479 31631 35485
rect 31573 35476 31585 35479
rect 31536 35448 31585 35476
rect 31536 35436 31542 35448
rect 31573 35445 31585 35448
rect 31619 35445 31631 35479
rect 31573 35439 31631 35445
rect 41233 35479 41291 35485
rect 41233 35445 41245 35479
rect 41279 35476 41291 35479
rect 41509 35479 41567 35485
rect 41509 35476 41521 35479
rect 41279 35448 41521 35476
rect 41279 35445 41291 35448
rect 41233 35439 41291 35445
rect 41509 35445 41521 35448
rect 41555 35445 41567 35479
rect 41509 35439 41567 35445
rect 47673 35479 47731 35485
rect 47673 35445 47685 35479
rect 47719 35476 47731 35479
rect 48774 35476 48780 35488
rect 47719 35448 48780 35476
rect 47719 35445 47731 35448
rect 47673 35439 47731 35445
rect 48774 35436 48780 35448
rect 48832 35436 48838 35488
rect 1104 35386 78844 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 78844 35386
rect 1104 35312 78844 35334
rect 34698 35232 34704 35284
rect 34756 35232 34762 35284
rect 44726 35232 44732 35284
rect 44784 35272 44790 35284
rect 45189 35275 45247 35281
rect 45189 35272 45201 35275
rect 44784 35244 45201 35272
rect 44784 35232 44790 35244
rect 45189 35241 45201 35244
rect 45235 35272 45247 35275
rect 45833 35275 45891 35281
rect 45235 35244 45554 35272
rect 45235 35241 45247 35244
rect 45189 35235 45247 35241
rect 43714 35164 43720 35216
rect 43772 35204 43778 35216
rect 43772 35176 44956 35204
rect 43772 35164 43778 35176
rect 28445 35139 28503 35145
rect 28445 35105 28457 35139
rect 28491 35136 28503 35139
rect 28626 35136 28632 35148
rect 28491 35108 28632 35136
rect 28491 35105 28503 35108
rect 28445 35099 28503 35105
rect 28626 35096 28632 35108
rect 28684 35096 28690 35148
rect 28718 35096 28724 35148
rect 28776 35096 28782 35148
rect 31478 35096 31484 35148
rect 31536 35096 31542 35148
rect 36170 35096 36176 35148
rect 36228 35136 36234 35148
rect 36265 35139 36323 35145
rect 36265 35136 36277 35139
rect 36228 35108 36277 35136
rect 36228 35096 36234 35108
rect 36265 35105 36277 35108
rect 36311 35105 36323 35139
rect 44082 35136 44088 35148
rect 36265 35099 36323 35105
rect 43548 35108 44088 35136
rect 43548 35080 43576 35108
rect 44082 35096 44088 35108
rect 44140 35096 44146 35148
rect 28353 35071 28411 35077
rect 28353 35037 28365 35071
rect 28399 35068 28411 35071
rect 29549 35071 29607 35077
rect 29549 35068 29561 35071
rect 28399 35040 29561 35068
rect 28399 35037 28411 35040
rect 28353 35031 28411 35037
rect 29549 35037 29561 35040
rect 29595 35037 29607 35071
rect 29549 35031 29607 35037
rect 29914 35028 29920 35080
rect 29972 35068 29978 35080
rect 30101 35071 30159 35077
rect 30101 35068 30113 35071
rect 29972 35040 30113 35068
rect 29972 35028 29978 35040
rect 30101 35037 30113 35040
rect 30147 35037 30159 35071
rect 30101 35031 30159 35037
rect 30190 35028 30196 35080
rect 30248 35068 30254 35080
rect 31205 35071 31263 35077
rect 31205 35068 31217 35071
rect 30248 35040 31217 35068
rect 30248 35028 30254 35040
rect 31205 35037 31217 35040
rect 31251 35037 31263 35071
rect 31205 35031 31263 35037
rect 34977 35071 35035 35077
rect 34977 35037 34989 35071
rect 35023 35037 35035 35071
rect 34977 35031 35035 35037
rect 35161 35071 35219 35077
rect 35161 35037 35173 35071
rect 35207 35068 35219 35071
rect 35434 35068 35440 35080
rect 35207 35040 35440 35068
rect 35207 35037 35219 35040
rect 35161 35031 35219 35037
rect 31570 34960 31576 35012
rect 31628 35000 31634 35012
rect 34992 35000 35020 35031
rect 35434 35028 35440 35040
rect 35492 35028 35498 35080
rect 35529 35071 35587 35077
rect 35529 35037 35541 35071
rect 35575 35068 35587 35071
rect 36541 35071 36599 35077
rect 36541 35068 36553 35071
rect 35575 35040 36553 35068
rect 35575 35037 35587 35040
rect 35529 35031 35587 35037
rect 36541 35037 36553 35040
rect 36587 35068 36599 35071
rect 38562 35068 38568 35080
rect 36587 35040 38568 35068
rect 36587 35037 36599 35040
rect 36541 35031 36599 35037
rect 38562 35028 38568 35040
rect 38620 35028 38626 35080
rect 43346 35028 43352 35080
rect 43404 35028 43410 35080
rect 43530 35028 43536 35080
rect 43588 35028 43594 35080
rect 43625 35071 43683 35077
rect 43625 35037 43637 35071
rect 43671 35068 43683 35071
rect 43993 35071 44051 35077
rect 43993 35068 44005 35071
rect 43671 35040 44005 35068
rect 43671 35037 43683 35040
rect 43625 35031 43683 35037
rect 43993 35037 44005 35040
rect 44039 35037 44051 35071
rect 43993 35031 44051 35037
rect 44266 35028 44272 35080
rect 44324 35068 44330 35080
rect 44545 35071 44603 35077
rect 44545 35068 44557 35071
rect 44324 35040 44557 35068
rect 44324 35028 44330 35040
rect 44545 35037 44557 35040
rect 44591 35037 44603 35071
rect 44928 35068 44956 35176
rect 45526 35136 45554 35244
rect 45833 35241 45845 35275
rect 45879 35272 45891 35275
rect 46106 35272 46112 35284
rect 45879 35244 46112 35272
rect 45879 35241 45891 35244
rect 45833 35235 45891 35241
rect 46106 35232 46112 35244
rect 46164 35232 46170 35284
rect 46474 35136 46480 35148
rect 45526 35108 46480 35136
rect 46032 35077 46060 35108
rect 46474 35096 46480 35108
rect 46532 35096 46538 35148
rect 45649 35071 45707 35077
rect 45649 35068 45661 35071
rect 44928 35040 45661 35068
rect 44545 35031 44603 35037
rect 45649 35037 45661 35040
rect 45695 35037 45707 35071
rect 45649 35031 45707 35037
rect 46017 35071 46075 35077
rect 46017 35037 46029 35071
rect 46063 35037 46075 35071
rect 46017 35031 46075 35037
rect 46109 35071 46167 35077
rect 46109 35037 46121 35071
rect 46155 35068 46167 35071
rect 46842 35068 46848 35080
rect 46155 35040 46848 35068
rect 46155 35037 46167 35040
rect 46109 35031 46167 35037
rect 36262 35000 36268 35012
rect 31628 34972 31970 35000
rect 34992 34972 36268 35000
rect 31628 34960 31634 34972
rect 36262 34960 36268 34972
rect 36320 34960 36326 35012
rect 44634 34960 44640 35012
rect 44692 35000 44698 35012
rect 45373 35003 45431 35009
rect 45373 35000 45385 35003
rect 44692 34972 45385 35000
rect 44692 34960 44698 34972
rect 45373 34969 45385 34972
rect 45419 34969 45431 35003
rect 45373 34963 45431 34969
rect 2038 34892 2044 34944
rect 2096 34892 2102 34944
rect 32490 34892 32496 34944
rect 32548 34932 32554 34944
rect 32766 34932 32772 34944
rect 32548 34904 32772 34932
rect 32548 34892 32554 34904
rect 32766 34892 32772 34904
rect 32824 34932 32830 34944
rect 32953 34935 33011 34941
rect 32953 34932 32965 34935
rect 32824 34904 32965 34932
rect 32824 34892 32830 34904
rect 32953 34901 32965 34904
rect 32999 34901 33011 34935
rect 32953 34895 33011 34901
rect 34514 34892 34520 34944
rect 34572 34932 34578 34944
rect 34885 34935 34943 34941
rect 34885 34932 34897 34935
rect 34572 34904 34897 34932
rect 34572 34892 34578 34904
rect 34885 34901 34897 34904
rect 34931 34901 34943 34935
rect 34885 34895 34943 34901
rect 35250 34892 35256 34944
rect 35308 34932 35314 34944
rect 35437 34935 35495 34941
rect 35437 34932 35449 34935
rect 35308 34904 35449 34932
rect 35308 34892 35314 34904
rect 35437 34901 35449 34904
rect 35483 34932 35495 34935
rect 38746 34932 38752 34944
rect 35483 34904 38752 34932
rect 35483 34901 35495 34904
rect 35437 34895 35495 34901
rect 38746 34892 38752 34904
rect 38804 34892 38810 34944
rect 42794 34892 42800 34944
rect 42852 34932 42858 34944
rect 43165 34935 43223 34941
rect 43165 34932 43177 34935
rect 42852 34904 43177 34932
rect 42852 34892 42858 34904
rect 43165 34901 43177 34904
rect 43211 34901 43223 34935
rect 43165 34895 43223 34901
rect 44082 34892 44088 34944
rect 44140 34932 44146 34944
rect 45005 34935 45063 34941
rect 45005 34932 45017 34935
rect 44140 34904 45017 34932
rect 44140 34892 44146 34904
rect 45005 34901 45017 34904
rect 45051 34901 45063 34935
rect 45005 34895 45063 34901
rect 45173 34935 45231 34941
rect 45173 34901 45185 34935
rect 45219 34932 45231 34935
rect 45738 34932 45744 34944
rect 45219 34904 45744 34932
rect 45219 34901 45231 34904
rect 45173 34895 45231 34901
rect 45738 34892 45744 34904
rect 45796 34932 45802 34944
rect 46124 34932 46152 35031
rect 46842 35028 46848 35040
rect 46900 35028 46906 35080
rect 45796 34904 46152 34932
rect 45796 34892 45802 34904
rect 1104 34842 78844 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 66314 34842
rect 66366 34790 66378 34842
rect 66430 34790 66442 34842
rect 66494 34790 66506 34842
rect 66558 34790 66570 34842
rect 66622 34790 78844 34842
rect 1104 34768 78844 34790
rect 1302 34688 1308 34740
rect 1360 34728 1366 34740
rect 1857 34731 1915 34737
rect 1857 34728 1869 34731
rect 1360 34700 1869 34728
rect 1360 34688 1366 34700
rect 1857 34697 1869 34700
rect 1903 34697 1915 34731
rect 30190 34728 30196 34740
rect 1857 34691 1915 34697
rect 28460 34700 30196 34728
rect 2038 34552 2044 34604
rect 2096 34552 2102 34604
rect 28460 34601 28488 34700
rect 30190 34688 30196 34700
rect 30248 34688 30254 34740
rect 34606 34688 34612 34740
rect 34664 34728 34670 34740
rect 34664 34700 35112 34728
rect 34664 34688 34670 34700
rect 28718 34620 28724 34672
rect 28776 34620 28782 34672
rect 31570 34660 31576 34672
rect 29946 34646 31576 34660
rect 29932 34632 31576 34646
rect 28445 34595 28503 34601
rect 28445 34561 28457 34595
rect 28491 34561 28503 34595
rect 28445 34555 28503 34561
rect 2130 34484 2136 34536
rect 2188 34484 2194 34536
rect 29932 34524 29960 34632
rect 31570 34620 31576 34632
rect 31628 34620 31634 34672
rect 33870 34660 33876 34672
rect 33520 34632 33876 34660
rect 32214 34552 32220 34604
rect 32272 34592 32278 34604
rect 33520 34601 33548 34632
rect 33870 34620 33876 34632
rect 33928 34620 33934 34672
rect 35084 34660 35112 34700
rect 36170 34688 36176 34740
rect 36228 34688 36234 34740
rect 36262 34688 36268 34740
rect 36320 34688 36326 34740
rect 45103 34731 45161 34737
rect 41386 34700 42932 34728
rect 35250 34660 35256 34672
rect 35006 34632 35256 34660
rect 35250 34620 35256 34632
rect 35308 34620 35314 34672
rect 35342 34620 35348 34672
rect 35400 34620 35406 34672
rect 36188 34660 36216 34688
rect 36188 34632 39068 34660
rect 32401 34595 32459 34601
rect 32401 34592 32413 34595
rect 32272 34564 32413 34592
rect 32272 34552 32278 34564
rect 32401 34561 32413 34564
rect 32447 34561 32459 34595
rect 32401 34555 32459 34561
rect 33505 34595 33563 34601
rect 33505 34561 33517 34595
rect 33551 34561 33563 34595
rect 35360 34592 35388 34620
rect 35526 34592 35532 34604
rect 35360 34564 35532 34592
rect 33505 34555 33563 34561
rect 35526 34552 35532 34564
rect 35584 34592 35590 34604
rect 36173 34595 36231 34601
rect 36173 34592 36185 34595
rect 35584 34564 36185 34592
rect 35584 34552 35590 34564
rect 36173 34561 36185 34564
rect 36219 34561 36231 34595
rect 36173 34555 36231 34561
rect 36357 34595 36415 34601
rect 36357 34561 36369 34595
rect 36403 34561 36415 34595
rect 36357 34555 36415 34561
rect 37921 34595 37979 34601
rect 37921 34561 37933 34595
rect 37967 34592 37979 34595
rect 38194 34592 38200 34604
rect 37967 34564 38200 34592
rect 37967 34561 37979 34564
rect 37921 34555 37979 34561
rect 30837 34527 30895 34533
rect 30837 34524 30849 34527
rect 28552 34496 29960 34524
rect 30392 34496 30849 34524
rect 28350 34416 28356 34468
rect 28408 34456 28414 34468
rect 28552 34456 28580 34496
rect 28408 34428 28580 34456
rect 28408 34416 28414 34428
rect 29730 34416 29736 34468
rect 29788 34456 29794 34468
rect 30285 34459 30343 34465
rect 30285 34456 30297 34459
rect 29788 34428 30297 34456
rect 29788 34416 29794 34428
rect 30285 34425 30297 34428
rect 30331 34425 30343 34459
rect 30285 34419 30343 34425
rect 29914 34348 29920 34400
rect 29972 34388 29978 34400
rect 30193 34391 30251 34397
rect 30193 34388 30205 34391
rect 29972 34360 30205 34388
rect 29972 34348 29978 34360
rect 30193 34357 30205 34360
rect 30239 34388 30251 34391
rect 30392 34388 30420 34496
rect 30837 34493 30849 34496
rect 30883 34493 30895 34527
rect 30837 34487 30895 34493
rect 32306 34484 32312 34536
rect 32364 34484 32370 34536
rect 32490 34484 32496 34536
rect 32548 34484 32554 34536
rect 32582 34484 32588 34536
rect 32640 34484 32646 34536
rect 35253 34527 35311 34533
rect 35253 34493 35265 34527
rect 35299 34524 35311 34527
rect 35342 34524 35348 34536
rect 35299 34496 35348 34524
rect 35299 34493 35311 34496
rect 35253 34487 35311 34493
rect 35342 34484 35348 34496
rect 35400 34524 35406 34536
rect 35437 34527 35495 34533
rect 35437 34524 35449 34527
rect 35400 34496 35449 34524
rect 35400 34484 35406 34496
rect 35437 34493 35449 34496
rect 35483 34493 35495 34527
rect 35437 34487 35495 34493
rect 36081 34527 36139 34533
rect 36081 34493 36093 34527
rect 36127 34524 36139 34527
rect 36372 34524 36400 34555
rect 38194 34552 38200 34564
rect 38252 34552 38258 34604
rect 39040 34601 39068 34632
rect 39025 34595 39083 34601
rect 39025 34561 39037 34595
rect 39071 34561 39083 34595
rect 39025 34555 39083 34561
rect 40402 34552 40408 34604
rect 40460 34592 40466 34604
rect 41230 34592 41236 34604
rect 40460 34564 41236 34592
rect 40460 34552 40466 34564
rect 41230 34552 41236 34564
rect 41288 34592 41294 34604
rect 41386 34592 41414 34700
rect 42705 34663 42763 34669
rect 42705 34629 42717 34663
rect 42751 34660 42763 34663
rect 42794 34660 42800 34672
rect 42751 34632 42800 34660
rect 42751 34629 42763 34632
rect 42705 34623 42763 34629
rect 42794 34620 42800 34632
rect 42852 34620 42858 34672
rect 42904 34660 42932 34700
rect 45103 34697 45115 34731
rect 45149 34728 45161 34731
rect 45830 34728 45836 34740
rect 45149 34700 45836 34728
rect 45149 34697 45161 34700
rect 45103 34691 45161 34697
rect 45830 34688 45836 34700
rect 45888 34688 45894 34740
rect 42904 34632 43194 34660
rect 44634 34620 44640 34672
rect 44692 34660 44698 34672
rect 45189 34663 45247 34669
rect 45189 34660 45201 34663
rect 44692 34632 45201 34660
rect 44692 34620 44698 34632
rect 45189 34629 45201 34632
rect 45235 34629 45247 34663
rect 45189 34623 45247 34629
rect 41288 34564 41414 34592
rect 41288 34552 41294 34564
rect 42242 34552 42248 34604
rect 42300 34592 42306 34604
rect 42429 34595 42487 34601
rect 42429 34592 42441 34595
rect 42300 34564 42441 34592
rect 42300 34552 42306 34564
rect 42429 34561 42441 34564
rect 42475 34561 42487 34595
rect 42429 34555 42487 34561
rect 44266 34552 44272 34604
rect 44324 34592 44330 34604
rect 45005 34595 45063 34601
rect 45005 34592 45017 34595
rect 44324 34564 45017 34592
rect 44324 34552 44330 34564
rect 45005 34561 45017 34564
rect 45051 34561 45063 34595
rect 45005 34555 45063 34561
rect 45281 34595 45339 34601
rect 45281 34561 45293 34595
rect 45327 34592 45339 34595
rect 46106 34592 46112 34604
rect 45327 34564 46112 34592
rect 45327 34561 45339 34564
rect 45281 34555 45339 34561
rect 46106 34552 46112 34564
rect 46164 34552 46170 34604
rect 36127 34496 36400 34524
rect 36127 34493 36139 34496
rect 36081 34487 36139 34493
rect 30239 34360 30420 34388
rect 30239 34357 30251 34360
rect 30193 34351 30251 34357
rect 31938 34348 31944 34400
rect 31996 34388 32002 34400
rect 32125 34391 32183 34397
rect 32125 34388 32137 34391
rect 31996 34360 32137 34388
rect 31996 34348 32002 34360
rect 32125 34357 32137 34360
rect 32171 34357 32183 34391
rect 32125 34351 32183 34357
rect 33768 34391 33826 34397
rect 33768 34357 33780 34391
rect 33814 34388 33826 34391
rect 34514 34388 34520 34400
rect 33814 34360 34520 34388
rect 33814 34357 33826 34360
rect 33768 34351 33826 34357
rect 34514 34348 34520 34360
rect 34572 34348 34578 34400
rect 37274 34348 37280 34400
rect 37332 34348 37338 34400
rect 39288 34391 39346 34397
rect 39288 34357 39300 34391
rect 39334 34388 39346 34391
rect 39482 34388 39488 34400
rect 39334 34360 39488 34388
rect 39334 34357 39346 34360
rect 39288 34351 39346 34357
rect 39482 34348 39488 34360
rect 39540 34348 39546 34400
rect 40034 34348 40040 34400
rect 40092 34388 40098 34400
rect 40773 34391 40831 34397
rect 40773 34388 40785 34391
rect 40092 34360 40785 34388
rect 40092 34348 40098 34360
rect 40773 34357 40785 34360
rect 40819 34357 40831 34391
rect 40773 34351 40831 34357
rect 44177 34391 44235 34397
rect 44177 34357 44189 34391
rect 44223 34388 44235 34391
rect 44266 34388 44272 34400
rect 44223 34360 44272 34388
rect 44223 34357 44235 34360
rect 44177 34351 44235 34357
rect 44266 34348 44272 34360
rect 44324 34348 44330 34400
rect 1104 34298 78844 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 78844 34298
rect 1104 34224 78844 34246
rect 38105 34187 38163 34193
rect 38105 34153 38117 34187
rect 38151 34184 38163 34187
rect 38194 34184 38200 34196
rect 38151 34156 38200 34184
rect 38151 34153 38163 34156
rect 38105 34147 38163 34153
rect 38194 34144 38200 34156
rect 38252 34144 38258 34196
rect 39114 34144 39120 34196
rect 39172 34184 39178 34196
rect 39301 34187 39359 34193
rect 39301 34184 39313 34187
rect 39172 34156 39313 34184
rect 39172 34144 39178 34156
rect 39301 34153 39313 34156
rect 39347 34153 39359 34187
rect 39301 34147 39359 34153
rect 39482 34144 39488 34196
rect 39540 34144 39546 34196
rect 41138 34144 41144 34196
rect 41196 34184 41202 34196
rect 41325 34187 41383 34193
rect 41325 34184 41337 34187
rect 41196 34156 41337 34184
rect 41196 34144 41202 34156
rect 41325 34153 41337 34156
rect 41371 34153 41383 34187
rect 41325 34147 41383 34153
rect 43346 34144 43352 34196
rect 43404 34144 43410 34196
rect 934 34076 940 34128
rect 992 34116 998 34128
rect 1857 34119 1915 34125
rect 1857 34116 1869 34119
rect 992 34088 1869 34116
rect 992 34076 998 34088
rect 1857 34085 1869 34088
rect 1903 34085 1915 34119
rect 1857 34079 1915 34085
rect 28442 34076 28448 34128
rect 28500 34116 28506 34128
rect 29089 34119 29147 34125
rect 29089 34116 29101 34119
rect 28500 34088 29101 34116
rect 28500 34076 28506 34088
rect 29089 34085 29101 34088
rect 29135 34085 29147 34119
rect 35526 34116 35532 34128
rect 29089 34079 29147 34085
rect 34900 34088 35532 34116
rect 30190 34008 30196 34060
rect 30248 34008 30254 34060
rect 31941 34051 31999 34057
rect 31941 34017 31953 34051
rect 31987 34048 31999 34051
rect 32582 34048 32588 34060
rect 31987 34020 32588 34048
rect 31987 34017 31999 34020
rect 31941 34011 31999 34017
rect 2041 33983 2099 33989
rect 2041 33949 2053 33983
rect 2087 33980 2099 33983
rect 2130 33980 2136 33992
rect 2087 33952 2136 33980
rect 2087 33949 2099 33952
rect 2041 33943 2099 33949
rect 2130 33940 2136 33952
rect 2188 33940 2194 33992
rect 26970 33940 26976 33992
rect 27028 33940 27034 33992
rect 28350 33940 28356 33992
rect 28408 33940 28414 33992
rect 28626 33940 28632 33992
rect 28684 33980 28690 33992
rect 28813 33983 28871 33989
rect 28813 33980 28825 33983
rect 28684 33952 28825 33980
rect 28684 33940 28690 33952
rect 28813 33949 28825 33952
rect 28859 33949 28871 33983
rect 28813 33943 28871 33949
rect 28905 33983 28963 33989
rect 28905 33949 28917 33983
rect 28951 33980 28963 33983
rect 29730 33980 29736 33992
rect 28951 33952 29736 33980
rect 28951 33949 28963 33952
rect 28905 33943 28963 33949
rect 29730 33940 29736 33952
rect 29788 33940 29794 33992
rect 31570 33940 31576 33992
rect 31628 33940 31634 33992
rect 32214 33940 32220 33992
rect 32272 33980 32278 33992
rect 32416 33989 32444 34020
rect 32582 34008 32588 34020
rect 32640 34008 32646 34060
rect 34900 33989 34928 34088
rect 35526 34076 35532 34088
rect 35584 34076 35590 34128
rect 38562 34076 38568 34128
rect 38620 34116 38626 34128
rect 45094 34116 45100 34128
rect 38620 34088 45100 34116
rect 38620 34076 38626 34088
rect 45094 34076 45100 34088
rect 45152 34076 45158 34128
rect 35713 34051 35771 34057
rect 35713 34048 35725 34051
rect 35360 34020 35725 34048
rect 35360 33992 35388 34020
rect 35713 34017 35725 34020
rect 35759 34017 35771 34051
rect 35713 34011 35771 34017
rect 36265 34051 36323 34057
rect 36265 34017 36277 34051
rect 36311 34048 36323 34051
rect 37274 34048 37280 34060
rect 36311 34020 37280 34048
rect 36311 34017 36323 34020
rect 36265 34011 36323 34017
rect 37274 34008 37280 34020
rect 37332 34008 37338 34060
rect 40954 34008 40960 34060
rect 41012 34048 41018 34060
rect 43165 34051 43223 34057
rect 43165 34048 43177 34051
rect 41012 34020 43177 34048
rect 41012 34008 41018 34020
rect 43165 34017 43177 34020
rect 43211 34017 43223 34051
rect 43165 34011 43223 34017
rect 32309 33983 32367 33989
rect 32309 33980 32321 33983
rect 32272 33952 32321 33980
rect 32272 33940 32278 33952
rect 32309 33949 32321 33952
rect 32355 33949 32367 33983
rect 32309 33943 32367 33949
rect 32401 33983 32459 33989
rect 32401 33949 32413 33983
rect 32447 33949 32459 33983
rect 34885 33983 34943 33989
rect 32401 33943 32459 33949
rect 32508 33952 32996 33980
rect 27246 33872 27252 33924
rect 27304 33872 27310 33924
rect 29086 33872 29092 33924
rect 29144 33872 29150 33924
rect 30374 33872 30380 33924
rect 30432 33912 30438 33924
rect 30469 33915 30527 33921
rect 30469 33912 30481 33915
rect 30432 33884 30481 33912
rect 30432 33872 30438 33884
rect 30469 33881 30481 33884
rect 30515 33881 30527 33915
rect 32508 33912 32536 33952
rect 30469 33875 30527 33881
rect 32232 33884 32536 33912
rect 32585 33915 32643 33921
rect 28721 33847 28779 33853
rect 28721 33813 28733 33847
rect 28767 33844 28779 33847
rect 29454 33844 29460 33856
rect 28767 33816 29460 33844
rect 28767 33813 28779 33816
rect 28721 33807 28779 33813
rect 29454 33804 29460 33816
rect 29512 33804 29518 33856
rect 32030 33804 32036 33856
rect 32088 33804 32094 33856
rect 32232 33853 32260 33884
rect 32585 33881 32597 33915
rect 32631 33881 32643 33915
rect 32585 33875 32643 33881
rect 32217 33847 32275 33853
rect 32217 33813 32229 33847
rect 32263 33844 32275 33847
rect 32306 33844 32312 33856
rect 32263 33816 32312 33844
rect 32263 33813 32275 33816
rect 32217 33807 32275 33813
rect 32306 33804 32312 33816
rect 32364 33804 32370 33856
rect 32398 33804 32404 33856
rect 32456 33844 32462 33856
rect 32600 33844 32628 33875
rect 32456 33816 32628 33844
rect 32968 33844 32996 33952
rect 34885 33949 34897 33983
rect 34931 33949 34943 33983
rect 34885 33943 34943 33949
rect 35069 33983 35127 33989
rect 35069 33949 35081 33983
rect 35115 33980 35127 33983
rect 35342 33980 35348 33992
rect 35115 33952 35348 33980
rect 35115 33949 35127 33952
rect 35069 33943 35127 33949
rect 35342 33940 35348 33952
rect 35400 33940 35406 33992
rect 35526 33940 35532 33992
rect 35584 33940 35590 33992
rect 35989 33983 36047 33989
rect 35989 33949 36001 33983
rect 36035 33949 36047 33983
rect 35989 33943 36047 33949
rect 33042 33872 33048 33924
rect 33100 33912 33106 33924
rect 34977 33915 35035 33921
rect 34977 33912 34989 33915
rect 33100 33884 34989 33912
rect 33100 33872 33106 33884
rect 34977 33881 34989 33884
rect 35023 33881 35035 33915
rect 34977 33875 35035 33881
rect 35250 33872 35256 33924
rect 35308 33872 35314 33924
rect 33686 33844 33692 33856
rect 32968 33816 33692 33844
rect 32456 33804 32462 33816
rect 33686 33804 33692 33816
rect 33744 33844 33750 33856
rect 34701 33847 34759 33853
rect 34701 33844 34713 33847
rect 33744 33816 34713 33844
rect 33744 33804 33750 33816
rect 34701 33813 34713 33816
rect 34747 33813 34759 33847
rect 34701 33807 34759 33813
rect 35345 33847 35403 33853
rect 35345 33813 35357 33847
rect 35391 33844 35403 33847
rect 35434 33844 35440 33856
rect 35391 33816 35440 33844
rect 35391 33813 35403 33816
rect 35345 33807 35403 33813
rect 35434 33804 35440 33816
rect 35492 33804 35498 33856
rect 36004 33844 36032 33943
rect 36078 33940 36084 33992
rect 36136 33940 36142 33992
rect 36170 33940 36176 33992
rect 36228 33980 36234 33992
rect 36357 33983 36415 33989
rect 36357 33980 36369 33983
rect 36228 33952 36369 33980
rect 36228 33940 36234 33952
rect 36357 33949 36369 33952
rect 36403 33949 36415 33983
rect 36357 33943 36415 33949
rect 38930 33940 38936 33992
rect 38988 33940 38994 33992
rect 39942 33940 39948 33992
rect 40000 33980 40006 33992
rect 40221 33983 40279 33989
rect 40221 33980 40233 33983
rect 40000 33952 40233 33980
rect 40000 33940 40006 33952
rect 40221 33949 40233 33952
rect 40267 33949 40279 33983
rect 40221 33943 40279 33949
rect 40862 33940 40868 33992
rect 40920 33940 40926 33992
rect 41046 33940 41052 33992
rect 41104 33980 41110 33992
rect 41141 33983 41199 33989
rect 41141 33980 41153 33983
rect 41104 33952 41153 33980
rect 41104 33940 41110 33952
rect 41141 33949 41153 33952
rect 41187 33949 41199 33983
rect 41322 33980 41328 33992
rect 41141 33943 41199 33949
rect 41248 33952 41328 33980
rect 36265 33915 36323 33921
rect 36265 33881 36277 33915
rect 36311 33912 36323 33915
rect 36633 33915 36691 33921
rect 36633 33912 36645 33915
rect 36311 33884 36645 33912
rect 36311 33881 36323 33884
rect 36265 33875 36323 33881
rect 36633 33881 36645 33884
rect 36679 33881 36691 33915
rect 36633 33875 36691 33881
rect 37366 33872 37372 33924
rect 37424 33872 37430 33924
rect 39301 33915 39359 33921
rect 39301 33881 39313 33915
rect 39347 33912 39359 33915
rect 39853 33915 39911 33921
rect 39853 33912 39865 33915
rect 39347 33884 39865 33912
rect 39347 33881 39359 33884
rect 39301 33875 39359 33881
rect 39853 33881 39865 33884
rect 39899 33881 39911 33915
rect 39853 33875 39911 33881
rect 40034 33872 40040 33924
rect 40092 33912 40098 33924
rect 41248 33912 41276 33952
rect 41322 33940 41328 33952
rect 41380 33980 41386 33992
rect 42426 33980 42432 33992
rect 41380 33952 42432 33980
rect 41380 33940 41386 33952
rect 42426 33940 42432 33952
rect 42484 33940 42490 33992
rect 43530 33940 43536 33992
rect 43588 33980 43594 33992
rect 43625 33983 43683 33989
rect 43625 33980 43637 33983
rect 43588 33952 43637 33980
rect 43588 33940 43594 33952
rect 43625 33949 43637 33952
rect 43671 33949 43683 33983
rect 43625 33943 43683 33949
rect 42150 33912 42156 33924
rect 40092 33884 41276 33912
rect 41340 33884 42156 33912
rect 40092 33872 40098 33884
rect 36354 33844 36360 33856
rect 36004 33816 36360 33844
rect 36354 33804 36360 33816
rect 36412 33804 36418 33856
rect 40678 33804 40684 33856
rect 40736 33844 40742 33856
rect 40957 33847 41015 33853
rect 40957 33844 40969 33847
rect 40736 33816 40969 33844
rect 40736 33804 40742 33816
rect 40957 33813 40969 33816
rect 41003 33844 41015 33847
rect 41340 33844 41368 33884
rect 42150 33872 42156 33884
rect 42208 33872 42214 33924
rect 41003 33816 41368 33844
rect 43533 33847 43591 33853
rect 41003 33813 41015 33816
rect 40957 33807 41015 33813
rect 43533 33813 43545 33847
rect 43579 33844 43591 33847
rect 44266 33844 44272 33856
rect 43579 33816 44272 33844
rect 43579 33813 43591 33816
rect 43533 33807 43591 33813
rect 44266 33804 44272 33816
rect 44324 33804 44330 33856
rect 45094 33804 45100 33856
rect 45152 33804 45158 33856
rect 1104 33754 78844 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 66314 33754
rect 66366 33702 66378 33754
rect 66430 33702 66442 33754
rect 66494 33702 66506 33754
rect 66558 33702 66570 33754
rect 66622 33702 78844 33754
rect 1104 33680 78844 33702
rect 27246 33600 27252 33652
rect 27304 33640 27310 33652
rect 28353 33643 28411 33649
rect 28353 33640 28365 33643
rect 27304 33612 28365 33640
rect 27304 33600 27310 33612
rect 28353 33609 28365 33612
rect 28399 33609 28411 33643
rect 28353 33603 28411 33609
rect 28813 33643 28871 33649
rect 28813 33609 28825 33643
rect 28859 33640 28871 33643
rect 29086 33640 29092 33652
rect 28859 33612 29092 33640
rect 28859 33609 28871 33612
rect 28813 33603 28871 33609
rect 29086 33600 29092 33612
rect 29144 33600 29150 33652
rect 29549 33643 29607 33649
rect 29549 33609 29561 33643
rect 29595 33609 29607 33643
rect 29549 33603 29607 33609
rect 28994 33572 29000 33584
rect 28276 33544 29000 33572
rect 28276 33513 28304 33544
rect 28994 33532 29000 33544
rect 29052 33572 29058 33584
rect 29564 33572 29592 33603
rect 30374 33600 30380 33652
rect 30432 33600 30438 33652
rect 38930 33600 38936 33652
rect 38988 33600 38994 33652
rect 39942 33600 39948 33652
rect 40000 33640 40006 33652
rect 40313 33643 40371 33649
rect 40313 33640 40325 33643
rect 40000 33612 40325 33640
rect 40000 33600 40006 33612
rect 40313 33609 40325 33612
rect 40359 33609 40371 33643
rect 40313 33603 40371 33609
rect 40481 33643 40539 33649
rect 40481 33609 40493 33643
rect 40527 33640 40539 33643
rect 40862 33640 40868 33652
rect 40527 33612 40868 33640
rect 40527 33609 40539 33612
rect 40481 33603 40539 33609
rect 29712 33575 29770 33581
rect 29712 33572 29724 33575
rect 29052 33544 29592 33572
rect 29656 33544 29724 33572
rect 29052 33532 29058 33544
rect 2041 33507 2099 33513
rect 2041 33473 2053 33507
rect 2087 33504 2099 33507
rect 2133 33507 2191 33513
rect 2133 33504 2145 33507
rect 2087 33476 2145 33504
rect 2087 33473 2099 33476
rect 2041 33467 2099 33473
rect 2133 33473 2145 33476
rect 2179 33473 2191 33507
rect 2133 33467 2191 33473
rect 28261 33507 28319 33513
rect 28261 33473 28273 33507
rect 28307 33473 28319 33507
rect 28261 33467 28319 33473
rect 28442 33464 28448 33516
rect 28500 33464 28506 33516
rect 28626 33464 28632 33516
rect 28684 33504 28690 33516
rect 29656 33504 29684 33544
rect 29712 33541 29724 33544
rect 29758 33541 29770 33575
rect 29712 33535 29770 33541
rect 29914 33532 29920 33584
rect 29972 33532 29978 33584
rect 32214 33532 32220 33584
rect 32272 33572 32278 33584
rect 32769 33575 32827 33581
rect 32769 33572 32781 33575
rect 32272 33544 32781 33572
rect 32272 33532 32278 33544
rect 32769 33541 32781 33544
rect 32815 33541 32827 33575
rect 32769 33535 32827 33541
rect 35250 33532 35256 33584
rect 35308 33572 35314 33584
rect 38948 33572 38976 33600
rect 35308 33544 35664 33572
rect 35308 33532 35314 33544
rect 30837 33507 30895 33513
rect 30837 33504 30849 33507
rect 28684 33476 30849 33504
rect 28684 33464 28690 33476
rect 30837 33473 30849 33476
rect 30883 33504 30895 33507
rect 32030 33504 32036 33516
rect 30883 33476 32036 33504
rect 30883 33473 30895 33476
rect 30837 33467 30895 33473
rect 32030 33464 32036 33476
rect 32088 33464 32094 33516
rect 32309 33507 32367 33513
rect 32309 33473 32321 33507
rect 32355 33504 32367 33507
rect 32398 33504 32404 33516
rect 32355 33476 32404 33504
rect 32355 33473 32367 33476
rect 32309 33467 32367 33473
rect 32398 33464 32404 33476
rect 32456 33464 32462 33516
rect 32493 33507 32551 33513
rect 32493 33473 32505 33507
rect 32539 33504 32551 33507
rect 32582 33504 32588 33516
rect 32539 33476 32588 33504
rect 32539 33473 32551 33476
rect 32493 33467 32551 33473
rect 32582 33464 32588 33476
rect 32640 33464 32646 33516
rect 35434 33464 35440 33516
rect 35492 33464 35498 33516
rect 35636 33513 35664 33544
rect 38396 33544 38976 33572
rect 35621 33507 35679 33513
rect 35621 33473 35633 33507
rect 35667 33504 35679 33507
rect 35986 33504 35992 33516
rect 35667 33476 35992 33504
rect 35667 33473 35679 33476
rect 35621 33467 35679 33473
rect 35986 33464 35992 33476
rect 36044 33464 36050 33516
rect 36354 33464 36360 33516
rect 36412 33464 36418 33516
rect 36541 33507 36599 33513
rect 36541 33473 36553 33507
rect 36587 33504 36599 33507
rect 36998 33504 37004 33516
rect 36587 33476 37004 33504
rect 36587 33473 36599 33476
rect 36541 33467 36599 33473
rect 29454 33396 29460 33448
rect 29512 33396 29518 33448
rect 35529 33439 35587 33445
rect 35529 33405 35541 33439
rect 35575 33436 35587 33439
rect 36078 33436 36084 33448
rect 35575 33408 36084 33436
rect 35575 33405 35587 33408
rect 35529 33399 35587 33405
rect 36078 33396 36084 33408
rect 36136 33436 36142 33448
rect 36556 33436 36584 33467
rect 36998 33464 37004 33476
rect 37056 33464 37062 33516
rect 38102 33464 38108 33516
rect 38160 33464 38166 33516
rect 38396 33513 38424 33544
rect 39482 33532 39488 33584
rect 39540 33572 39546 33584
rect 39821 33575 39879 33581
rect 39821 33572 39833 33575
rect 39540 33544 39833 33572
rect 39540 33532 39546 33544
rect 39821 33541 39833 33544
rect 39867 33572 39879 33575
rect 39960 33572 39988 33600
rect 39867 33544 39988 33572
rect 40037 33575 40095 33581
rect 39867 33541 39879 33544
rect 39821 33535 39879 33541
rect 40037 33541 40049 33575
rect 40083 33572 40095 33575
rect 40083 33544 40172 33572
rect 40083 33541 40095 33544
rect 40037 33535 40095 33541
rect 38381 33507 38439 33513
rect 38381 33473 38393 33507
rect 38427 33473 38439 33507
rect 38381 33467 38439 33473
rect 38565 33507 38623 33513
rect 38565 33473 38577 33507
rect 38611 33504 38623 33507
rect 38933 33507 38991 33513
rect 38933 33504 38945 33507
rect 38611 33476 38945 33504
rect 38611 33473 38623 33476
rect 38565 33467 38623 33473
rect 38933 33473 38945 33476
rect 38979 33473 38991 33507
rect 38933 33467 38991 33473
rect 36136 33408 36584 33436
rect 36136 33396 36142 33408
rect 39206 33396 39212 33448
rect 39264 33436 39270 33448
rect 39577 33439 39635 33445
rect 39577 33436 39589 33439
rect 39264 33408 39589 33436
rect 39264 33396 39270 33408
rect 39577 33405 39589 33408
rect 39623 33436 39635 33439
rect 40144 33436 40172 33544
rect 40328 33504 40356 33603
rect 40862 33600 40868 33612
rect 40920 33600 40926 33652
rect 41046 33640 41052 33652
rect 40972 33612 41052 33640
rect 40678 33532 40684 33584
rect 40736 33572 40742 33584
rect 40972 33572 41000 33612
rect 41046 33600 41052 33612
rect 41104 33640 41110 33652
rect 41969 33643 42027 33649
rect 41104 33612 41414 33640
rect 41104 33600 41110 33612
rect 40736 33544 41000 33572
rect 41141 33575 41199 33581
rect 40736 33532 40742 33544
rect 41141 33541 41153 33575
rect 41187 33541 41199 33575
rect 41386 33572 41414 33612
rect 41969 33609 41981 33643
rect 42015 33640 42027 33643
rect 43806 33640 43812 33652
rect 42015 33612 43812 33640
rect 42015 33609 42027 33612
rect 41969 33603 42027 33609
rect 43806 33600 43812 33612
rect 43864 33600 43870 33652
rect 44174 33600 44180 33652
rect 44232 33640 44238 33652
rect 44453 33643 44511 33649
rect 44453 33640 44465 33643
rect 44232 33612 44465 33640
rect 44232 33600 44238 33612
rect 44453 33609 44465 33612
rect 44499 33609 44511 33643
rect 45922 33640 45928 33652
rect 44453 33603 44511 33609
rect 44652 33612 45928 33640
rect 41386 33544 42748 33572
rect 41141 33535 41199 33541
rect 40773 33507 40831 33513
rect 40773 33504 40785 33507
rect 40328 33476 40785 33504
rect 40773 33473 40785 33476
rect 40819 33473 40831 33507
rect 40773 33467 40831 33473
rect 40954 33464 40960 33516
rect 41012 33504 41018 33516
rect 41156 33504 41184 33535
rect 41012 33476 41184 33504
rect 41012 33464 41018 33476
rect 41322 33464 41328 33516
rect 41380 33504 41386 33516
rect 41509 33507 41567 33513
rect 41509 33504 41521 33507
rect 41380 33476 41521 33504
rect 41380 33464 41386 33476
rect 41509 33473 41521 33476
rect 41555 33473 41567 33507
rect 41509 33467 41567 33473
rect 41785 33510 41843 33513
rect 41892 33510 41920 33544
rect 41785 33507 41920 33510
rect 41785 33473 41797 33507
rect 41831 33482 41920 33507
rect 41831 33473 41843 33482
rect 41785 33467 41843 33473
rect 42150 33464 42156 33516
rect 42208 33464 42214 33516
rect 42426 33464 42432 33516
rect 42484 33464 42490 33516
rect 42720 33513 42748 33544
rect 42705 33507 42763 33513
rect 42705 33473 42717 33507
rect 42751 33473 42763 33507
rect 42705 33467 42763 33473
rect 44266 33464 44272 33516
rect 44324 33464 44330 33516
rect 44652 33513 44680 33612
rect 45922 33600 45928 33612
rect 45980 33600 45986 33652
rect 46106 33600 46112 33652
rect 46164 33600 46170 33652
rect 46198 33600 46204 33652
rect 46256 33640 46262 33652
rect 46256 33612 46612 33640
rect 46256 33600 46262 33612
rect 45094 33532 45100 33584
rect 45152 33532 45158 33584
rect 46584 33572 46612 33612
rect 47670 33572 47676 33584
rect 45526 33544 46336 33572
rect 44637 33507 44695 33513
rect 44637 33473 44649 33507
rect 44683 33473 44695 33507
rect 44637 33467 44695 33473
rect 44726 33464 44732 33516
rect 44784 33504 44790 33516
rect 44821 33507 44879 33513
rect 44821 33504 44833 33507
rect 44784 33476 44833 33504
rect 44784 33464 44790 33476
rect 44821 33473 44833 33476
rect 44867 33473 44879 33507
rect 44821 33467 44879 33473
rect 42521 33439 42579 33445
rect 42521 33436 42533 33439
rect 39623 33408 42533 33436
rect 39623 33405 39635 33408
rect 39577 33399 39635 33405
rect 934 33328 940 33380
rect 992 33368 998 33380
rect 1857 33371 1915 33377
rect 1857 33368 1869 33371
rect 992 33340 1869 33368
rect 992 33328 998 33340
rect 1857 33337 1869 33340
rect 1903 33337 1915 33371
rect 1857 33331 1915 33337
rect 29472 33300 29500 33396
rect 30561 33371 30619 33377
rect 30561 33337 30573 33371
rect 30607 33368 30619 33371
rect 31938 33368 31944 33380
rect 30607 33340 31944 33368
rect 30607 33337 30619 33340
rect 30561 33331 30619 33337
rect 31938 33328 31944 33340
rect 31996 33328 32002 33380
rect 41325 33371 41383 33377
rect 41325 33337 41337 33371
rect 41371 33368 41383 33371
rect 41598 33368 41604 33380
rect 41371 33340 41604 33368
rect 41371 33337 41383 33340
rect 41325 33331 41383 33337
rect 41598 33328 41604 33340
rect 41656 33328 41662 33380
rect 29730 33300 29736 33312
rect 29472 33272 29736 33300
rect 29730 33260 29736 33272
rect 29788 33260 29794 33312
rect 32030 33260 32036 33312
rect 32088 33300 32094 33312
rect 32125 33303 32183 33309
rect 32125 33300 32137 33303
rect 32088 33272 32137 33300
rect 32088 33260 32094 33272
rect 32125 33269 32137 33272
rect 32171 33269 32183 33303
rect 32125 33263 32183 33269
rect 32677 33303 32735 33309
rect 32677 33269 32689 33303
rect 32723 33300 32735 33303
rect 33042 33300 33048 33312
rect 32723 33272 33048 33300
rect 32723 33269 32735 33272
rect 32677 33263 32735 33269
rect 33042 33260 33048 33272
rect 33100 33260 33106 33312
rect 36541 33303 36599 33309
rect 36541 33269 36553 33303
rect 36587 33300 36599 33303
rect 37274 33300 37280 33312
rect 36587 33272 37280 33300
rect 36587 33269 36599 33272
rect 36541 33263 36599 33269
rect 37274 33260 37280 33272
rect 37332 33260 37338 33312
rect 37734 33260 37740 33312
rect 37792 33300 37798 33312
rect 37921 33303 37979 33309
rect 37921 33300 37933 33303
rect 37792 33272 37933 33300
rect 37792 33260 37798 33272
rect 37921 33269 37933 33272
rect 37967 33269 37979 33303
rect 37921 33263 37979 33269
rect 39666 33260 39672 33312
rect 39724 33260 39730 33312
rect 39850 33260 39856 33312
rect 39908 33260 39914 33312
rect 40497 33303 40555 33309
rect 40497 33269 40509 33303
rect 40543 33300 40555 33303
rect 40586 33300 40592 33312
rect 40543 33272 40592 33300
rect 40543 33269 40555 33272
rect 40497 33263 40555 33269
rect 40586 33260 40592 33272
rect 40644 33260 40650 33312
rect 41138 33260 41144 33312
rect 41196 33260 41202 33312
rect 41785 33303 41843 33309
rect 41785 33269 41797 33303
rect 41831 33300 41843 33303
rect 41892 33300 41920 33408
rect 42521 33405 42533 33408
rect 42567 33405 42579 33439
rect 45526 33436 45554 33544
rect 46308 33513 46336 33544
rect 46584 33544 47676 33572
rect 46293 33507 46351 33513
rect 46293 33473 46305 33507
rect 46339 33473 46351 33507
rect 46293 33467 46351 33473
rect 46382 33464 46388 33516
rect 46440 33464 46446 33516
rect 46584 33513 46612 33544
rect 47670 33532 47676 33544
rect 47728 33532 47734 33584
rect 48774 33532 48780 33584
rect 48832 33532 48838 33584
rect 46569 33507 46627 33513
rect 46569 33473 46581 33507
rect 46615 33473 46627 33507
rect 46569 33467 46627 33473
rect 46661 33507 46719 33513
rect 46661 33473 46673 33507
rect 46707 33473 46719 33507
rect 46661 33467 46719 33473
rect 42521 33399 42579 33405
rect 42904 33408 45554 33436
rect 45925 33439 45983 33445
rect 42904 33377 42932 33408
rect 45925 33405 45937 33439
rect 45971 33436 45983 33439
rect 46014 33436 46020 33448
rect 45971 33408 46020 33436
rect 45971 33405 45983 33408
rect 45925 33399 45983 33405
rect 46014 33396 46020 33408
rect 46072 33396 46078 33448
rect 46676 33436 46704 33467
rect 46842 33464 46848 33516
rect 46900 33504 46906 33516
rect 46937 33507 46995 33513
rect 46937 33504 46949 33507
rect 46900 33476 46949 33504
rect 46900 33464 46906 33476
rect 46937 33473 46949 33476
rect 46983 33473 46995 33507
rect 46937 33467 46995 33473
rect 46124 33408 46704 33436
rect 42889 33371 42947 33377
rect 42889 33337 42901 33371
rect 42935 33337 42947 33371
rect 42889 33331 42947 33337
rect 44726 33328 44732 33380
rect 44784 33368 44790 33380
rect 45186 33368 45192 33380
rect 44784 33340 45192 33368
rect 44784 33328 44790 33340
rect 45186 33328 45192 33340
rect 45244 33368 45250 33380
rect 46124 33368 46152 33408
rect 47762 33396 47768 33448
rect 47820 33396 47826 33448
rect 48038 33396 48044 33448
rect 48096 33396 48102 33448
rect 47780 33368 47808 33396
rect 45244 33340 46152 33368
rect 46860 33340 47808 33368
rect 45244 33328 45250 33340
rect 41831 33272 41920 33300
rect 41831 33269 41843 33272
rect 41785 33263 41843 33269
rect 42150 33260 42156 33312
rect 42208 33300 42214 33312
rect 42429 33303 42487 33309
rect 42429 33300 42441 33303
rect 42208 33272 42441 33300
rect 42208 33260 42214 33272
rect 42429 33269 42441 33272
rect 42475 33269 42487 33303
rect 42429 33263 42487 33269
rect 44634 33260 44640 33312
rect 44692 33260 44698 33312
rect 46014 33260 46020 33312
rect 46072 33300 46078 33312
rect 46860 33300 46888 33340
rect 46072 33272 46888 33300
rect 47029 33303 47087 33309
rect 46072 33260 46078 33272
rect 47029 33269 47041 33303
rect 47075 33300 47087 33303
rect 47486 33300 47492 33312
rect 47075 33272 47492 33300
rect 47075 33269 47087 33272
rect 47029 33263 47087 33269
rect 47486 33260 47492 33272
rect 47544 33260 47550 33312
rect 47670 33260 47676 33312
rect 47728 33300 47734 33312
rect 49513 33303 49571 33309
rect 49513 33300 49525 33303
rect 47728 33272 49525 33300
rect 47728 33260 47734 33272
rect 49513 33269 49525 33272
rect 49559 33269 49571 33303
rect 49513 33263 49571 33269
rect 49602 33260 49608 33312
rect 49660 33300 49666 33312
rect 49697 33303 49755 33309
rect 49697 33300 49709 33303
rect 49660 33272 49709 33300
rect 49660 33260 49666 33272
rect 49697 33269 49709 33272
rect 49743 33269 49755 33303
rect 49697 33263 49755 33269
rect 1104 33210 78844 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 78844 33210
rect 1104 33136 78844 33158
rect 30282 33056 30288 33108
rect 30340 33096 30346 33108
rect 32033 33099 32091 33105
rect 32033 33096 32045 33099
rect 30340 33068 32045 33096
rect 30340 33056 30346 33068
rect 32033 33065 32045 33068
rect 32079 33065 32091 33099
rect 32033 33059 32091 33065
rect 33689 33099 33747 33105
rect 33689 33065 33701 33099
rect 33735 33096 33747 33099
rect 33962 33096 33968 33108
rect 33735 33068 33968 33096
rect 33735 33065 33747 33068
rect 33689 33059 33747 33065
rect 33962 33056 33968 33068
rect 34020 33056 34026 33108
rect 36354 33096 36360 33108
rect 35544 33068 36360 33096
rect 32401 33031 32459 33037
rect 32401 32997 32413 33031
rect 32447 33028 32459 33031
rect 35544 33028 35572 33068
rect 36354 33056 36360 33068
rect 36412 33096 36418 33108
rect 36906 33096 36912 33108
rect 36412 33068 36912 33096
rect 36412 33056 36418 33068
rect 36906 33056 36912 33068
rect 36964 33056 36970 33108
rect 36998 33056 37004 33108
rect 37056 33056 37062 33108
rect 37369 33099 37427 33105
rect 37369 33065 37381 33099
rect 37415 33096 37427 33099
rect 38102 33096 38108 33108
rect 37415 33068 38108 33096
rect 37415 33065 37427 33068
rect 37369 33059 37427 33065
rect 38102 33056 38108 33068
rect 38160 33056 38166 33108
rect 38930 33056 38936 33108
rect 38988 33096 38994 33108
rect 39301 33099 39359 33105
rect 39301 33096 39313 33099
rect 38988 33068 39313 33096
rect 38988 33056 38994 33068
rect 39301 33065 39313 33068
rect 39347 33065 39359 33099
rect 39301 33059 39359 33065
rect 40678 33056 40684 33108
rect 40736 33096 40742 33108
rect 40865 33099 40923 33105
rect 40865 33096 40877 33099
rect 40736 33068 40877 33096
rect 40736 33056 40742 33068
rect 40865 33065 40877 33068
rect 40911 33065 40923 33099
rect 40865 33059 40923 33065
rect 43806 33056 43812 33108
rect 43864 33056 43870 33108
rect 44266 33056 44272 33108
rect 44324 33096 44330 33108
rect 44324 33068 45140 33096
rect 44324 33056 44330 33068
rect 37016 33028 37044 33056
rect 32447 33000 35572 33028
rect 32447 32997 32459 33000
rect 32401 32991 32459 32997
rect 28994 32960 29000 32972
rect 28276 32932 29000 32960
rect 28276 32901 28304 32932
rect 28994 32920 29000 32932
rect 29052 32920 29058 32972
rect 30190 32920 30196 32972
rect 30248 32960 30254 32972
rect 30285 32963 30343 32969
rect 30285 32960 30297 32963
rect 30248 32932 30297 32960
rect 30248 32920 30254 32932
rect 30285 32929 30297 32932
rect 30331 32929 30343 32963
rect 30285 32923 30343 32929
rect 33042 32920 33048 32972
rect 33100 32920 33106 32972
rect 33597 32963 33655 32969
rect 33597 32929 33609 32963
rect 33643 32960 33655 32963
rect 33643 32932 34100 32960
rect 33643 32929 33655 32932
rect 33597 32923 33655 32929
rect 2041 32895 2099 32901
rect 2041 32861 2053 32895
rect 2087 32892 2099 32895
rect 2133 32895 2191 32901
rect 2133 32892 2145 32895
rect 2087 32864 2145 32892
rect 2087 32861 2099 32864
rect 2041 32855 2099 32861
rect 2133 32861 2145 32864
rect 2179 32861 2191 32895
rect 2133 32855 2191 32861
rect 28261 32895 28319 32901
rect 28261 32861 28273 32895
rect 28307 32861 28319 32895
rect 28261 32855 28319 32861
rect 28445 32895 28503 32901
rect 28445 32861 28457 32895
rect 28491 32892 28503 32895
rect 28629 32895 28687 32901
rect 28629 32892 28641 32895
rect 28491 32864 28641 32892
rect 28491 32861 28503 32864
rect 28445 32855 28503 32861
rect 28629 32861 28641 32864
rect 28675 32861 28687 32895
rect 28629 32855 28687 32861
rect 29178 32852 29184 32904
rect 29236 32852 29242 32904
rect 32030 32852 32036 32904
rect 32088 32852 32094 32904
rect 32122 32852 32128 32904
rect 32180 32852 32186 32904
rect 33686 32852 33692 32904
rect 33744 32852 33750 32904
rect 34072 32901 34100 32932
rect 33965 32895 34023 32901
rect 33965 32861 33977 32895
rect 34011 32861 34023 32895
rect 33965 32855 34023 32861
rect 34057 32895 34115 32901
rect 34057 32861 34069 32895
rect 34103 32861 34115 32895
rect 35544 32892 35572 33000
rect 36096 33000 37044 33028
rect 35651 32895 35709 32901
rect 35651 32892 35663 32895
rect 35544 32864 35663 32892
rect 34057 32855 34115 32861
rect 35651 32861 35663 32864
rect 35697 32861 35709 32895
rect 35651 32855 35709 32861
rect 35805 32895 35863 32901
rect 35805 32861 35817 32895
rect 35851 32892 35863 32895
rect 36096 32892 36124 33000
rect 39206 32988 39212 33040
rect 39264 32988 39270 33040
rect 45005 33031 45063 33037
rect 45005 33028 45017 33031
rect 44100 33000 45017 33028
rect 36170 32920 36176 32972
rect 36228 32960 36234 32972
rect 37461 32963 37519 32969
rect 37461 32960 37473 32963
rect 36228 32932 37473 32960
rect 36228 32920 36234 32932
rect 37461 32929 37473 32932
rect 37507 32929 37519 32963
rect 37461 32923 37519 32929
rect 37734 32920 37740 32972
rect 37792 32920 37798 32972
rect 38746 32920 38752 32972
rect 38804 32960 38810 32972
rect 39669 32963 39727 32969
rect 38804 32932 39620 32960
rect 38804 32920 38810 32932
rect 35851 32864 36124 32892
rect 37001 32895 37059 32901
rect 35851 32861 35863 32864
rect 35805 32855 35863 32861
rect 37001 32861 37013 32895
rect 37047 32861 37059 32895
rect 37001 32855 37059 32861
rect 29362 32784 29368 32836
rect 29420 32824 29426 32836
rect 29549 32827 29607 32833
rect 29549 32824 29561 32827
rect 29420 32796 29561 32824
rect 29420 32784 29426 32796
rect 29549 32793 29561 32796
rect 29595 32793 29607 32827
rect 33980 32824 34008 32855
rect 33980 32796 35388 32824
rect 29549 32787 29607 32793
rect 35360 32768 35388 32796
rect 934 32716 940 32768
rect 992 32756 998 32768
rect 1857 32759 1915 32765
rect 1857 32756 1869 32759
rect 992 32728 1869 32756
rect 992 32716 998 32728
rect 1857 32725 1869 32728
rect 1903 32725 1915 32759
rect 1857 32719 1915 32725
rect 27982 32716 27988 32768
rect 28040 32756 28046 32768
rect 28353 32759 28411 32765
rect 28353 32756 28365 32759
rect 28040 32728 28365 32756
rect 28040 32716 28046 32728
rect 28353 32725 28365 32728
rect 28399 32725 28411 32759
rect 28353 32719 28411 32725
rect 33873 32759 33931 32765
rect 33873 32725 33885 32759
rect 33919 32756 33931 32759
rect 34149 32759 34207 32765
rect 34149 32756 34161 32759
rect 33919 32728 34161 32756
rect 33919 32725 33931 32728
rect 33873 32719 33931 32725
rect 34149 32725 34161 32728
rect 34195 32725 34207 32759
rect 34149 32719 34207 32725
rect 35342 32716 35348 32768
rect 35400 32756 35406 32768
rect 35437 32759 35495 32765
rect 35437 32756 35449 32759
rect 35400 32728 35449 32756
rect 35400 32716 35406 32728
rect 35437 32725 35449 32728
rect 35483 32725 35495 32759
rect 37016 32756 37044 32855
rect 37090 32852 37096 32904
rect 37148 32852 37154 32904
rect 38856 32878 38884 32932
rect 39482 32852 39488 32904
rect 39540 32852 39546 32904
rect 39592 32892 39620 32932
rect 39669 32929 39681 32963
rect 39715 32960 39727 32963
rect 39850 32960 39856 32972
rect 39715 32932 39856 32960
rect 39715 32929 39727 32932
rect 39669 32923 39727 32929
rect 39850 32920 39856 32932
rect 39908 32920 39914 32972
rect 42242 32920 42248 32972
rect 42300 32960 42306 32972
rect 42613 32963 42671 32969
rect 42613 32960 42625 32963
rect 42300 32932 42625 32960
rect 42300 32920 42306 32932
rect 42613 32929 42625 32932
rect 42659 32960 42671 32963
rect 42702 32960 42708 32972
rect 42659 32932 42708 32960
rect 42659 32929 42671 32932
rect 42613 32923 42671 32929
rect 42702 32920 42708 32932
rect 42760 32920 42766 32972
rect 44100 32969 44128 33000
rect 45005 32997 45017 33000
rect 45051 32997 45063 33031
rect 45112 33028 45140 33068
rect 45186 33056 45192 33108
rect 45244 33056 45250 33108
rect 46569 33099 46627 33105
rect 46569 33096 46581 33099
rect 45526 33068 46581 33096
rect 45370 33028 45376 33040
rect 45112 33000 45376 33028
rect 45005 32991 45063 32997
rect 45370 32988 45376 33000
rect 45428 32988 45434 33040
rect 44085 32963 44143 32969
rect 44085 32929 44097 32963
rect 44131 32929 44143 32963
rect 45186 32960 45192 32972
rect 44085 32923 44143 32929
rect 44652 32932 45192 32960
rect 39592 32864 39988 32892
rect 39040 32796 39712 32824
rect 39040 32756 39068 32796
rect 39684 32768 39712 32796
rect 39960 32768 39988 32864
rect 41230 32852 41236 32904
rect 41288 32852 41294 32904
rect 44177 32895 44235 32901
rect 44177 32861 44189 32895
rect 44223 32892 44235 32895
rect 44542 32892 44548 32904
rect 44223 32864 44548 32892
rect 44223 32861 44235 32864
rect 44177 32855 44235 32861
rect 44542 32852 44548 32864
rect 44600 32852 44606 32904
rect 44652 32901 44680 32932
rect 45186 32920 45192 32932
rect 45244 32960 45250 32972
rect 45526 32960 45554 33068
rect 46569 33065 46581 33068
rect 46615 33065 46627 33099
rect 46569 33059 46627 33065
rect 47949 33099 48007 33105
rect 47949 33065 47961 33099
rect 47995 33096 48007 33099
rect 48038 33096 48044 33108
rect 47995 33068 48044 33096
rect 47995 33065 48007 33068
rect 47949 33059 48007 33065
rect 48038 33056 48044 33068
rect 48096 33056 48102 33108
rect 46385 33031 46443 33037
rect 46385 32997 46397 33031
rect 46431 33028 46443 33031
rect 46842 33028 46848 33040
rect 46431 33000 46848 33028
rect 46431 32997 46443 33000
rect 46385 32991 46443 32997
rect 46842 32988 46848 33000
rect 46900 32988 46906 33040
rect 45244 32932 45554 32960
rect 45244 32920 45250 32932
rect 45922 32920 45928 32972
rect 45980 32960 45986 32972
rect 46293 32963 46351 32969
rect 46293 32960 46305 32963
rect 45980 32932 46305 32960
rect 45980 32920 45986 32932
rect 46293 32929 46305 32932
rect 46339 32929 46351 32963
rect 46293 32923 46351 32929
rect 47044 32932 47624 32960
rect 44637 32895 44695 32901
rect 44637 32861 44649 32895
rect 44683 32861 44695 32895
rect 44637 32855 44695 32861
rect 44726 32852 44732 32904
rect 44784 32892 44790 32904
rect 45281 32895 45339 32901
rect 45281 32892 45293 32895
rect 44784 32864 45293 32892
rect 44784 32852 44790 32864
rect 45281 32861 45293 32864
rect 45327 32861 45339 32895
rect 45281 32855 45339 32861
rect 45370 32852 45376 32904
rect 45428 32892 45434 32904
rect 45557 32895 45615 32901
rect 45557 32892 45569 32895
rect 45428 32864 45569 32892
rect 45428 32852 45434 32864
rect 45557 32861 45569 32864
rect 45603 32861 45615 32895
rect 45557 32855 45615 32861
rect 45808 32895 45866 32901
rect 45808 32861 45820 32895
rect 45854 32892 45866 32895
rect 46014 32892 46020 32904
rect 45854 32864 46020 32892
rect 45854 32861 45866 32864
rect 45808 32855 45866 32861
rect 46014 32852 46020 32864
rect 46072 32852 46078 32904
rect 42337 32827 42395 32833
rect 42337 32793 42349 32827
rect 42383 32793 42395 32827
rect 42337 32787 42395 32793
rect 43717 32827 43775 32833
rect 43717 32793 43729 32827
rect 43763 32824 43775 32827
rect 45925 32827 45983 32833
rect 43763 32796 45554 32824
rect 43763 32793 43775 32796
rect 43717 32787 43775 32793
rect 37016 32728 39068 32756
rect 35437 32719 35495 32725
rect 39666 32716 39672 32768
rect 39724 32716 39730 32768
rect 39942 32716 39948 32768
rect 40000 32716 40006 32768
rect 41598 32716 41604 32768
rect 41656 32756 41662 32768
rect 42352 32756 42380 32787
rect 41656 32728 42380 32756
rect 41656 32716 41662 32728
rect 44358 32716 44364 32768
rect 44416 32716 44422 32768
rect 44450 32716 44456 32768
rect 44508 32756 44514 32768
rect 44545 32759 44603 32765
rect 44545 32756 44557 32759
rect 44508 32728 44557 32756
rect 44508 32716 44514 32728
rect 44545 32725 44557 32728
rect 44591 32725 44603 32759
rect 45526 32756 45554 32796
rect 45925 32793 45937 32827
rect 45971 32824 45983 32827
rect 46198 32824 46204 32836
rect 45971 32796 46204 32824
rect 45971 32793 45983 32796
rect 45925 32787 45983 32793
rect 46198 32784 46204 32796
rect 46256 32784 46262 32836
rect 46308 32824 46336 32923
rect 47044 32901 47072 32932
rect 47596 32904 47624 32932
rect 47762 32920 47768 32972
rect 47820 32960 47826 32972
rect 48041 32963 48099 32969
rect 48041 32960 48053 32963
rect 47820 32932 48053 32960
rect 47820 32920 47826 32932
rect 48041 32929 48053 32932
rect 48087 32929 48099 32963
rect 48041 32923 48099 32929
rect 48774 32920 48780 32972
rect 48832 32960 48838 32972
rect 49602 32960 49608 32972
rect 48832 32932 49608 32960
rect 48832 32920 48838 32932
rect 49602 32920 49608 32932
rect 49660 32960 49666 32972
rect 49881 32963 49939 32969
rect 49881 32960 49893 32963
rect 49660 32932 49893 32960
rect 49660 32920 49666 32932
rect 49881 32929 49893 32932
rect 49927 32929 49939 32963
rect 49881 32923 49939 32929
rect 47029 32895 47087 32901
rect 47029 32861 47041 32895
rect 47075 32861 47087 32895
rect 47029 32855 47087 32861
rect 47210 32852 47216 32904
rect 47268 32852 47274 32904
rect 47302 32852 47308 32904
rect 47360 32852 47366 32904
rect 47486 32852 47492 32904
rect 47544 32852 47550 32904
rect 47578 32852 47584 32904
rect 47636 32852 47642 32904
rect 47670 32852 47676 32904
rect 47728 32852 47734 32904
rect 46753 32827 46811 32833
rect 46753 32824 46765 32827
rect 46308 32796 46765 32824
rect 46753 32793 46765 32796
rect 46799 32793 46811 32827
rect 46753 32787 46811 32793
rect 47121 32827 47179 32833
rect 47121 32793 47133 32827
rect 47167 32824 47179 32827
rect 48317 32827 48375 32833
rect 48317 32824 48329 32827
rect 47167 32796 48329 32824
rect 47167 32793 47179 32796
rect 47121 32787 47179 32793
rect 48317 32793 48329 32796
rect 48363 32793 48375 32827
rect 48317 32787 48375 32793
rect 48774 32784 48780 32836
rect 48832 32784 48838 32836
rect 45649 32759 45707 32765
rect 45649 32756 45661 32759
rect 45526 32728 45661 32756
rect 44545 32719 44603 32725
rect 45649 32725 45661 32728
rect 45695 32725 45707 32759
rect 45649 32719 45707 32725
rect 46017 32759 46075 32765
rect 46017 32725 46029 32759
rect 46063 32756 46075 32759
rect 46106 32756 46112 32768
rect 46063 32728 46112 32756
rect 46063 32725 46075 32728
rect 46017 32719 46075 32725
rect 46106 32716 46112 32728
rect 46164 32716 46170 32768
rect 46566 32765 46572 32768
rect 46553 32759 46572 32765
rect 46553 32725 46565 32759
rect 46553 32719 46572 32725
rect 46566 32716 46572 32719
rect 46624 32716 46630 32768
rect 49786 32716 49792 32768
rect 49844 32716 49850 32768
rect 1104 32666 78844 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 66314 32666
rect 66366 32614 66378 32666
rect 66430 32614 66442 32666
rect 66494 32614 66506 32666
rect 66558 32614 66570 32666
rect 66622 32614 78844 32666
rect 1104 32592 78844 32614
rect 27338 32552 27344 32564
rect 26988 32524 27344 32552
rect 17678 32484 17684 32496
rect 17144 32456 17684 32484
rect 17144 32425 17172 32456
rect 17678 32444 17684 32456
rect 17736 32444 17742 32496
rect 18690 32484 18696 32496
rect 18630 32456 18696 32484
rect 18690 32444 18696 32456
rect 18748 32484 18754 32496
rect 18969 32487 19027 32493
rect 18969 32484 18981 32487
rect 18748 32456 18981 32484
rect 18748 32444 18754 32456
rect 18969 32453 18981 32456
rect 19015 32453 19027 32487
rect 18969 32447 19027 32453
rect 26988 32425 27016 32524
rect 27338 32512 27344 32524
rect 27396 32552 27402 32564
rect 30190 32552 30196 32564
rect 27396 32524 30196 32552
rect 27396 32512 27402 32524
rect 30190 32512 30196 32524
rect 30248 32512 30254 32564
rect 30282 32512 30288 32564
rect 30340 32512 30346 32564
rect 32493 32555 32551 32561
rect 32493 32521 32505 32555
rect 32539 32552 32551 32555
rect 33042 32552 33048 32564
rect 32539 32524 33048 32552
rect 32539 32521 32551 32524
rect 32493 32515 32551 32521
rect 33042 32512 33048 32524
rect 33100 32512 33106 32564
rect 36170 32552 36176 32564
rect 34348 32524 36176 32552
rect 33962 32444 33968 32496
rect 34020 32444 34026 32496
rect 17129 32419 17187 32425
rect 17129 32385 17141 32419
rect 17175 32385 17187 32419
rect 17129 32379 17187 32385
rect 26973 32419 27031 32425
rect 26973 32385 26985 32419
rect 27019 32385 27031 32419
rect 26973 32379 27031 32385
rect 28350 32376 28356 32428
rect 28408 32376 28414 32428
rect 28994 32376 29000 32428
rect 29052 32376 29058 32428
rect 29730 32376 29736 32428
rect 29788 32376 29794 32428
rect 30006 32376 30012 32428
rect 30064 32416 30070 32428
rect 30101 32419 30159 32425
rect 30101 32416 30113 32419
rect 30064 32388 30113 32416
rect 30064 32376 30070 32388
rect 30101 32385 30113 32388
rect 30147 32385 30159 32419
rect 30101 32379 30159 32385
rect 31021 32419 31079 32425
rect 31021 32385 31033 32419
rect 31067 32416 31079 32419
rect 31113 32419 31171 32425
rect 31113 32416 31125 32419
rect 31067 32388 31125 32416
rect 31067 32385 31079 32388
rect 31021 32379 31079 32385
rect 31113 32385 31125 32388
rect 31159 32385 31171 32419
rect 31113 32379 31171 32385
rect 31294 32376 31300 32428
rect 31352 32376 31358 32428
rect 32858 32376 32864 32428
rect 32916 32376 32922 32428
rect 34348 32425 34376 32524
rect 36170 32512 36176 32524
rect 36228 32512 36234 32564
rect 45186 32512 45192 32564
rect 45244 32512 45250 32564
rect 46201 32555 46259 32561
rect 46201 32521 46213 32555
rect 46247 32552 46259 32555
rect 46382 32552 46388 32564
rect 46247 32524 46388 32552
rect 46247 32521 46259 32524
rect 46201 32515 46259 32521
rect 46382 32512 46388 32524
rect 46440 32512 46446 32564
rect 47578 32512 47584 32564
rect 47636 32512 47642 32564
rect 37366 32484 37372 32496
rect 35834 32456 37372 32484
rect 37366 32444 37372 32456
rect 37424 32444 37430 32496
rect 45357 32487 45415 32493
rect 45357 32453 45369 32487
rect 45403 32484 45415 32487
rect 45403 32456 45508 32484
rect 45403 32453 45415 32456
rect 45357 32447 45415 32453
rect 34241 32419 34299 32425
rect 34241 32385 34253 32419
rect 34287 32416 34299 32419
rect 34333 32419 34391 32425
rect 34333 32416 34345 32419
rect 34287 32388 34345 32416
rect 34287 32385 34299 32388
rect 34241 32379 34299 32385
rect 34333 32385 34345 32388
rect 34379 32385 34391 32419
rect 34333 32379 34391 32385
rect 43717 32419 43775 32425
rect 43717 32385 43729 32419
rect 43763 32416 43775 32419
rect 43806 32416 43812 32428
rect 43763 32388 43812 32416
rect 43763 32385 43775 32388
rect 43717 32379 43775 32385
rect 43806 32376 43812 32388
rect 43864 32376 43870 32428
rect 44085 32419 44143 32425
rect 44085 32385 44097 32419
rect 44131 32416 44143 32419
rect 44174 32416 44180 32428
rect 44131 32388 44180 32416
rect 44131 32385 44143 32388
rect 44085 32379 44143 32385
rect 44174 32376 44180 32388
rect 44232 32376 44238 32428
rect 44450 32376 44456 32428
rect 44508 32376 44514 32428
rect 44634 32376 44640 32428
rect 44692 32376 44698 32428
rect 45480 32416 45508 32456
rect 45554 32444 45560 32496
rect 45612 32444 45618 32496
rect 45833 32487 45891 32493
rect 45833 32453 45845 32487
rect 45879 32484 45891 32487
rect 45922 32484 45928 32496
rect 45879 32456 45928 32484
rect 45879 32453 45891 32456
rect 45833 32447 45891 32453
rect 45922 32444 45928 32456
rect 45980 32444 45986 32496
rect 46014 32444 46020 32496
rect 46072 32493 46078 32496
rect 46072 32487 46107 32493
rect 46095 32484 46107 32487
rect 46095 32456 47164 32484
rect 46095 32453 46107 32456
rect 46072 32447 46107 32453
rect 46072 32444 46078 32447
rect 46032 32416 46060 32444
rect 45480 32388 46060 32416
rect 2038 32308 2044 32360
rect 2096 32308 2102 32360
rect 17402 32308 17408 32360
rect 17460 32308 17466 32360
rect 27246 32308 27252 32360
rect 27304 32308 27310 32360
rect 28721 32351 28779 32357
rect 28721 32317 28733 32351
rect 28767 32348 28779 32351
rect 29178 32348 29184 32360
rect 28767 32320 29184 32348
rect 28767 32317 28779 32320
rect 28721 32311 28779 32317
rect 29178 32308 29184 32320
rect 29236 32308 29242 32360
rect 29641 32351 29699 32357
rect 29641 32317 29653 32351
rect 29687 32348 29699 32351
rect 29914 32348 29920 32360
rect 29687 32320 29920 32348
rect 29687 32317 29699 32320
rect 29641 32311 29699 32317
rect 29914 32308 29920 32320
rect 29972 32308 29978 32360
rect 30374 32308 30380 32360
rect 30432 32308 30438 32360
rect 34609 32351 34667 32357
rect 34609 32317 34621 32351
rect 34655 32348 34667 32351
rect 34698 32348 34704 32360
rect 34655 32320 34704 32348
rect 34655 32317 34667 32320
rect 34609 32311 34667 32317
rect 34698 32308 34704 32320
rect 34756 32308 34762 32360
rect 35986 32308 35992 32360
rect 36044 32348 36050 32360
rect 36081 32351 36139 32357
rect 36081 32348 36093 32351
rect 36044 32320 36093 32348
rect 36044 32308 36050 32320
rect 36081 32317 36093 32320
rect 36127 32348 36139 32351
rect 36725 32351 36783 32357
rect 36725 32348 36737 32351
rect 36127 32320 36737 32348
rect 36127 32317 36139 32320
rect 36081 32311 36139 32317
rect 36725 32317 36737 32320
rect 36771 32317 36783 32351
rect 36725 32311 36783 32317
rect 39666 32308 39672 32360
rect 39724 32348 39730 32360
rect 46566 32348 46572 32360
rect 39724 32320 46572 32348
rect 39724 32308 39730 32320
rect 46566 32308 46572 32320
rect 46624 32308 46630 32360
rect 47136 32348 47164 32456
rect 47210 32444 47216 32496
rect 47268 32484 47274 32496
rect 48041 32487 48099 32493
rect 48041 32484 48053 32487
rect 47268 32456 48053 32484
rect 47268 32444 47274 32456
rect 48041 32453 48053 32456
rect 48087 32453 48099 32487
rect 48041 32447 48099 32453
rect 47762 32376 47768 32428
rect 47820 32416 47826 32428
rect 48225 32419 48283 32425
rect 48225 32416 48237 32419
rect 47820 32388 48237 32416
rect 47820 32376 47826 32388
rect 48225 32385 48237 32388
rect 48271 32385 48283 32419
rect 48225 32379 48283 32385
rect 48317 32419 48375 32425
rect 48317 32385 48329 32419
rect 48363 32416 48375 32419
rect 49786 32416 49792 32428
rect 48363 32388 49792 32416
rect 48363 32385 48375 32388
rect 48317 32379 48375 32385
rect 47949 32351 48007 32357
rect 47949 32348 47961 32351
rect 47136 32320 47961 32348
rect 47949 32317 47961 32320
rect 47995 32317 48007 32351
rect 47949 32311 48007 32317
rect 29196 32280 29224 32308
rect 29196 32252 30052 32280
rect 18506 32172 18512 32224
rect 18564 32212 18570 32224
rect 18877 32215 18935 32221
rect 18877 32212 18889 32215
rect 18564 32184 18889 32212
rect 18564 32172 18570 32184
rect 18877 32181 18889 32184
rect 18923 32181 18935 32215
rect 18877 32175 18935 32181
rect 27706 32172 27712 32224
rect 27764 32212 27770 32224
rect 28810 32212 28816 32224
rect 27764 32184 28816 32212
rect 27764 32172 27770 32184
rect 28810 32172 28816 32184
rect 28868 32172 28874 32224
rect 29362 32172 29368 32224
rect 29420 32172 29426 32224
rect 30024 32221 30052 32252
rect 43530 32240 43536 32292
rect 43588 32240 43594 32292
rect 46198 32280 46204 32292
rect 45388 32252 46204 32280
rect 30009 32215 30067 32221
rect 30009 32181 30021 32215
rect 30055 32181 30067 32215
rect 30009 32175 30067 32181
rect 31113 32215 31171 32221
rect 31113 32181 31125 32215
rect 31159 32212 31171 32215
rect 31386 32212 31392 32224
rect 31159 32184 31392 32212
rect 31159 32181 31171 32184
rect 31113 32175 31171 32181
rect 31386 32172 31392 32184
rect 31444 32172 31450 32224
rect 36170 32172 36176 32224
rect 36228 32172 36234 32224
rect 45388 32221 45416 32252
rect 46198 32240 46204 32252
rect 46256 32240 46262 32292
rect 47964 32280 47992 32311
rect 48038 32308 48044 32360
rect 48096 32308 48102 32360
rect 48332 32280 48360 32379
rect 49786 32376 49792 32388
rect 49844 32376 49850 32428
rect 47964 32252 48360 32280
rect 45373 32215 45431 32221
rect 45373 32181 45385 32215
rect 45419 32181 45431 32215
rect 45373 32175 45431 32181
rect 45554 32172 45560 32224
rect 45612 32212 45618 32224
rect 46017 32215 46075 32221
rect 46017 32212 46029 32215
rect 45612 32184 46029 32212
rect 45612 32172 45618 32184
rect 46017 32181 46029 32184
rect 46063 32212 46075 32215
rect 46106 32212 46112 32224
rect 46063 32184 46112 32212
rect 46063 32181 46075 32184
rect 46017 32175 46075 32181
rect 46106 32172 46112 32184
rect 46164 32212 46170 32224
rect 46382 32212 46388 32224
rect 46164 32184 46388 32212
rect 46164 32172 46170 32184
rect 46382 32172 46388 32184
rect 46440 32172 46446 32224
rect 47302 32172 47308 32224
rect 47360 32212 47366 32224
rect 48038 32212 48044 32224
rect 47360 32184 48044 32212
rect 47360 32172 47366 32184
rect 48038 32172 48044 32184
rect 48096 32172 48102 32224
rect 1104 32122 78844 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 78844 32122
rect 1104 32048 78844 32070
rect 1302 31968 1308 32020
rect 1360 32008 1366 32020
rect 1857 32011 1915 32017
rect 1857 32008 1869 32011
rect 1360 31980 1869 32008
rect 1360 31968 1366 31980
rect 1857 31977 1869 31980
rect 1903 31977 1915 32011
rect 1857 31971 1915 31977
rect 17129 32011 17187 32017
rect 17129 31977 17141 32011
rect 17175 32008 17187 32011
rect 17402 32008 17408 32020
rect 17175 31980 17408 32008
rect 17175 31977 17187 31980
rect 17129 31971 17187 31977
rect 17402 31968 17408 31980
rect 17460 31968 17466 32020
rect 27246 31968 27252 32020
rect 27304 32008 27310 32020
rect 27985 32011 28043 32017
rect 27985 32008 27997 32011
rect 27304 31980 27997 32008
rect 27304 31968 27310 31980
rect 27985 31977 27997 31980
rect 28031 31977 28043 32011
rect 27985 31971 28043 31977
rect 29825 32011 29883 32017
rect 29825 31977 29837 32011
rect 29871 32008 29883 32011
rect 30374 32008 30380 32020
rect 29871 31980 30380 32008
rect 29871 31977 29883 31980
rect 29825 31971 29883 31977
rect 30374 31968 30380 31980
rect 30432 31968 30438 32020
rect 31386 31968 31392 32020
rect 31444 32017 31450 32020
rect 31444 32011 31459 32017
rect 31447 31977 31459 32011
rect 31444 31971 31459 31977
rect 31444 31968 31450 31971
rect 34698 31968 34704 32020
rect 34756 31968 34762 32020
rect 35069 32011 35127 32017
rect 35069 31977 35081 32011
rect 35115 32008 35127 32011
rect 35434 32008 35440 32020
rect 35115 31980 35440 32008
rect 35115 31977 35127 31980
rect 35069 31971 35127 31977
rect 35434 31968 35440 31980
rect 35492 31968 35498 32020
rect 43993 32011 44051 32017
rect 43993 31977 44005 32011
rect 44039 32008 44051 32011
rect 44450 32008 44456 32020
rect 44039 31980 44456 32008
rect 44039 31977 44051 31980
rect 43993 31971 44051 31977
rect 44450 31968 44456 31980
rect 44508 31968 44514 32020
rect 46293 32011 46351 32017
rect 46293 31977 46305 32011
rect 46339 32008 46351 32011
rect 46382 32008 46388 32020
rect 46339 31980 46388 32008
rect 46339 31977 46351 31980
rect 46293 31971 46351 31977
rect 46382 31968 46388 31980
rect 46440 31968 46446 32020
rect 46477 32011 46535 32017
rect 46477 31977 46489 32011
rect 46523 32008 46535 32011
rect 47118 32008 47124 32020
rect 46523 31980 47124 32008
rect 46523 31977 46535 31980
rect 46477 31971 46535 31977
rect 47118 31968 47124 31980
rect 47176 32008 47182 32020
rect 47762 32008 47768 32020
rect 47176 31980 47768 32008
rect 47176 31968 47182 31980
rect 47762 31968 47768 31980
rect 47820 31968 47826 32020
rect 28350 31900 28356 31952
rect 28408 31940 28414 31952
rect 43882 31943 43940 31949
rect 28408 31912 30328 31940
rect 28408 31900 28414 31912
rect 16669 31875 16727 31881
rect 16669 31841 16681 31875
rect 16715 31841 16727 31875
rect 16669 31835 16727 31841
rect 2038 31764 2044 31816
rect 2096 31764 2102 31816
rect 11330 31764 11336 31816
rect 11388 31804 11394 31816
rect 12069 31807 12127 31813
rect 12069 31804 12081 31807
rect 11388 31776 12081 31804
rect 11388 31764 11394 31776
rect 12069 31773 12081 31776
rect 12115 31773 12127 31807
rect 12069 31767 12127 31773
rect 15378 31764 15384 31816
rect 15436 31764 15442 31816
rect 15565 31807 15623 31813
rect 15565 31773 15577 31807
rect 15611 31804 15623 31807
rect 16684 31804 16712 31835
rect 17678 31832 17684 31884
rect 17736 31872 17742 31884
rect 21450 31872 21456 31884
rect 17736 31844 21456 31872
rect 17736 31832 17742 31844
rect 21450 31832 21456 31844
rect 21508 31872 21514 31884
rect 26970 31872 26976 31884
rect 21508 31844 26976 31872
rect 21508 31832 21514 31844
rect 26970 31832 26976 31844
rect 27028 31832 27034 31884
rect 15611 31776 16712 31804
rect 16761 31807 16819 31813
rect 15611 31773 15623 31776
rect 15565 31767 15623 31773
rect 12342 31696 12348 31748
rect 12400 31696 12406 31748
rect 13630 31736 13636 31748
rect 13570 31708 13636 31736
rect 13630 31696 13636 31708
rect 13688 31736 13694 31748
rect 14185 31739 14243 31745
rect 14185 31736 14197 31739
rect 13688 31708 14197 31736
rect 13688 31696 13694 31708
rect 14185 31705 14197 31708
rect 14231 31736 14243 31739
rect 14734 31736 14740 31748
rect 14231 31708 14740 31736
rect 14231 31705 14243 31708
rect 14185 31699 14243 31705
rect 14734 31696 14740 31708
rect 14792 31736 14798 31748
rect 16298 31736 16304 31748
rect 14792 31708 16304 31736
rect 14792 31696 14798 31708
rect 16298 31696 16304 31708
rect 16356 31696 16362 31748
rect 16546 31736 16574 31776
rect 16761 31773 16773 31807
rect 16807 31804 16819 31807
rect 17865 31807 17923 31813
rect 17865 31804 17877 31807
rect 16807 31776 17877 31804
rect 16807 31773 16819 31776
rect 16761 31767 16819 31773
rect 17865 31773 17877 31776
rect 17911 31773 17923 31807
rect 17865 31767 17923 31773
rect 18506 31764 18512 31816
rect 18564 31804 18570 31816
rect 18782 31804 18788 31816
rect 18564 31776 18788 31804
rect 18564 31764 18570 31776
rect 18782 31764 18788 31776
rect 18840 31764 18846 31816
rect 27706 31764 27712 31816
rect 27764 31804 27770 31816
rect 27801 31807 27859 31813
rect 27801 31804 27813 31807
rect 27764 31776 27813 31804
rect 27764 31764 27770 31776
rect 27801 31773 27813 31776
rect 27847 31773 27859 31807
rect 27801 31767 27859 31773
rect 27982 31764 27988 31816
rect 28040 31764 28046 31816
rect 28810 31764 28816 31816
rect 28868 31804 28874 31816
rect 29549 31807 29607 31813
rect 29549 31804 29561 31807
rect 28868 31776 29561 31804
rect 28868 31764 28874 31776
rect 29549 31773 29561 31776
rect 29595 31773 29607 31807
rect 29549 31767 29607 31773
rect 29825 31807 29883 31813
rect 29825 31773 29837 31807
rect 29871 31804 29883 31807
rect 29871 31776 30144 31804
rect 30300 31790 30328 31912
rect 43882 31909 43894 31943
rect 43928 31940 43940 31943
rect 44174 31940 44180 31952
rect 43928 31912 44180 31940
rect 43928 31909 43940 31912
rect 43882 31903 43940 31909
rect 44174 31900 44180 31912
rect 44232 31900 44238 31952
rect 44361 31943 44419 31949
rect 44361 31909 44373 31943
rect 44407 31940 44419 31943
rect 44542 31940 44548 31952
rect 44407 31912 44548 31940
rect 44407 31909 44419 31912
rect 44361 31903 44419 31909
rect 44542 31900 44548 31912
rect 44600 31900 44606 31952
rect 30374 31832 30380 31884
rect 30432 31872 30438 31884
rect 31665 31875 31723 31881
rect 31665 31872 31677 31875
rect 30432 31844 31677 31872
rect 30432 31832 30438 31844
rect 31665 31841 31677 31844
rect 31711 31841 31723 31875
rect 31665 31835 31723 31841
rect 35161 31875 35219 31881
rect 35161 31841 35173 31875
rect 35207 31872 35219 31875
rect 36170 31872 36176 31884
rect 35207 31844 36176 31872
rect 35207 31841 35219 31844
rect 35161 31835 35219 31841
rect 36170 31832 36176 31844
rect 36228 31832 36234 31884
rect 40678 31832 40684 31884
rect 40736 31872 40742 31884
rect 44085 31875 44143 31881
rect 44085 31872 44097 31875
rect 40736 31844 44097 31872
rect 40736 31832 40742 31844
rect 44085 31841 44097 31844
rect 44131 31872 44143 31875
rect 44634 31872 44640 31884
rect 44131 31844 44640 31872
rect 44131 31841 44143 31844
rect 44085 31835 44143 31841
rect 44634 31832 44640 31844
rect 44692 31832 44698 31884
rect 34885 31807 34943 31813
rect 29871 31773 29883 31776
rect 29825 31767 29883 31773
rect 17126 31736 17132 31748
rect 16546 31708 17132 31736
rect 17126 31696 17132 31708
rect 17184 31696 17190 31748
rect 20162 31696 20168 31748
rect 20220 31736 20226 31748
rect 20625 31739 20683 31745
rect 20625 31736 20637 31739
rect 20220 31708 20637 31736
rect 20220 31696 20226 31708
rect 20625 31705 20637 31708
rect 20671 31736 20683 31739
rect 21637 31739 21695 31745
rect 21637 31736 21649 31739
rect 20671 31708 21649 31736
rect 20671 31705 20683 31708
rect 20625 31699 20683 31705
rect 21637 31705 21649 31708
rect 21683 31705 21695 31739
rect 21637 31699 21695 31705
rect 29641 31739 29699 31745
rect 29641 31705 29653 31739
rect 29687 31736 29699 31739
rect 30006 31736 30012 31748
rect 29687 31708 30012 31736
rect 29687 31705 29699 31708
rect 29641 31699 29699 31705
rect 30006 31696 30012 31708
rect 30064 31696 30070 31748
rect 2038 31628 2044 31680
rect 2096 31668 2102 31680
rect 2133 31671 2191 31677
rect 2133 31668 2145 31671
rect 2096 31640 2145 31668
rect 2096 31628 2102 31640
rect 2133 31637 2145 31640
rect 2179 31637 2191 31671
rect 2133 31631 2191 31637
rect 13814 31628 13820 31680
rect 13872 31628 13878 31680
rect 15286 31628 15292 31680
rect 15344 31668 15350 31680
rect 15473 31671 15531 31677
rect 15473 31668 15485 31671
rect 15344 31640 15485 31668
rect 15344 31628 15350 31640
rect 15473 31637 15485 31640
rect 15519 31637 15531 31671
rect 15473 31631 15531 31637
rect 29914 31628 29920 31680
rect 29972 31628 29978 31680
rect 30116 31668 30144 31776
rect 34885 31773 34897 31807
rect 34931 31804 34943 31807
rect 35342 31804 35348 31816
rect 34931 31776 35348 31804
rect 34931 31773 34943 31776
rect 34885 31767 34943 31773
rect 35342 31764 35348 31776
rect 35400 31764 35406 31816
rect 37274 31764 37280 31816
rect 37332 31804 37338 31816
rect 41414 31804 41420 31816
rect 37332 31776 41420 31804
rect 37332 31764 37338 31776
rect 41414 31764 41420 31776
rect 41472 31804 41478 31816
rect 41690 31804 41696 31816
rect 41472 31776 41696 31804
rect 41472 31764 41478 31776
rect 41690 31764 41696 31776
rect 41748 31764 41754 31816
rect 43717 31807 43775 31813
rect 43717 31773 43729 31807
rect 43763 31804 43775 31807
rect 43806 31804 43812 31816
rect 43763 31776 43812 31804
rect 43763 31773 43775 31776
rect 43717 31767 43775 31773
rect 43806 31764 43812 31776
rect 43864 31764 43870 31816
rect 44358 31764 44364 31816
rect 44416 31804 44422 31816
rect 45370 31804 45376 31816
rect 44416 31776 45376 31804
rect 44416 31764 44422 31776
rect 45370 31764 45376 31776
rect 45428 31764 45434 31816
rect 46106 31696 46112 31748
rect 46164 31696 46170 31748
rect 46290 31696 46296 31748
rect 46348 31745 46354 31748
rect 46348 31739 46383 31745
rect 46371 31736 46383 31739
rect 46566 31736 46572 31748
rect 46371 31708 46572 31736
rect 46371 31705 46383 31708
rect 46348 31699 46383 31705
rect 46348 31696 46354 31699
rect 46566 31696 46572 31708
rect 46624 31696 46630 31748
rect 30742 31668 30748 31680
rect 30116 31640 30748 31668
rect 30742 31628 30748 31640
rect 30800 31628 30806 31680
rect 36722 31628 36728 31680
rect 36780 31668 36786 31680
rect 37461 31671 37519 31677
rect 37461 31668 37473 31671
rect 36780 31640 37473 31668
rect 36780 31628 36786 31640
rect 37461 31637 37473 31640
rect 37507 31668 37519 31671
rect 39114 31668 39120 31680
rect 37507 31640 39120 31668
rect 37507 31637 37519 31640
rect 37461 31631 37519 31637
rect 39114 31628 39120 31640
rect 39172 31668 39178 31680
rect 40494 31668 40500 31680
rect 39172 31640 40500 31668
rect 39172 31628 39178 31640
rect 40494 31628 40500 31640
rect 40552 31668 40558 31680
rect 45094 31668 45100 31680
rect 40552 31640 45100 31668
rect 40552 31628 40558 31640
rect 45094 31628 45100 31640
rect 45152 31628 45158 31680
rect 1104 31578 78844 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 66314 31578
rect 66366 31526 66378 31578
rect 66430 31526 66442 31578
rect 66494 31526 66506 31578
rect 66558 31526 66570 31578
rect 66622 31526 78844 31578
rect 1104 31504 78844 31526
rect 934 31424 940 31476
rect 992 31464 998 31476
rect 1857 31467 1915 31473
rect 1857 31464 1869 31467
rect 992 31436 1869 31464
rect 992 31424 998 31436
rect 1857 31433 1869 31436
rect 1903 31433 1915 31467
rect 1857 31427 1915 31433
rect 12345 31467 12403 31473
rect 12345 31433 12357 31467
rect 12391 31464 12403 31467
rect 13630 31464 13636 31476
rect 12391 31436 13636 31464
rect 12391 31433 12403 31436
rect 12345 31427 12403 31433
rect 11606 31396 11612 31408
rect 11086 31368 11612 31396
rect 11606 31356 11612 31368
rect 11664 31396 11670 31408
rect 12360 31396 12388 31427
rect 13630 31424 13636 31436
rect 13688 31424 13694 31476
rect 17497 31467 17555 31473
rect 17497 31433 17509 31467
rect 17543 31464 17555 31467
rect 18690 31464 18696 31476
rect 17543 31436 18696 31464
rect 17543 31433 17555 31436
rect 17497 31427 17555 31433
rect 11664 31368 12388 31396
rect 15013 31399 15071 31405
rect 11664 31356 11670 31368
rect 15013 31365 15025 31399
rect 15059 31396 15071 31399
rect 15286 31396 15292 31408
rect 15059 31368 15292 31396
rect 15059 31365 15071 31368
rect 15013 31359 15071 31365
rect 15286 31356 15292 31368
rect 15344 31356 15350 31408
rect 16298 31396 16304 31408
rect 16238 31368 16304 31396
rect 16298 31356 16304 31368
rect 16356 31396 16362 31408
rect 17512 31396 17540 31427
rect 18690 31424 18696 31436
rect 18748 31424 18754 31476
rect 28810 31424 28816 31476
rect 28868 31464 28874 31476
rect 29799 31467 29857 31473
rect 29799 31464 29811 31467
rect 28868 31436 29811 31464
rect 28868 31424 28874 31436
rect 29799 31433 29811 31436
rect 29845 31433 29857 31467
rect 29799 31427 29857 31433
rect 30742 31424 30748 31476
rect 30800 31464 30806 31476
rect 30837 31467 30895 31473
rect 30837 31464 30849 31467
rect 30800 31436 30849 31464
rect 30800 31424 30806 31436
rect 30837 31433 30849 31436
rect 30883 31433 30895 31467
rect 30837 31427 30895 31433
rect 37384 31436 38654 31464
rect 37384 31408 37412 31436
rect 20346 31396 20352 31408
rect 16356 31368 17540 31396
rect 19182 31368 20352 31396
rect 16356 31356 16362 31368
rect 20346 31356 20352 31368
rect 20404 31356 20410 31408
rect 30006 31396 30012 31408
rect 29196 31368 30012 31396
rect 2038 31288 2044 31340
rect 2096 31288 2102 31340
rect 11422 31288 11428 31340
rect 11480 31328 11486 31340
rect 14737 31331 14795 31337
rect 14737 31328 14749 31331
rect 11480 31300 14749 31328
rect 11480 31288 11486 31300
rect 14737 31297 14749 31300
rect 14783 31297 14795 31331
rect 14737 31291 14795 31297
rect 17678 31288 17684 31340
rect 17736 31288 17742 31340
rect 27801 31331 27859 31337
rect 27801 31297 27813 31331
rect 27847 31328 27859 31331
rect 28537 31331 28595 31337
rect 28537 31328 28549 31331
rect 27847 31300 28549 31328
rect 27847 31297 27859 31300
rect 27801 31291 27859 31297
rect 28537 31297 28549 31300
rect 28583 31297 28595 31331
rect 28537 31291 28595 31297
rect 29086 31288 29092 31340
rect 29144 31328 29150 31340
rect 29196 31337 29224 31368
rect 30006 31356 30012 31368
rect 30064 31356 30070 31408
rect 35986 31356 35992 31408
rect 36044 31396 36050 31408
rect 36722 31396 36728 31408
rect 36044 31368 36728 31396
rect 36044 31356 36050 31368
rect 36722 31356 36728 31368
rect 36780 31356 36786 31408
rect 36941 31399 36999 31405
rect 36941 31365 36953 31399
rect 36987 31396 36999 31399
rect 37366 31396 37372 31408
rect 36987 31368 37372 31396
rect 36987 31365 36999 31368
rect 36941 31359 36999 31365
rect 37366 31356 37372 31368
rect 37424 31356 37430 31408
rect 38626 31396 38654 31436
rect 40052 31436 40632 31464
rect 40052 31405 40080 31436
rect 40037 31399 40095 31405
rect 40037 31396 40049 31399
rect 38626 31368 40049 31396
rect 29181 31331 29239 31337
rect 29181 31328 29193 31331
rect 29144 31300 29193 31328
rect 29144 31288 29150 31300
rect 29181 31297 29193 31300
rect 29227 31297 29239 31331
rect 29181 31291 29239 31297
rect 37274 31288 37280 31340
rect 37332 31328 37338 31340
rect 39776 31337 39804 31368
rect 40037 31365 40049 31368
rect 40083 31365 40095 31399
rect 40037 31359 40095 31365
rect 40494 31356 40500 31408
rect 40552 31356 40558 31408
rect 40604 31396 40632 31436
rect 40678 31424 40684 31476
rect 40736 31473 40742 31476
rect 40736 31467 40755 31473
rect 40743 31433 40755 31467
rect 40736 31427 40755 31433
rect 40736 31424 40742 31427
rect 40862 31424 40868 31476
rect 40920 31464 40926 31476
rect 41049 31467 41107 31473
rect 41049 31464 41061 31467
rect 40920 31436 41061 31464
rect 40920 31424 40926 31436
rect 41049 31433 41061 31436
rect 41095 31433 41107 31467
rect 41049 31427 41107 31433
rect 42886 31396 42892 31408
rect 40604 31368 40724 31396
rect 39761 31331 39819 31337
rect 37332 31300 37674 31328
rect 37332 31288 37338 31300
rect 39761 31297 39773 31331
rect 39807 31297 39819 31331
rect 39761 31291 39819 31297
rect 39945 31331 40003 31337
rect 39945 31297 39957 31331
rect 39991 31297 40003 31331
rect 39945 31291 40003 31297
rect 40221 31331 40279 31337
rect 40221 31297 40233 31331
rect 40267 31297 40279 31331
rect 40696 31328 40724 31368
rect 41524 31368 42892 31396
rect 41524 31337 41552 31368
rect 42886 31356 42892 31368
rect 42944 31396 42950 31408
rect 44542 31396 44548 31408
rect 42944 31368 44548 31396
rect 42944 31356 42950 31368
rect 44542 31356 44548 31368
rect 44600 31356 44606 31408
rect 45097 31399 45155 31405
rect 45097 31365 45109 31399
rect 45143 31396 45155 31399
rect 45373 31399 45431 31405
rect 45373 31396 45385 31399
rect 45143 31368 45385 31396
rect 45143 31365 45155 31368
rect 45097 31359 45155 31365
rect 45373 31365 45385 31368
rect 45419 31365 45431 31399
rect 45833 31399 45891 31405
rect 45833 31396 45845 31399
rect 45373 31359 45431 31365
rect 45480 31368 45845 31396
rect 40957 31331 41015 31337
rect 40957 31328 40969 31331
rect 40696 31300 40969 31328
rect 40221 31291 40279 31297
rect 40957 31297 40969 31300
rect 41003 31297 41015 31331
rect 40957 31291 41015 31297
rect 41141 31331 41199 31337
rect 41141 31297 41153 31331
rect 41187 31297 41199 31331
rect 41141 31291 41199 31297
rect 41509 31331 41567 31337
rect 41509 31297 41521 31331
rect 41555 31297 41567 31331
rect 41509 31291 41567 31297
rect 9585 31263 9643 31269
rect 9585 31229 9597 31263
rect 9631 31260 9643 31263
rect 9631 31232 9720 31260
rect 9631 31229 9643 31232
rect 9585 31223 9643 31229
rect 9692 31136 9720 31232
rect 9858 31220 9864 31272
rect 9916 31220 9922 31272
rect 11333 31263 11391 31269
rect 11333 31229 11345 31263
rect 11379 31260 11391 31263
rect 11882 31260 11888 31272
rect 11379 31232 11888 31260
rect 11379 31229 11391 31232
rect 11333 31223 11391 31229
rect 11882 31220 11888 31232
rect 11940 31260 11946 31272
rect 12069 31263 12127 31269
rect 12069 31260 12081 31263
rect 11940 31232 12081 31260
rect 11940 31220 11946 31232
rect 12069 31229 12081 31232
rect 12115 31229 12127 31263
rect 12069 31223 12127 31229
rect 12250 31220 12256 31272
rect 12308 31260 12314 31272
rect 13357 31263 13415 31269
rect 13357 31260 13369 31263
rect 12308 31232 13369 31260
rect 12308 31220 12314 31232
rect 13357 31229 13369 31232
rect 13403 31260 13415 31263
rect 13814 31260 13820 31272
rect 13403 31232 13820 31260
rect 13403 31229 13415 31232
rect 13357 31223 13415 31229
rect 13814 31220 13820 31232
rect 13872 31260 13878 31272
rect 14093 31263 14151 31269
rect 14093 31260 14105 31263
rect 13872 31232 14105 31260
rect 13872 31220 13878 31232
rect 14093 31229 14105 31232
rect 14139 31229 14151 31263
rect 17221 31263 17279 31269
rect 17221 31260 17233 31263
rect 14093 31223 14151 31229
rect 16500 31232 17233 31260
rect 16500 31136 16528 31232
rect 17221 31229 17233 31232
rect 17267 31229 17279 31263
rect 17221 31223 17279 31229
rect 17957 31263 18015 31269
rect 17957 31229 17969 31263
rect 18003 31260 18015 31263
rect 18506 31260 18512 31272
rect 18003 31232 18512 31260
rect 18003 31229 18015 31232
rect 17957 31223 18015 31229
rect 18506 31220 18512 31232
rect 18564 31220 18570 31272
rect 18690 31220 18696 31272
rect 18748 31260 18754 31272
rect 19429 31263 19487 31269
rect 19429 31260 19441 31263
rect 18748 31232 19441 31260
rect 18748 31220 18754 31232
rect 19429 31229 19441 31232
rect 19475 31260 19487 31263
rect 20073 31263 20131 31269
rect 20073 31260 20085 31263
rect 19475 31232 20085 31260
rect 19475 31229 19487 31232
rect 19429 31223 19487 31229
rect 20073 31229 20085 31232
rect 20119 31229 20131 31263
rect 20073 31223 20131 31229
rect 27706 31220 27712 31272
rect 27764 31220 27770 31272
rect 29914 31220 29920 31272
rect 29972 31260 29978 31272
rect 31389 31263 31447 31269
rect 31389 31260 31401 31263
rect 29972 31232 31401 31260
rect 29972 31220 29978 31232
rect 31389 31229 31401 31232
rect 31435 31260 31447 31263
rect 31570 31260 31576 31272
rect 31435 31232 31576 31260
rect 31435 31229 31447 31232
rect 31389 31223 31447 31229
rect 31570 31220 31576 31232
rect 31628 31220 31634 31272
rect 38749 31263 38807 31269
rect 38749 31260 38761 31263
rect 37108 31232 38761 31260
rect 29641 31195 29699 31201
rect 29641 31161 29653 31195
rect 29687 31192 29699 31195
rect 29730 31192 29736 31204
rect 29687 31164 29736 31192
rect 29687 31161 29699 31164
rect 29641 31155 29699 31161
rect 29730 31152 29736 31164
rect 29788 31192 29794 31204
rect 31294 31192 31300 31204
rect 29788 31164 31300 31192
rect 29788 31152 29794 31164
rect 31294 31152 31300 31164
rect 31352 31152 31358 31204
rect 37108 31201 37136 31232
rect 38749 31229 38761 31232
rect 38795 31229 38807 31263
rect 39025 31263 39083 31269
rect 39025 31260 39037 31263
rect 38749 31223 38807 31229
rect 38948 31232 39037 31260
rect 37093 31195 37151 31201
rect 37093 31161 37105 31195
rect 37139 31161 37151 31195
rect 37093 31155 37151 31161
rect 9674 31084 9680 31136
rect 9732 31124 9738 31136
rect 11330 31124 11336 31136
rect 9732 31096 11336 31124
rect 9732 31084 9738 31096
rect 11330 31084 11336 31096
rect 11388 31084 11394 31136
rect 11422 31084 11428 31136
rect 11480 31124 11486 31136
rect 11517 31127 11575 31133
rect 11517 31124 11529 31127
rect 11480 31096 11529 31124
rect 11480 31084 11486 31096
rect 11517 31093 11529 31096
rect 11563 31093 11575 31127
rect 11517 31087 11575 31093
rect 12802 31084 12808 31136
rect 12860 31084 12866 31136
rect 13538 31084 13544 31136
rect 13596 31084 13602 31136
rect 16482 31084 16488 31136
rect 16540 31084 16546 31136
rect 16666 31084 16672 31136
rect 16724 31084 16730 31136
rect 19518 31084 19524 31136
rect 19576 31084 19582 31136
rect 20346 31084 20352 31136
rect 20404 31084 20410 31136
rect 27433 31127 27491 31133
rect 27433 31093 27445 31127
rect 27479 31124 27491 31127
rect 27614 31124 27620 31136
rect 27479 31096 27620 31124
rect 27479 31093 27491 31096
rect 27433 31087 27491 31093
rect 27614 31084 27620 31096
rect 27672 31084 27678 31136
rect 29825 31127 29883 31133
rect 29825 31093 29837 31127
rect 29871 31124 29883 31127
rect 29914 31124 29920 31136
rect 29871 31096 29920 31124
rect 29871 31093 29883 31096
rect 29825 31087 29883 31093
rect 29914 31084 29920 31096
rect 29972 31084 29978 31136
rect 36906 31084 36912 31136
rect 36964 31084 36970 31136
rect 37277 31127 37335 31133
rect 37277 31093 37289 31127
rect 37323 31124 37335 31127
rect 37458 31124 37464 31136
rect 37323 31096 37464 31124
rect 37323 31093 37335 31096
rect 37277 31087 37335 31093
rect 37458 31084 37464 31096
rect 37516 31084 37522 31136
rect 38654 31084 38660 31136
rect 38712 31124 38718 31136
rect 38948 31124 38976 31232
rect 39025 31229 39037 31232
rect 39071 31229 39083 31263
rect 39960 31260 39988 31291
rect 40236 31260 40264 31291
rect 40678 31260 40684 31272
rect 39960 31232 40684 31260
rect 39025 31223 39083 31229
rect 40678 31220 40684 31232
rect 40736 31260 40742 31272
rect 41156 31260 41184 31291
rect 41690 31288 41696 31340
rect 41748 31288 41754 31340
rect 42518 31288 42524 31340
rect 42576 31328 42582 31340
rect 44266 31328 44272 31340
rect 42576 31300 44272 31328
rect 42576 31288 42582 31300
rect 44266 31288 44272 31300
rect 44324 31288 44330 31340
rect 44729 31331 44787 31337
rect 44729 31297 44741 31331
rect 44775 31328 44787 31331
rect 45480 31328 45508 31368
rect 45833 31365 45845 31368
rect 45879 31396 45891 31399
rect 46845 31399 46903 31405
rect 45879 31368 46704 31396
rect 45879 31365 45891 31368
rect 45833 31359 45891 31365
rect 44775 31300 45508 31328
rect 45557 31331 45615 31337
rect 44775 31297 44787 31300
rect 44729 31291 44787 31297
rect 45557 31297 45569 31331
rect 45603 31297 45615 31331
rect 45557 31291 45615 31297
rect 45741 31331 45799 31337
rect 45741 31297 45753 31331
rect 45787 31328 45799 31331
rect 46017 31331 46075 31337
rect 46017 31328 46029 31331
rect 45787 31300 46029 31328
rect 45787 31297 45799 31300
rect 45741 31291 45799 31297
rect 46017 31297 46029 31300
rect 46063 31328 46075 31331
rect 46290 31328 46296 31340
rect 46063 31300 46296 31328
rect 46063 31297 46075 31300
rect 46017 31291 46075 31297
rect 40736 31232 41184 31260
rect 45572 31260 45600 31291
rect 46290 31288 46296 31300
rect 46348 31288 46354 31340
rect 46382 31288 46388 31340
rect 46440 31328 46446 31340
rect 46566 31328 46572 31340
rect 46440 31300 46572 31328
rect 46440 31288 46446 31300
rect 46566 31288 46572 31300
rect 46624 31288 46630 31340
rect 46676 31337 46704 31368
rect 46845 31365 46857 31399
rect 46891 31365 46903 31399
rect 46845 31359 46903 31365
rect 46661 31331 46719 31337
rect 46661 31297 46673 31331
rect 46707 31297 46719 31331
rect 46860 31328 46888 31359
rect 46937 31331 46995 31337
rect 46937 31328 46949 31331
rect 46860 31300 46949 31328
rect 46661 31291 46719 31297
rect 46937 31297 46949 31300
rect 46983 31297 46995 31331
rect 46937 31291 46995 31297
rect 47118 31288 47124 31340
rect 47176 31288 47182 31340
rect 46106 31260 46112 31272
rect 45572 31232 46112 31260
rect 40736 31220 40742 31232
rect 46106 31220 46112 31232
rect 46164 31260 46170 31272
rect 46201 31263 46259 31269
rect 46201 31260 46213 31263
rect 46164 31232 46213 31260
rect 46164 31220 46170 31232
rect 46201 31229 46213 31232
rect 46247 31260 46259 31263
rect 46750 31260 46756 31272
rect 46247 31232 46756 31260
rect 46247 31229 46259 31232
rect 46201 31223 46259 31229
rect 46750 31220 46756 31232
rect 46808 31220 46814 31272
rect 46845 31263 46903 31269
rect 46845 31229 46857 31263
rect 46891 31260 46903 31263
rect 47302 31260 47308 31272
rect 46891 31232 47308 31260
rect 46891 31229 46903 31232
rect 46845 31223 46903 31229
rect 39853 31195 39911 31201
rect 39853 31161 39865 31195
rect 39899 31192 39911 31195
rect 39899 31164 40724 31192
rect 39899 31161 39911 31164
rect 39853 31155 39911 31161
rect 38712 31096 38976 31124
rect 40313 31127 40371 31133
rect 38712 31084 38718 31096
rect 40313 31093 40325 31127
rect 40359 31124 40371 31127
rect 40586 31124 40592 31136
rect 40359 31096 40592 31124
rect 40359 31093 40371 31096
rect 40313 31087 40371 31093
rect 40586 31084 40592 31096
rect 40644 31084 40650 31136
rect 40696 31133 40724 31164
rect 40954 31152 40960 31204
rect 41012 31192 41018 31204
rect 41325 31195 41383 31201
rect 41325 31192 41337 31195
rect 41012 31164 41337 31192
rect 41012 31152 41018 31164
rect 41325 31161 41337 31164
rect 41371 31192 41383 31195
rect 46860 31192 46888 31223
rect 47302 31220 47308 31232
rect 47360 31220 47366 31272
rect 41371 31164 46888 31192
rect 41371 31161 41383 31164
rect 41325 31155 41383 31161
rect 40681 31127 40739 31133
rect 40681 31093 40693 31127
rect 40727 31093 40739 31127
rect 40681 31087 40739 31093
rect 40770 31084 40776 31136
rect 40828 31124 40834 31136
rect 40865 31127 40923 31133
rect 40865 31124 40877 31127
rect 40828 31096 40877 31124
rect 40828 31084 40834 31096
rect 40865 31093 40877 31096
rect 40911 31093 40923 31127
rect 40865 31087 40923 31093
rect 42794 31084 42800 31136
rect 42852 31124 42858 31136
rect 43073 31127 43131 31133
rect 43073 31124 43085 31127
rect 42852 31096 43085 31124
rect 42852 31084 42858 31096
rect 43073 31093 43085 31096
rect 43119 31093 43131 31127
rect 43073 31087 43131 31093
rect 45094 31084 45100 31136
rect 45152 31084 45158 31136
rect 45278 31084 45284 31136
rect 45336 31084 45342 31136
rect 46937 31127 46995 31133
rect 46937 31093 46949 31127
rect 46983 31124 46995 31127
rect 47210 31124 47216 31136
rect 46983 31096 47216 31124
rect 46983 31093 46995 31096
rect 46937 31087 46995 31093
rect 47210 31084 47216 31096
rect 47268 31084 47274 31136
rect 1104 31034 78844 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 78844 31034
rect 1104 30960 78844 30982
rect 9858 30880 9864 30932
rect 9916 30920 9922 30932
rect 10965 30923 11023 30929
rect 10965 30920 10977 30923
rect 9916 30892 10977 30920
rect 9916 30880 9922 30892
rect 10965 30889 10977 30892
rect 11011 30889 11023 30923
rect 10965 30883 11023 30889
rect 12161 30923 12219 30929
rect 12161 30889 12173 30923
rect 12207 30920 12219 30923
rect 12342 30920 12348 30932
rect 12207 30892 12348 30920
rect 12207 30889 12219 30892
rect 12161 30883 12219 30889
rect 12342 30880 12348 30892
rect 12400 30880 12406 30932
rect 15378 30880 15384 30932
rect 15436 30920 15442 30932
rect 15473 30923 15531 30929
rect 15473 30920 15485 30923
rect 15436 30892 15485 30920
rect 15436 30880 15442 30892
rect 15473 30889 15485 30892
rect 15519 30889 15531 30923
rect 15473 30883 15531 30889
rect 18506 30880 18512 30932
rect 18564 30880 18570 30932
rect 29086 30880 29092 30932
rect 29144 30880 29150 30932
rect 31570 30880 31576 30932
rect 31628 30880 31634 30932
rect 36906 30880 36912 30932
rect 36964 30920 36970 30932
rect 37277 30923 37335 30929
rect 37277 30920 37289 30923
rect 36964 30892 37289 30920
rect 36964 30880 36970 30892
rect 37277 30889 37289 30892
rect 37323 30889 37335 30923
rect 37277 30883 37335 30889
rect 37366 30880 37372 30932
rect 37424 30920 37430 30932
rect 37829 30923 37887 30929
rect 37829 30920 37841 30923
rect 37424 30892 37841 30920
rect 37424 30880 37430 30892
rect 37829 30889 37841 30892
rect 37875 30889 37887 30923
rect 37829 30883 37887 30889
rect 40678 30880 40684 30932
rect 40736 30880 40742 30932
rect 41601 30923 41659 30929
rect 41601 30889 41613 30923
rect 41647 30920 41659 30923
rect 42518 30920 42524 30932
rect 41647 30892 42524 30920
rect 41647 30889 41659 30892
rect 41601 30883 41659 30889
rect 42518 30880 42524 30892
rect 42576 30880 42582 30932
rect 46750 30880 46756 30932
rect 46808 30880 46814 30932
rect 48685 30923 48743 30929
rect 48685 30920 48697 30923
rect 46860 30892 48697 30920
rect 17405 30855 17463 30861
rect 17405 30821 17417 30855
rect 17451 30852 17463 30855
rect 31389 30855 31447 30861
rect 17451 30824 17632 30852
rect 17451 30821 17463 30824
rect 17405 30815 17463 30821
rect 11333 30787 11391 30793
rect 11333 30784 11345 30787
rect 10980 30756 11345 30784
rect 10980 30725 11008 30756
rect 11333 30753 11345 30756
rect 11379 30753 11391 30787
rect 11333 30747 11391 30753
rect 11698 30744 11704 30796
rect 11756 30744 11762 30796
rect 17604 30793 17632 30824
rect 31389 30821 31401 30855
rect 31435 30852 31447 30855
rect 32122 30852 32128 30864
rect 31435 30824 32128 30852
rect 31435 30821 31447 30824
rect 31389 30815 31447 30821
rect 32122 30812 32128 30824
rect 32180 30812 32186 30864
rect 46566 30812 46572 30864
rect 46624 30852 46630 30864
rect 46860 30852 46888 30892
rect 48685 30889 48697 30892
rect 48731 30889 48743 30923
rect 48685 30883 48743 30889
rect 46624 30824 46888 30852
rect 46624 30812 46630 30824
rect 17589 30787 17647 30793
rect 17589 30753 17601 30787
rect 17635 30753 17647 30787
rect 19518 30784 19524 30796
rect 17589 30747 17647 30753
rect 18156 30756 19524 30784
rect 2041 30719 2099 30725
rect 2041 30685 2053 30719
rect 2087 30716 2099 30719
rect 2133 30719 2191 30725
rect 2133 30716 2145 30719
rect 2087 30688 2145 30716
rect 2087 30685 2099 30688
rect 2041 30679 2099 30685
rect 2133 30685 2145 30688
rect 2179 30685 2191 30719
rect 2133 30679 2191 30685
rect 10965 30719 11023 30725
rect 10965 30685 10977 30719
rect 11011 30685 11023 30719
rect 10965 30679 11023 30685
rect 11149 30719 11207 30725
rect 11149 30685 11161 30719
rect 11195 30685 11207 30719
rect 11149 30679 11207 30685
rect 11164 30648 11192 30679
rect 11238 30676 11244 30728
rect 11296 30676 11302 30728
rect 11422 30676 11428 30728
rect 11480 30676 11486 30728
rect 11793 30719 11851 30725
rect 11793 30685 11805 30719
rect 11839 30716 11851 30719
rect 12802 30716 12808 30728
rect 11839 30688 12808 30716
rect 11839 30685 11851 30688
rect 11793 30679 11851 30685
rect 12802 30676 12808 30688
rect 12860 30676 12866 30728
rect 15194 30676 15200 30728
rect 15252 30676 15258 30728
rect 15473 30719 15531 30725
rect 15473 30685 15485 30719
rect 15519 30716 15531 30719
rect 16666 30716 16672 30728
rect 15519 30688 16672 30716
rect 15519 30685 15531 30688
rect 15473 30679 15531 30685
rect 16666 30676 16672 30688
rect 16724 30676 16730 30728
rect 17126 30676 17132 30728
rect 17184 30676 17190 30728
rect 17405 30719 17463 30725
rect 17405 30685 17417 30719
rect 17451 30716 17463 30719
rect 18156 30716 18184 30756
rect 19518 30744 19524 30756
rect 19576 30744 19582 30796
rect 27338 30744 27344 30796
rect 27396 30744 27402 30796
rect 27614 30744 27620 30796
rect 27672 30744 27678 30796
rect 37476 30756 38148 30784
rect 37476 30728 37504 30756
rect 17451 30688 18184 30716
rect 18233 30719 18291 30725
rect 17451 30685 17463 30688
rect 17405 30679 17463 30685
rect 18233 30685 18245 30719
rect 18279 30716 18291 30719
rect 18325 30719 18383 30725
rect 18325 30716 18337 30719
rect 18279 30688 18337 30716
rect 18279 30685 18291 30688
rect 18233 30679 18291 30685
rect 18325 30685 18337 30688
rect 18371 30685 18383 30719
rect 18325 30679 18383 30685
rect 18414 30676 18420 30728
rect 18472 30716 18478 30728
rect 18509 30719 18567 30725
rect 18509 30716 18521 30719
rect 18472 30688 18521 30716
rect 18472 30676 18478 30688
rect 18509 30685 18521 30688
rect 18555 30685 18567 30719
rect 18509 30679 18567 30685
rect 31294 30676 31300 30728
rect 31352 30716 31358 30728
rect 31573 30719 31631 30725
rect 31573 30716 31585 30719
rect 31352 30688 31585 30716
rect 31352 30676 31358 30688
rect 31573 30685 31585 30688
rect 31619 30685 31631 30719
rect 31573 30679 31631 30685
rect 31941 30719 31999 30725
rect 31941 30685 31953 30719
rect 31987 30685 31999 30719
rect 31941 30679 31999 30685
rect 32033 30719 32091 30725
rect 32033 30685 32045 30719
rect 32079 30716 32091 30719
rect 32122 30716 32128 30728
rect 32079 30688 32128 30716
rect 32079 30685 32091 30688
rect 32033 30679 32091 30685
rect 11698 30648 11704 30660
rect 11164 30620 11704 30648
rect 11698 30608 11704 30620
rect 11756 30608 11762 30660
rect 28350 30608 28356 30660
rect 28408 30608 28414 30660
rect 934 30540 940 30592
rect 992 30580 998 30592
rect 1857 30583 1915 30589
rect 1857 30580 1869 30583
rect 992 30552 1869 30580
rect 992 30540 998 30552
rect 1857 30549 1869 30552
rect 1903 30549 1915 30583
rect 1857 30543 1915 30549
rect 15286 30540 15292 30592
rect 15344 30540 15350 30592
rect 17221 30583 17279 30589
rect 17221 30549 17233 30583
rect 17267 30580 17279 30583
rect 17954 30580 17960 30592
rect 17267 30552 17960 30580
rect 17267 30549 17279 30552
rect 17221 30543 17279 30549
rect 17954 30540 17960 30552
rect 18012 30540 18018 30592
rect 30374 30540 30380 30592
rect 30432 30580 30438 30592
rect 30653 30583 30711 30589
rect 30653 30580 30665 30583
rect 30432 30552 30665 30580
rect 30432 30540 30438 30552
rect 30653 30549 30665 30552
rect 30699 30549 30711 30583
rect 31956 30580 31984 30679
rect 32122 30676 32128 30688
rect 32180 30676 32186 30728
rect 34238 30676 34244 30728
rect 34296 30676 34302 30728
rect 37458 30676 37464 30728
rect 37516 30676 37522 30728
rect 37734 30716 37740 30728
rect 37568 30688 37740 30716
rect 32950 30608 32956 30660
rect 33008 30608 33014 30660
rect 33962 30608 33968 30660
rect 34020 30608 34026 30660
rect 36265 30651 36323 30657
rect 36265 30617 36277 30651
rect 36311 30617 36323 30651
rect 36265 30611 36323 30617
rect 32493 30583 32551 30589
rect 32493 30580 32505 30583
rect 31956 30552 32505 30580
rect 30653 30543 30711 30549
rect 32493 30549 32505 30552
rect 32539 30580 32551 30583
rect 33134 30580 33140 30592
rect 32539 30552 33140 30580
rect 32539 30549 32551 30552
rect 32493 30543 32551 30549
rect 33134 30540 33140 30552
rect 33192 30540 33198 30592
rect 36078 30540 36084 30592
rect 36136 30540 36142 30592
rect 36280 30580 36308 30611
rect 36446 30608 36452 30660
rect 36504 30648 36510 30660
rect 37568 30648 37596 30688
rect 37734 30676 37740 30688
rect 37792 30676 37798 30728
rect 37826 30676 37832 30728
rect 37884 30676 37890 30728
rect 38120 30725 38148 30756
rect 42702 30744 42708 30796
rect 42760 30784 42766 30796
rect 43349 30787 43407 30793
rect 43349 30784 43361 30787
rect 42760 30756 43361 30784
rect 42760 30744 42766 30756
rect 43349 30753 43361 30756
rect 43395 30784 43407 30787
rect 45005 30787 45063 30793
rect 45005 30784 45017 30787
rect 43395 30756 45017 30784
rect 43395 30753 43407 30756
rect 43349 30747 43407 30753
rect 45005 30753 45017 30756
rect 45051 30784 45063 30787
rect 46937 30787 46995 30793
rect 46937 30784 46949 30787
rect 45051 30756 46949 30784
rect 45051 30753 45063 30756
rect 45005 30747 45063 30753
rect 46937 30753 46949 30756
rect 46983 30753 46995 30787
rect 46937 30747 46995 30753
rect 47210 30744 47216 30796
rect 47268 30744 47274 30796
rect 38105 30719 38163 30725
rect 38105 30685 38117 30719
rect 38151 30685 38163 30719
rect 38105 30679 38163 30685
rect 40586 30676 40592 30728
rect 40644 30676 40650 30728
rect 36504 30620 37596 30648
rect 37921 30651 37979 30657
rect 36504 30608 36510 30620
rect 37921 30617 37933 30651
rect 37967 30617 37979 30651
rect 37921 30611 37979 30617
rect 36538 30580 36544 30592
rect 36280 30552 36544 30580
rect 36538 30540 36544 30552
rect 36596 30580 36602 30592
rect 37642 30580 37648 30592
rect 36596 30552 37648 30580
rect 36596 30540 36602 30552
rect 37642 30540 37648 30552
rect 37700 30540 37706 30592
rect 37734 30540 37740 30592
rect 37792 30580 37798 30592
rect 37936 30580 37964 30611
rect 40218 30608 40224 30660
rect 40276 30648 40282 30660
rect 41230 30648 41236 30660
rect 40276 30620 41236 30648
rect 40276 30608 40282 30620
rect 41230 30608 41236 30620
rect 41288 30648 41294 30660
rect 41288 30620 41906 30648
rect 41288 30608 41294 30620
rect 43070 30608 43076 30660
rect 43128 30608 43134 30660
rect 45278 30608 45284 30660
rect 45336 30608 45342 30660
rect 46934 30648 46940 30660
rect 46506 30620 46940 30648
rect 46934 30608 46940 30620
rect 46992 30608 46998 30660
rect 48438 30620 48544 30648
rect 37792 30552 37964 30580
rect 37792 30540 37798 30552
rect 43622 30540 43628 30592
rect 43680 30580 43686 30592
rect 43717 30583 43775 30589
rect 43717 30580 43729 30583
rect 43680 30552 43729 30580
rect 43680 30540 43686 30552
rect 43717 30549 43729 30552
rect 43763 30549 43775 30583
rect 43717 30543 43775 30549
rect 48222 30540 48228 30592
rect 48280 30580 48286 30592
rect 48516 30580 48544 30620
rect 48774 30580 48780 30592
rect 48280 30552 48780 30580
rect 48280 30540 48286 30552
rect 48774 30540 48780 30552
rect 48832 30540 48838 30592
rect 1104 30490 78844 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 66314 30490
rect 66366 30438 66378 30490
rect 66430 30438 66442 30490
rect 66494 30438 66506 30490
rect 66558 30438 66570 30490
rect 66622 30438 78844 30490
rect 1104 30416 78844 30438
rect 11238 30336 11244 30388
rect 11296 30376 11302 30388
rect 13081 30379 13139 30385
rect 11296 30348 12572 30376
rect 11296 30336 11302 30348
rect 11808 30249 11836 30348
rect 12437 30311 12495 30317
rect 12437 30277 12449 30311
rect 12483 30277 12495 30311
rect 12544 30308 12572 30348
rect 13081 30345 13093 30379
rect 13127 30376 13139 30379
rect 13538 30376 13544 30388
rect 13127 30348 13544 30376
rect 13127 30345 13139 30348
rect 13081 30339 13139 30345
rect 13538 30336 13544 30348
rect 13596 30336 13602 30388
rect 15194 30336 15200 30388
rect 15252 30376 15258 30388
rect 15949 30379 16007 30385
rect 15949 30376 15961 30379
rect 15252 30348 15961 30376
rect 15252 30336 15258 30348
rect 15949 30345 15961 30348
rect 15995 30345 16007 30379
rect 15949 30339 16007 30345
rect 17589 30379 17647 30385
rect 17589 30345 17601 30379
rect 17635 30376 17647 30379
rect 17954 30376 17960 30388
rect 17635 30348 17960 30376
rect 17635 30345 17647 30348
rect 17589 30339 17647 30345
rect 17954 30336 17960 30348
rect 18012 30376 18018 30388
rect 18782 30376 18788 30388
rect 18012 30348 18788 30376
rect 18012 30336 18018 30348
rect 18782 30336 18788 30348
rect 18840 30336 18846 30388
rect 39942 30376 39948 30388
rect 39408 30348 39948 30376
rect 12621 30311 12679 30317
rect 12621 30308 12633 30311
rect 12544 30280 12633 30308
rect 12437 30271 12495 30277
rect 12621 30277 12633 30280
rect 12667 30277 12679 30311
rect 12621 30271 12679 30277
rect 13265 30311 13323 30317
rect 13265 30277 13277 30311
rect 13311 30308 13323 30311
rect 14001 30311 14059 30317
rect 14001 30308 14013 30311
rect 13311 30280 14013 30308
rect 13311 30277 13323 30280
rect 13265 30271 13323 30277
rect 14001 30277 14013 30280
rect 14047 30277 14059 30311
rect 14001 30271 14059 30277
rect 2041 30243 2099 30249
rect 2041 30209 2053 30243
rect 2087 30240 2099 30243
rect 2133 30243 2191 30249
rect 2133 30240 2145 30243
rect 2087 30212 2145 30240
rect 2087 30209 2099 30212
rect 2041 30203 2099 30209
rect 2133 30209 2145 30212
rect 2179 30209 2191 30243
rect 2133 30203 2191 30209
rect 11793 30243 11851 30249
rect 11793 30209 11805 30243
rect 11839 30209 11851 30243
rect 11793 30203 11851 30209
rect 11882 30200 11888 30252
rect 11940 30240 11946 30252
rect 12452 30240 12480 30271
rect 15470 30268 15476 30320
rect 15528 30308 15534 30320
rect 15749 30311 15807 30317
rect 15749 30308 15761 30311
rect 15528 30280 15761 30308
rect 15528 30268 15534 30280
rect 15749 30277 15761 30280
rect 15795 30277 15807 30311
rect 15749 30271 15807 30277
rect 17497 30311 17555 30317
rect 17497 30277 17509 30311
rect 17543 30308 17555 30311
rect 18690 30308 18696 30320
rect 17543 30280 18696 30308
rect 17543 30277 17555 30280
rect 17497 30271 17555 30277
rect 11940 30212 12480 30240
rect 11940 30200 11946 30212
rect 12526 30200 12532 30252
rect 12584 30200 12590 30252
rect 12989 30243 13047 30249
rect 12989 30209 13001 30243
rect 13035 30209 13047 30243
rect 12989 30203 13047 30209
rect 13363 30243 13421 30249
rect 13363 30209 13375 30243
rect 13409 30240 13421 30243
rect 13409 30212 13492 30240
rect 13409 30209 13421 30212
rect 13363 30203 13421 30209
rect 13004 30172 13032 30203
rect 12084 30144 13032 30172
rect 11609 30107 11667 30113
rect 11609 30073 11621 30107
rect 11655 30104 11667 30107
rect 11698 30104 11704 30116
rect 11655 30076 11704 30104
rect 11655 30073 11667 30076
rect 11609 30067 11667 30073
rect 11698 30064 11704 30076
rect 11756 30104 11762 30116
rect 12084 30104 12112 30144
rect 11756 30076 12112 30104
rect 11756 30064 11762 30076
rect 12250 30064 12256 30116
rect 12308 30064 12314 30116
rect 12805 30107 12863 30113
rect 12805 30073 12817 30107
rect 12851 30104 12863 30107
rect 13078 30104 13084 30116
rect 12851 30076 13084 30104
rect 12851 30073 12863 30076
rect 12805 30067 12863 30073
rect 13078 30064 13084 30076
rect 13136 30064 13142 30116
rect 13354 30064 13360 30116
rect 13412 30064 13418 30116
rect 934 29996 940 30048
rect 992 30036 998 30048
rect 1857 30039 1915 30045
rect 1857 30036 1869 30039
rect 992 30008 1869 30036
rect 992 29996 998 30008
rect 1857 30005 1869 30008
rect 1903 30005 1915 30039
rect 1857 29999 1915 30005
rect 13265 30039 13323 30045
rect 13265 30005 13277 30039
rect 13311 30036 13323 30039
rect 13464 30036 13492 30212
rect 13538 30200 13544 30252
rect 13596 30240 13602 30252
rect 15194 30240 15200 30252
rect 13596 30212 15200 30240
rect 13596 30200 13602 30212
rect 15194 30200 15200 30212
rect 15252 30200 15258 30252
rect 15764 30240 15792 30271
rect 18690 30268 18696 30280
rect 18748 30268 18754 30320
rect 30653 30311 30711 30317
rect 30653 30308 30665 30311
rect 29380 30280 30665 30308
rect 16482 30240 16488 30252
rect 15764 30212 16488 30240
rect 16482 30200 16488 30212
rect 16540 30240 16546 30252
rect 17221 30243 17279 30249
rect 17221 30240 17233 30243
rect 16540 30212 17233 30240
rect 16540 30200 16546 30212
rect 17221 30209 17233 30212
rect 17267 30209 17279 30243
rect 17221 30203 17279 30209
rect 17402 30200 17408 30252
rect 17460 30200 17466 30252
rect 18414 30200 18420 30252
rect 18472 30200 18478 30252
rect 29380 30249 29408 30280
rect 30653 30277 30665 30280
rect 30699 30277 30711 30311
rect 32493 30311 32551 30317
rect 32493 30308 32505 30311
rect 30653 30271 30711 30277
rect 31588 30280 32505 30308
rect 18601 30243 18659 30249
rect 18601 30209 18613 30243
rect 18647 30240 18659 30243
rect 18785 30243 18843 30249
rect 18785 30240 18797 30243
rect 18647 30212 18797 30240
rect 18647 30209 18659 30212
rect 18601 30203 18659 30209
rect 18785 30209 18797 30212
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 29365 30243 29423 30249
rect 29365 30209 29377 30243
rect 29411 30209 29423 30243
rect 29365 30203 29423 30209
rect 29549 30243 29607 30249
rect 29549 30209 29561 30243
rect 29595 30240 29607 30243
rect 29730 30240 29736 30252
rect 29595 30212 29736 30240
rect 29595 30209 29607 30212
rect 29549 30203 29607 30209
rect 29730 30200 29736 30212
rect 29788 30240 29794 30252
rect 29825 30243 29883 30249
rect 29825 30240 29837 30243
rect 29788 30212 29837 30240
rect 29788 30200 29794 30212
rect 29825 30209 29837 30212
rect 29871 30209 29883 30243
rect 29825 30203 29883 30209
rect 30193 30243 30251 30249
rect 30193 30209 30205 30243
rect 30239 30240 30251 30243
rect 30374 30240 30380 30252
rect 30239 30212 30380 30240
rect 30239 30209 30251 30212
rect 30193 30203 30251 30209
rect 30374 30200 30380 30212
rect 30432 30200 30438 30252
rect 31588 30249 31616 30280
rect 32493 30277 32505 30280
rect 32539 30277 32551 30311
rect 32493 30271 32551 30277
rect 32950 30268 32956 30320
rect 33008 30308 33014 30320
rect 33008 30280 35006 30308
rect 33008 30268 33014 30280
rect 35986 30268 35992 30320
rect 36044 30308 36050 30320
rect 36081 30311 36139 30317
rect 36081 30308 36093 30311
rect 36044 30280 36093 30308
rect 36044 30268 36050 30280
rect 36081 30277 36093 30280
rect 36127 30277 36139 30311
rect 36081 30271 36139 30277
rect 36297 30311 36355 30317
rect 36297 30277 36309 30311
rect 36343 30308 36355 30311
rect 36633 30311 36691 30317
rect 36633 30308 36645 30311
rect 36343 30280 36645 30308
rect 36343 30277 36355 30280
rect 36297 30271 36355 30277
rect 36633 30277 36645 30280
rect 36679 30277 36691 30311
rect 36633 30271 36691 30277
rect 37369 30311 37427 30317
rect 37369 30277 37381 30311
rect 37415 30308 37427 30311
rect 37921 30311 37979 30317
rect 37921 30308 37933 30311
rect 37415 30280 37933 30308
rect 37415 30277 37427 30280
rect 37369 30271 37427 30277
rect 37921 30277 37933 30280
rect 37967 30308 37979 30311
rect 39408 30308 39436 30348
rect 39942 30336 39948 30348
rect 40000 30376 40006 30388
rect 40000 30348 40908 30376
rect 40000 30336 40006 30348
rect 37967 30280 39436 30308
rect 37967 30277 37979 30280
rect 37921 30271 37979 30277
rect 40218 30268 40224 30320
rect 40276 30268 40282 30320
rect 40681 30311 40739 30317
rect 40681 30277 40693 30311
rect 40727 30308 40739 30311
rect 40770 30308 40776 30320
rect 40727 30280 40776 30308
rect 40727 30277 40739 30280
rect 40681 30271 40739 30277
rect 40770 30268 40776 30280
rect 40828 30268 40834 30320
rect 40880 30308 40908 30348
rect 43070 30336 43076 30388
rect 43128 30336 43134 30388
rect 44361 30379 44419 30385
rect 44361 30345 44373 30379
rect 44407 30345 44419 30379
rect 44361 30339 44419 30345
rect 44085 30311 44143 30317
rect 44085 30308 44097 30311
rect 40880 30280 44097 30308
rect 44085 30277 44097 30280
rect 44131 30308 44143 30311
rect 44376 30308 44404 30339
rect 44729 30311 44787 30317
rect 44729 30308 44741 30311
rect 44131 30280 44741 30308
rect 44131 30277 44143 30280
rect 44085 30271 44143 30277
rect 44729 30277 44741 30280
rect 44775 30308 44787 30311
rect 44910 30308 44916 30320
rect 44775 30280 44916 30308
rect 44775 30277 44787 30280
rect 44729 30271 44787 30277
rect 44910 30268 44916 30280
rect 44968 30268 44974 30320
rect 31573 30243 31631 30249
rect 31573 30209 31585 30243
rect 31619 30209 31631 30243
rect 31573 30203 31631 30209
rect 32122 30200 32128 30252
rect 32180 30200 32186 30252
rect 32309 30243 32367 30249
rect 32309 30209 32321 30243
rect 32355 30209 32367 30243
rect 32309 30203 32367 30209
rect 14550 30132 14556 30184
rect 14608 30132 14614 30184
rect 19058 30132 19064 30184
rect 19116 30172 19122 30184
rect 19337 30175 19395 30181
rect 19337 30172 19349 30175
rect 19116 30144 19349 30172
rect 19116 30132 19122 30144
rect 19337 30141 19349 30144
rect 19383 30141 19395 30175
rect 19337 30135 19395 30141
rect 29641 30175 29699 30181
rect 29641 30141 29653 30175
rect 29687 30172 29699 30175
rect 31205 30175 31263 30181
rect 31205 30172 31217 30175
rect 29687 30144 31217 30172
rect 29687 30141 29699 30144
rect 29641 30135 29699 30141
rect 31205 30141 31217 30144
rect 31251 30172 31263 30175
rect 31294 30172 31300 30184
rect 31251 30144 31300 30172
rect 31251 30141 31263 30144
rect 31205 30135 31263 30141
rect 31294 30132 31300 30144
rect 31352 30132 31358 30184
rect 31665 30175 31723 30181
rect 31665 30141 31677 30175
rect 31711 30172 31723 30175
rect 32217 30175 32275 30181
rect 32217 30172 32229 30175
rect 31711 30144 32229 30172
rect 31711 30141 31723 30144
rect 31665 30135 31723 30141
rect 32217 30141 32229 30144
rect 32263 30141 32275 30175
rect 32217 30135 32275 30141
rect 16117 30107 16175 30113
rect 16117 30073 16129 30107
rect 16163 30104 16175 30107
rect 17126 30104 17132 30116
rect 16163 30076 17132 30104
rect 16163 30073 16175 30076
rect 16117 30067 16175 30073
rect 17126 30064 17132 30076
rect 17184 30064 17190 30116
rect 28350 30064 28356 30116
rect 28408 30104 28414 30116
rect 30009 30107 30067 30113
rect 28408 30076 29684 30104
rect 28408 30064 28414 30076
rect 13311 30008 13492 30036
rect 13311 30005 13323 30008
rect 13265 29999 13323 30005
rect 15286 29996 15292 30048
rect 15344 30036 15350 30048
rect 15838 30036 15844 30048
rect 15344 30008 15844 30036
rect 15344 29996 15350 30008
rect 15838 29996 15844 30008
rect 15896 30036 15902 30048
rect 15933 30039 15991 30045
rect 15933 30036 15945 30039
rect 15896 30008 15945 30036
rect 15896 29996 15902 30008
rect 15933 30005 15945 30008
rect 15979 30005 15991 30039
rect 15933 29999 15991 30005
rect 17678 29996 17684 30048
rect 17736 30036 17742 30048
rect 17773 30039 17831 30045
rect 17773 30036 17785 30039
rect 17736 30008 17785 30036
rect 17736 29996 17742 30008
rect 17773 30005 17785 30008
rect 17819 30005 17831 30039
rect 17773 29999 17831 30005
rect 18417 30039 18475 30045
rect 18417 30005 18429 30039
rect 18463 30036 18475 30039
rect 19242 30036 19248 30048
rect 18463 30008 19248 30036
rect 18463 30005 18475 30008
rect 18417 29999 18475 30005
rect 19242 29996 19248 30008
rect 19300 29996 19306 30048
rect 29546 29996 29552 30048
rect 29604 29996 29610 30048
rect 29656 30036 29684 30076
rect 30009 30073 30021 30107
rect 30055 30104 30067 30107
rect 32324 30104 32352 30203
rect 33134 30200 33140 30252
rect 33192 30200 33198 30252
rect 34238 30200 34244 30252
rect 34296 30200 34302 30252
rect 36538 30200 36544 30252
rect 36596 30200 36602 30252
rect 36725 30243 36783 30249
rect 36725 30209 36737 30243
rect 36771 30209 36783 30243
rect 36725 30203 36783 30209
rect 34514 30132 34520 30184
rect 34572 30132 34578 30184
rect 36446 30172 36452 30184
rect 36004 30144 36452 30172
rect 30055 30076 31064 30104
rect 30055 30073 30067 30076
rect 30009 30067 30067 30073
rect 30282 30036 30288 30048
rect 29656 30008 30288 30036
rect 30282 29996 30288 30008
rect 30340 30036 30346 30048
rect 30469 30039 30527 30045
rect 30469 30036 30481 30039
rect 30340 30008 30481 30036
rect 30340 29996 30346 30008
rect 30469 30005 30481 30008
rect 30515 30005 30527 30039
rect 31036 30036 31064 30076
rect 31726 30076 32352 30104
rect 31726 30048 31754 30076
rect 31726 30036 31760 30048
rect 31036 30008 31760 30036
rect 30469 29999 30527 30005
rect 31754 29996 31760 30008
rect 31812 29996 31818 30048
rect 31849 30039 31907 30045
rect 31849 30005 31861 30039
rect 31895 30036 31907 30039
rect 33962 30036 33968 30048
rect 31895 30008 33968 30036
rect 31895 30005 31907 30008
rect 31849 29999 31907 30005
rect 33962 29996 33968 30008
rect 34020 29996 34026 30048
rect 35894 29996 35900 30048
rect 35952 30036 35958 30048
rect 36004 30045 36032 30144
rect 36446 30132 36452 30144
rect 36504 30172 36510 30184
rect 36740 30172 36768 30203
rect 42794 30200 42800 30252
rect 42852 30200 42858 30252
rect 42886 30200 42892 30252
rect 42944 30200 42950 30252
rect 43622 30200 43628 30252
rect 43680 30200 43686 30252
rect 44545 30243 44603 30249
rect 44545 30209 44557 30243
rect 44591 30240 44603 30243
rect 44818 30240 44824 30252
rect 44591 30212 44824 30240
rect 44591 30209 44603 30212
rect 44545 30203 44603 30209
rect 44818 30200 44824 30212
rect 44876 30200 44882 30252
rect 36504 30144 36768 30172
rect 39209 30175 39267 30181
rect 36504 30132 36510 30144
rect 39209 30141 39221 30175
rect 39255 30172 39267 30175
rect 40586 30172 40592 30184
rect 39255 30144 40592 30172
rect 39255 30141 39267 30144
rect 39209 30135 39267 30141
rect 40586 30132 40592 30144
rect 40644 30132 40650 30184
rect 40957 30175 41015 30181
rect 40957 30141 40969 30175
rect 41003 30141 41015 30175
rect 40957 30135 41015 30141
rect 40972 30048 41000 30135
rect 42426 30132 42432 30184
rect 42484 30132 42490 30184
rect 43438 30132 43444 30184
rect 43496 30132 43502 30184
rect 35989 30039 36047 30045
rect 35989 30036 36001 30039
rect 35952 30008 36001 30036
rect 35952 29996 35958 30008
rect 35989 30005 36001 30008
rect 36035 30005 36047 30039
rect 35989 29999 36047 30005
rect 36078 29996 36084 30048
rect 36136 30036 36142 30048
rect 36265 30039 36323 30045
rect 36265 30036 36277 30039
rect 36136 30008 36277 30036
rect 36136 29996 36142 30008
rect 36265 30005 36277 30008
rect 36311 30005 36323 30039
rect 36265 29999 36323 30005
rect 36354 29996 36360 30048
rect 36412 30036 36418 30048
rect 36449 30039 36507 30045
rect 36449 30036 36461 30039
rect 36412 30008 36461 30036
rect 36412 29996 36418 30008
rect 36449 30005 36461 30008
rect 36495 30005 36507 30039
rect 36449 29999 36507 30005
rect 37274 29996 37280 30048
rect 37332 30036 37338 30048
rect 37461 30039 37519 30045
rect 37461 30036 37473 30039
rect 37332 30008 37473 30036
rect 37332 29996 37338 30008
rect 37461 30005 37473 30008
rect 37507 30005 37519 30039
rect 37461 29999 37519 30005
rect 38654 29996 38660 30048
rect 38712 30036 38718 30048
rect 40954 30036 40960 30048
rect 38712 30008 40960 30036
rect 38712 29996 38718 30008
rect 40954 29996 40960 30008
rect 41012 29996 41018 30048
rect 43806 29996 43812 30048
rect 43864 29996 43870 30048
rect 44818 29996 44824 30048
rect 44876 29996 44882 30048
rect 46934 29996 46940 30048
rect 46992 30036 46998 30048
rect 48222 30036 48228 30048
rect 46992 30008 48228 30036
rect 46992 29996 46998 30008
rect 48222 29996 48228 30008
rect 48280 29996 48286 30048
rect 1104 29946 78844 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 78844 29946
rect 1104 29872 78844 29894
rect 11606 29792 11612 29844
rect 11664 29792 11670 29844
rect 15470 29792 15476 29844
rect 15528 29792 15534 29844
rect 15838 29792 15844 29844
rect 15896 29792 15902 29844
rect 16482 29792 16488 29844
rect 16540 29832 16546 29844
rect 17681 29835 17739 29841
rect 17681 29832 17693 29835
rect 16540 29804 17693 29832
rect 16540 29792 16546 29804
rect 17681 29801 17693 29804
rect 17727 29832 17739 29835
rect 17770 29832 17776 29844
rect 17727 29804 17776 29832
rect 17727 29801 17739 29804
rect 17681 29795 17739 29801
rect 17770 29792 17776 29804
rect 17828 29792 17834 29844
rect 17865 29835 17923 29841
rect 17865 29801 17877 29835
rect 17911 29832 17923 29835
rect 18414 29832 18420 29844
rect 17911 29804 18420 29832
rect 17911 29801 17923 29804
rect 17865 29795 17923 29801
rect 18414 29792 18420 29804
rect 18472 29792 18478 29844
rect 18782 29792 18788 29844
rect 18840 29792 18846 29844
rect 20254 29792 20260 29844
rect 20312 29832 20318 29844
rect 22281 29835 22339 29841
rect 22281 29832 22293 29835
rect 20312 29804 22293 29832
rect 20312 29792 20318 29804
rect 22281 29801 22293 29804
rect 22327 29832 22339 29835
rect 22370 29832 22376 29844
rect 22327 29804 22376 29832
rect 22327 29801 22339 29804
rect 22281 29795 22339 29801
rect 22370 29792 22376 29804
rect 22428 29792 22434 29844
rect 31294 29792 31300 29844
rect 31352 29792 31358 29844
rect 34514 29792 34520 29844
rect 34572 29832 34578 29844
rect 34701 29835 34759 29841
rect 34701 29832 34713 29835
rect 34572 29804 34713 29832
rect 34572 29792 34578 29804
rect 34701 29801 34713 29804
rect 34747 29801 34759 29835
rect 34701 29795 34759 29801
rect 37642 29792 37648 29844
rect 37700 29832 37706 29844
rect 37737 29835 37795 29841
rect 37737 29832 37749 29835
rect 37700 29804 37749 29832
rect 37700 29792 37706 29804
rect 37737 29801 37749 29804
rect 37783 29801 37795 29835
rect 37737 29795 37795 29801
rect 18601 29767 18659 29773
rect 15304 29736 17540 29764
rect 8941 29699 8999 29705
rect 8941 29665 8953 29699
rect 8987 29696 8999 29699
rect 9674 29696 9680 29708
rect 8987 29668 9680 29696
rect 8987 29665 8999 29668
rect 8941 29659 8999 29665
rect 9674 29656 9680 29668
rect 9732 29696 9738 29708
rect 10226 29696 10232 29708
rect 9732 29668 10232 29696
rect 9732 29656 9738 29668
rect 10226 29656 10232 29668
rect 10284 29656 10290 29708
rect 10689 29699 10747 29705
rect 10689 29665 10701 29699
rect 10735 29696 10747 29699
rect 11146 29696 11152 29708
rect 10735 29668 11152 29696
rect 10735 29665 10747 29668
rect 10689 29659 10747 29665
rect 11146 29656 11152 29668
rect 11204 29696 11210 29708
rect 15304 29705 15332 29736
rect 11333 29699 11391 29705
rect 11333 29696 11345 29699
rect 11204 29668 11345 29696
rect 11204 29656 11210 29668
rect 11333 29665 11345 29668
rect 11379 29665 11391 29699
rect 11333 29659 11391 29665
rect 15289 29699 15347 29705
rect 15289 29665 15301 29699
rect 15335 29665 15347 29699
rect 17402 29696 17408 29708
rect 15289 29659 15347 29665
rect 16040 29668 17408 29696
rect 14642 29588 14648 29640
rect 14700 29628 14706 29640
rect 15105 29631 15163 29637
rect 15105 29628 15117 29631
rect 14700 29600 15117 29628
rect 14700 29588 14706 29600
rect 15105 29597 15117 29600
rect 15151 29597 15163 29631
rect 15105 29591 15163 29597
rect 15565 29631 15623 29637
rect 15565 29597 15577 29631
rect 15611 29628 15623 29631
rect 15838 29628 15844 29640
rect 15611 29600 15844 29628
rect 15611 29597 15623 29600
rect 15565 29591 15623 29597
rect 15838 29588 15844 29600
rect 15896 29588 15902 29640
rect 16040 29637 16068 29668
rect 17402 29656 17408 29668
rect 17460 29656 17466 29708
rect 17512 29696 17540 29736
rect 18601 29733 18613 29767
rect 18647 29733 18659 29767
rect 20272 29764 20300 29792
rect 18601 29727 18659 29733
rect 18892 29736 20300 29764
rect 34885 29767 34943 29773
rect 18616 29696 18644 29727
rect 17512 29668 18644 29696
rect 16025 29631 16083 29637
rect 16025 29597 16037 29631
rect 16071 29597 16083 29631
rect 16025 29591 16083 29597
rect 16209 29631 16267 29637
rect 16209 29597 16221 29631
rect 16255 29597 16267 29631
rect 18325 29631 18383 29637
rect 18325 29628 18337 29631
rect 16209 29591 16267 29597
rect 17880 29600 18337 29628
rect 9214 29520 9220 29572
rect 9272 29520 9278 29572
rect 11606 29560 11612 29572
rect 10442 29532 11612 29560
rect 11606 29520 11612 29532
rect 11664 29520 11670 29572
rect 16224 29560 16252 29591
rect 16298 29560 16304 29572
rect 16224 29532 16304 29560
rect 16298 29520 16304 29532
rect 16356 29560 16362 29572
rect 17497 29563 17555 29569
rect 17497 29560 17509 29563
rect 16356 29532 17509 29560
rect 16356 29520 16362 29532
rect 17497 29529 17509 29532
rect 17543 29529 17555 29563
rect 17497 29523 17555 29529
rect 2038 29452 2044 29504
rect 2096 29452 2102 29504
rect 10778 29452 10784 29504
rect 10836 29452 10842 29504
rect 14550 29452 14556 29504
rect 14608 29492 14614 29504
rect 14921 29495 14979 29501
rect 14921 29492 14933 29495
rect 14608 29464 14933 29492
rect 14608 29452 14614 29464
rect 14921 29461 14933 29464
rect 14967 29461 14979 29495
rect 17512 29492 17540 29523
rect 17678 29520 17684 29572
rect 17736 29569 17742 29572
rect 17736 29563 17760 29569
rect 17748 29560 17760 29563
rect 17880 29560 17908 29600
rect 18325 29597 18337 29600
rect 18371 29597 18383 29631
rect 18325 29591 18383 29597
rect 18690 29588 18696 29640
rect 18748 29628 18754 29640
rect 18892 29637 18920 29736
rect 34885 29733 34897 29767
rect 34931 29764 34943 29767
rect 35986 29764 35992 29776
rect 34931 29736 35992 29764
rect 34931 29733 34943 29736
rect 34885 29727 34943 29733
rect 35986 29724 35992 29736
rect 36044 29724 36050 29776
rect 19978 29696 19984 29708
rect 19444 29668 19984 29696
rect 18785 29631 18843 29637
rect 18785 29628 18797 29631
rect 18748 29600 18797 29628
rect 18748 29588 18754 29600
rect 18785 29597 18797 29600
rect 18831 29597 18843 29631
rect 18785 29591 18843 29597
rect 18877 29631 18935 29637
rect 18877 29597 18889 29631
rect 18923 29597 18935 29631
rect 18877 29591 18935 29597
rect 19058 29588 19064 29640
rect 19116 29588 19122 29640
rect 19242 29588 19248 29640
rect 19300 29588 19306 29640
rect 19444 29637 19472 29668
rect 19978 29656 19984 29668
rect 20036 29656 20042 29708
rect 20441 29699 20499 29705
rect 20441 29665 20453 29699
rect 20487 29665 20499 29699
rect 20441 29659 20499 29665
rect 20533 29699 20591 29705
rect 20533 29665 20545 29699
rect 20579 29696 20591 29699
rect 20806 29696 20812 29708
rect 20579 29668 20812 29696
rect 20579 29665 20591 29668
rect 20533 29659 20591 29665
rect 19429 29631 19487 29637
rect 19429 29597 19441 29631
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 17748 29532 17908 29560
rect 17748 29529 17760 29532
rect 17736 29523 17760 29529
rect 17736 29520 17742 29523
rect 17954 29520 17960 29572
rect 18012 29520 18018 29572
rect 18141 29563 18199 29569
rect 18141 29529 18153 29563
rect 18187 29560 18199 29563
rect 19076 29560 19104 29588
rect 19444 29560 19472 29591
rect 20070 29588 20076 29640
rect 20128 29588 20134 29640
rect 18187 29532 19104 29560
rect 19260 29532 19472 29560
rect 20456 29560 20484 29659
rect 20806 29656 20812 29668
rect 20864 29696 20870 29708
rect 21450 29696 21456 29708
rect 20864 29668 21456 29696
rect 20864 29656 20870 29668
rect 21450 29656 21456 29668
rect 21508 29656 21514 29708
rect 29549 29699 29607 29705
rect 29549 29665 29561 29699
rect 29595 29696 29607 29699
rect 30190 29696 30196 29708
rect 29595 29668 30196 29696
rect 29595 29665 29607 29668
rect 29549 29659 29607 29665
rect 30190 29656 30196 29668
rect 30248 29656 30254 29708
rect 32122 29656 32128 29708
rect 32180 29696 32186 29708
rect 32401 29699 32459 29705
rect 32401 29696 32413 29699
rect 32180 29668 32413 29696
rect 32180 29656 32186 29668
rect 32401 29665 32413 29668
rect 32447 29665 32459 29699
rect 32401 29659 32459 29665
rect 35161 29699 35219 29705
rect 35161 29665 35173 29699
rect 35207 29696 35219 29699
rect 35894 29696 35900 29708
rect 35207 29668 35900 29696
rect 35207 29665 35219 29668
rect 35161 29659 35219 29665
rect 35894 29656 35900 29668
rect 35952 29656 35958 29708
rect 36265 29699 36323 29705
rect 36265 29665 36277 29699
rect 36311 29696 36323 29699
rect 36354 29696 36360 29708
rect 36311 29668 36360 29696
rect 36311 29665 36323 29668
rect 36265 29659 36323 29665
rect 36354 29656 36360 29668
rect 36412 29656 36418 29708
rect 40954 29656 40960 29708
rect 41012 29696 41018 29708
rect 42245 29699 42303 29705
rect 42245 29696 42257 29699
rect 41012 29668 42257 29696
rect 41012 29656 41018 29668
rect 42245 29665 42257 29668
rect 42291 29665 42303 29699
rect 42245 29659 42303 29665
rect 34238 29588 34244 29640
rect 34296 29628 34302 29640
rect 35986 29628 35992 29640
rect 34296 29600 35992 29628
rect 34296 29588 34302 29600
rect 35986 29588 35992 29600
rect 36044 29588 36050 29640
rect 43806 29628 43812 29640
rect 43654 29614 43812 29628
rect 43640 29600 43812 29614
rect 20809 29563 20867 29569
rect 20809 29560 20821 29563
rect 20456 29532 20821 29560
rect 18187 29529 18199 29532
rect 18141 29523 18199 29529
rect 17972 29492 18000 29520
rect 17512 29464 18000 29492
rect 14921 29455 14979 29461
rect 18046 29452 18052 29504
rect 18104 29492 18110 29504
rect 18233 29495 18291 29501
rect 18233 29492 18245 29495
rect 18104 29464 18245 29492
rect 18104 29452 18110 29464
rect 18233 29461 18245 29464
rect 18279 29461 18291 29495
rect 18233 29455 18291 29461
rect 18509 29495 18567 29501
rect 18509 29461 18521 29495
rect 18555 29492 18567 29495
rect 19260 29492 19288 29532
rect 20809 29529 20821 29532
rect 20855 29529 20867 29563
rect 28350 29560 28356 29572
rect 22034 29532 28356 29560
rect 20809 29523 20867 29529
rect 28350 29520 28356 29532
rect 28408 29520 28414 29572
rect 29825 29563 29883 29569
rect 29825 29529 29837 29563
rect 29871 29560 29883 29563
rect 30098 29560 30104 29572
rect 29871 29532 30104 29560
rect 29871 29529 29883 29532
rect 29825 29523 29883 29529
rect 30098 29520 30104 29532
rect 30156 29520 30162 29572
rect 30282 29520 30288 29572
rect 30340 29520 30346 29572
rect 32950 29520 32956 29572
rect 33008 29560 33014 29572
rect 37829 29563 37887 29569
rect 33008 29532 36754 29560
rect 33008 29520 33014 29532
rect 18555 29464 19288 29492
rect 19337 29495 19395 29501
rect 18555 29461 18567 29464
rect 18509 29455 18567 29461
rect 19337 29461 19349 29495
rect 19383 29492 19395 29495
rect 20438 29492 20444 29504
rect 19383 29464 20444 29492
rect 19383 29461 19395 29464
rect 19337 29455 19395 29461
rect 20438 29452 20444 29464
rect 20496 29452 20502 29504
rect 31570 29452 31576 29504
rect 31628 29492 31634 29504
rect 31849 29495 31907 29501
rect 31849 29492 31861 29495
rect 31628 29464 31861 29492
rect 31628 29452 31634 29464
rect 31849 29461 31861 29464
rect 31895 29461 31907 29495
rect 36648 29492 36676 29532
rect 37829 29529 37841 29563
rect 37875 29529 37887 29563
rect 37829 29523 37887 29529
rect 38565 29563 38623 29569
rect 38565 29529 38577 29563
rect 38611 29560 38623 29563
rect 38654 29560 38660 29572
rect 38611 29532 38660 29560
rect 38611 29529 38623 29532
rect 38565 29523 38623 29529
rect 37274 29492 37280 29504
rect 36648 29464 37280 29492
rect 31849 29455 31907 29461
rect 37274 29452 37280 29464
rect 37332 29452 37338 29504
rect 37844 29492 37872 29523
rect 38654 29520 38660 29532
rect 38712 29520 38718 29572
rect 42521 29563 42579 29569
rect 42521 29529 42533 29563
rect 42567 29560 42579 29563
rect 42610 29560 42616 29572
rect 42567 29532 42616 29560
rect 42567 29529 42579 29532
rect 42521 29523 42579 29529
rect 42610 29520 42616 29532
rect 42668 29520 42674 29572
rect 38470 29492 38476 29504
rect 37844 29464 38476 29492
rect 38470 29452 38476 29464
rect 38528 29492 38534 29504
rect 38838 29492 38844 29504
rect 38528 29464 38844 29492
rect 38528 29452 38534 29464
rect 38838 29452 38844 29464
rect 38896 29452 38902 29504
rect 40218 29452 40224 29504
rect 40276 29492 40282 29504
rect 43640 29492 43668 29600
rect 43806 29588 43812 29600
rect 43864 29588 43870 29640
rect 44269 29563 44327 29569
rect 44269 29529 44281 29563
rect 44315 29560 44327 29563
rect 44358 29560 44364 29572
rect 44315 29532 44364 29560
rect 44315 29529 44327 29532
rect 44269 29523 44327 29529
rect 44358 29520 44364 29532
rect 44416 29520 44422 29572
rect 40276 29464 43668 29492
rect 40276 29452 40282 29464
rect 1104 29402 78844 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 66314 29402
rect 66366 29350 66378 29402
rect 66430 29350 66442 29402
rect 66494 29350 66506 29402
rect 66558 29350 66570 29402
rect 66622 29350 78844 29402
rect 1104 29328 78844 29350
rect 1302 29248 1308 29300
rect 1360 29288 1366 29300
rect 1857 29291 1915 29297
rect 1857 29288 1869 29291
rect 1360 29260 1869 29288
rect 1360 29248 1366 29260
rect 1857 29257 1869 29260
rect 1903 29257 1915 29291
rect 1857 29251 1915 29257
rect 10781 29291 10839 29297
rect 10781 29257 10793 29291
rect 10827 29257 10839 29291
rect 10781 29251 10839 29257
rect 10796 29220 10824 29251
rect 11146 29248 11152 29300
rect 11204 29248 11210 29300
rect 12161 29291 12219 29297
rect 12161 29257 12173 29291
rect 12207 29288 12219 29291
rect 13354 29288 13360 29300
rect 12207 29260 13360 29288
rect 12207 29257 12219 29260
rect 12161 29251 12219 29257
rect 13354 29248 13360 29260
rect 13412 29248 13418 29300
rect 14734 29248 14740 29300
rect 14792 29248 14798 29300
rect 18969 29291 19027 29297
rect 18969 29257 18981 29291
rect 19015 29288 19027 29291
rect 19058 29288 19064 29300
rect 19015 29260 19064 29288
rect 19015 29257 19027 29260
rect 18969 29251 19027 29257
rect 19058 29248 19064 29260
rect 19116 29248 19122 29300
rect 20070 29248 20076 29300
rect 20128 29288 20134 29300
rect 21821 29291 21879 29297
rect 21821 29288 21833 29291
rect 20128 29260 21833 29288
rect 20128 29248 20134 29260
rect 21821 29257 21833 29260
rect 21867 29257 21879 29291
rect 21821 29251 21879 29257
rect 30098 29248 30104 29300
rect 30156 29248 30162 29300
rect 32122 29248 32128 29300
rect 32180 29248 32186 29300
rect 39390 29248 39396 29300
rect 39448 29248 39454 29300
rect 42610 29248 42616 29300
rect 42668 29248 42674 29300
rect 42978 29288 42984 29300
rect 42939 29260 42984 29288
rect 42978 29248 42984 29260
rect 43036 29288 43042 29300
rect 44358 29288 44364 29300
rect 43036 29260 44364 29288
rect 43036 29248 43042 29260
rect 44358 29248 44364 29260
rect 44416 29248 44422 29300
rect 11164 29220 11192 29248
rect 13173 29223 13231 29229
rect 10796 29192 11008 29220
rect 11164 29192 12020 29220
rect 2038 29112 2044 29164
rect 2096 29112 2102 29164
rect 10689 29155 10747 29161
rect 10689 29121 10701 29155
rect 10735 29152 10747 29155
rect 10778 29152 10784 29164
rect 10735 29124 10784 29152
rect 10735 29121 10747 29124
rect 10689 29115 10747 29121
rect 10778 29112 10784 29124
rect 10836 29112 10842 29164
rect 10870 29112 10876 29164
rect 10928 29112 10934 29164
rect 10980 29161 11008 29192
rect 10965 29155 11023 29161
rect 10965 29121 10977 29155
rect 11011 29121 11023 29155
rect 10965 29115 11023 29121
rect 11149 29155 11207 29161
rect 11149 29121 11161 29155
rect 11195 29152 11207 29155
rect 11238 29152 11244 29164
rect 11195 29124 11244 29152
rect 11195 29121 11207 29124
rect 11149 29115 11207 29121
rect 11238 29112 11244 29124
rect 11296 29112 11302 29164
rect 11330 29112 11336 29164
rect 11388 29152 11394 29164
rect 11517 29155 11575 29161
rect 11517 29152 11529 29155
rect 11388 29124 11529 29152
rect 11388 29112 11394 29124
rect 11517 29121 11529 29124
rect 11563 29121 11575 29155
rect 11517 29115 11575 29121
rect 11882 29112 11888 29164
rect 11940 29112 11946 29164
rect 11992 29161 12020 29192
rect 13173 29189 13185 29223
rect 13219 29220 13231 29223
rect 13262 29220 13268 29232
rect 13219 29192 13268 29220
rect 13219 29189 13231 29192
rect 13173 29183 13231 29189
rect 13262 29180 13268 29192
rect 13320 29180 13326 29232
rect 14752 29220 14780 29248
rect 14398 29192 14780 29220
rect 20438 29180 20444 29232
rect 20496 29180 20502 29232
rect 32950 29180 32956 29232
rect 33008 29180 33014 29232
rect 38654 29220 38660 29232
rect 38028 29192 38660 29220
rect 11977 29155 12035 29161
rect 11977 29121 11989 29155
rect 12023 29121 12035 29155
rect 11977 29115 12035 29121
rect 15194 29112 15200 29164
rect 15252 29152 15258 29164
rect 15381 29155 15439 29161
rect 15381 29152 15393 29155
rect 15252 29124 15393 29152
rect 15252 29112 15258 29124
rect 15381 29121 15393 29124
rect 15427 29121 15439 29155
rect 15381 29115 15439 29121
rect 15565 29155 15623 29161
rect 15565 29121 15577 29155
rect 15611 29152 15623 29155
rect 15838 29152 15844 29164
rect 15611 29124 15844 29152
rect 15611 29121 15623 29124
rect 15565 29115 15623 29121
rect 2130 29044 2136 29096
rect 2188 29044 2194 29096
rect 9214 29044 9220 29096
rect 9272 29084 9278 29096
rect 11057 29087 11115 29093
rect 11057 29084 11069 29087
rect 9272 29056 11069 29084
rect 9272 29044 9278 29056
rect 11057 29053 11069 29056
rect 11103 29053 11115 29087
rect 12897 29087 12955 29093
rect 12897 29084 12909 29087
rect 11057 29047 11115 29053
rect 12406 29056 12909 29084
rect 10226 28976 10232 29028
rect 10284 29016 10290 29028
rect 12406 29016 12434 29056
rect 12897 29053 12909 29056
rect 12943 29084 12955 29087
rect 13262 29084 13268 29096
rect 12943 29056 13268 29084
rect 12943 29053 12955 29056
rect 12897 29047 12955 29053
rect 13262 29044 13268 29056
rect 13320 29044 13326 29096
rect 14642 29044 14648 29096
rect 14700 29044 14706 29096
rect 15396 29084 15424 29115
rect 15838 29112 15844 29124
rect 15896 29112 15902 29164
rect 16666 29112 16672 29164
rect 16724 29112 16730 29164
rect 19334 29112 19340 29164
rect 19392 29112 19398 29164
rect 20717 29155 20775 29161
rect 20717 29121 20729 29155
rect 20763 29152 20775 29155
rect 20806 29152 20812 29164
rect 20763 29124 20812 29152
rect 20763 29121 20775 29124
rect 20717 29115 20775 29121
rect 20806 29112 20812 29124
rect 20864 29112 20870 29164
rect 22370 29112 22376 29164
rect 22428 29112 22434 29164
rect 29546 29112 29552 29164
rect 29604 29152 29610 29164
rect 30009 29155 30067 29161
rect 30009 29152 30021 29155
rect 29604 29124 30021 29152
rect 29604 29112 29610 29124
rect 30009 29121 30021 29124
rect 30055 29121 30067 29155
rect 30009 29115 30067 29121
rect 30193 29155 30251 29161
rect 30193 29121 30205 29155
rect 30239 29121 30251 29155
rect 30193 29115 30251 29121
rect 16482 29084 16488 29096
rect 15396 29056 16488 29084
rect 16482 29044 16488 29056
rect 16540 29044 16546 29096
rect 19352 29084 19380 29112
rect 20346 29084 20352 29096
rect 19352 29056 20352 29084
rect 20346 29044 20352 29056
rect 20404 29084 20410 29096
rect 20901 29087 20959 29093
rect 20901 29084 20913 29087
rect 20404 29056 20913 29084
rect 20404 29044 20410 29056
rect 20901 29053 20913 29056
rect 20947 29084 20959 29087
rect 30208 29084 30236 29115
rect 31570 29112 31576 29164
rect 31628 29112 31634 29164
rect 31754 29152 31760 29164
rect 31680 29124 31760 29152
rect 31680 29093 31708 29124
rect 31754 29112 31760 29124
rect 31812 29112 31818 29164
rect 33873 29155 33931 29161
rect 33873 29121 33885 29155
rect 33919 29152 33931 29155
rect 34238 29152 34244 29164
rect 33919 29124 34244 29152
rect 33919 29121 33931 29124
rect 33873 29115 33931 29121
rect 34238 29112 34244 29124
rect 34296 29112 34302 29164
rect 31665 29087 31723 29093
rect 31665 29084 31677 29087
rect 20947 29056 22094 29084
rect 30208 29056 31677 29084
rect 20947 29053 20959 29056
rect 20901 29047 20959 29053
rect 10284 28988 12434 29016
rect 10284 28976 10290 28988
rect 15286 28976 15292 29028
rect 15344 29016 15350 29028
rect 16298 29016 16304 29028
rect 15344 28988 16304 29016
rect 15344 28976 15350 28988
rect 16298 28976 16304 28988
rect 16356 28976 16362 29028
rect 22066 29016 22094 29056
rect 31665 29053 31677 29056
rect 31711 29053 31723 29087
rect 31665 29047 31723 29053
rect 31941 29087 31999 29093
rect 31941 29053 31953 29087
rect 31987 29084 31999 29087
rect 33597 29087 33655 29093
rect 33597 29084 33609 29087
rect 31987 29056 33609 29084
rect 31987 29053 31999 29056
rect 31941 29047 31999 29053
rect 33597 29053 33609 29056
rect 33643 29053 33655 29087
rect 33597 29047 33655 29053
rect 35986 29044 35992 29096
rect 36044 29084 36050 29096
rect 38028 29093 38056 29192
rect 38654 29180 38660 29192
rect 38712 29180 38718 29232
rect 38286 29161 38292 29164
rect 38280 29115 38292 29161
rect 38286 29112 38292 29115
rect 38344 29112 38350 29164
rect 39408 29152 39436 29248
rect 41138 29180 41144 29232
rect 41196 29220 41202 29232
rect 41417 29223 41475 29229
rect 41417 29220 41429 29223
rect 41196 29192 41429 29220
rect 41196 29180 41202 29192
rect 41417 29189 41429 29192
rect 41463 29220 41475 29223
rect 43438 29220 43444 29232
rect 41463 29192 43444 29220
rect 41463 29189 41475 29192
rect 41417 29183 41475 29189
rect 40037 29155 40095 29161
rect 40037 29152 40049 29155
rect 39408 29124 40049 29152
rect 40037 29121 40049 29124
rect 40083 29121 40095 29155
rect 40037 29115 40095 29121
rect 40862 29112 40868 29164
rect 40920 29112 40926 29164
rect 40957 29155 41015 29161
rect 40957 29121 40969 29155
rect 41003 29152 41015 29155
rect 42702 29152 42708 29164
rect 41003 29124 42708 29152
rect 41003 29121 41015 29124
rect 40957 29115 41015 29121
rect 42702 29112 42708 29124
rect 42760 29112 42766 29164
rect 38013 29087 38071 29093
rect 38013 29084 38025 29087
rect 36044 29056 38025 29084
rect 36044 29044 36050 29056
rect 38013 29053 38025 29056
rect 38059 29053 38071 29087
rect 38013 29047 38071 29053
rect 41138 29044 41144 29096
rect 41196 29044 41202 29096
rect 43070 29044 43076 29096
rect 43128 29044 43134 29096
rect 43272 29093 43300 29192
rect 43438 29180 43444 29192
rect 43496 29220 43502 29232
rect 43533 29223 43591 29229
rect 43533 29220 43545 29223
rect 43496 29192 43545 29220
rect 43496 29180 43502 29192
rect 43533 29189 43545 29192
rect 43579 29220 43591 29223
rect 47670 29220 47676 29232
rect 43579 29192 47676 29220
rect 43579 29189 43591 29192
rect 43533 29183 43591 29189
rect 47670 29180 47676 29192
rect 47728 29180 47734 29232
rect 44085 29155 44143 29161
rect 44085 29121 44097 29155
rect 44131 29121 44143 29155
rect 44266 29152 44272 29164
rect 44085 29115 44143 29121
rect 44192 29124 44272 29152
rect 43257 29087 43315 29093
rect 43257 29053 43269 29087
rect 43303 29053 43315 29087
rect 43990 29084 43996 29096
rect 43257 29047 43315 29053
rect 43364 29056 43996 29084
rect 30374 29016 30380 29028
rect 22066 28988 30380 29016
rect 30374 28976 30380 28988
rect 30432 28976 30438 29028
rect 42794 28976 42800 29028
rect 42852 29016 42858 29028
rect 43364 29016 43392 29056
rect 43990 29044 43996 29056
rect 44048 29044 44054 29096
rect 42852 28988 43392 29016
rect 44100 29016 44128 29115
rect 44192 29093 44220 29124
rect 44266 29112 44272 29124
rect 44324 29112 44330 29164
rect 45094 29112 45100 29164
rect 45152 29152 45158 29164
rect 45649 29155 45707 29161
rect 45649 29152 45661 29155
rect 45152 29124 45661 29152
rect 45152 29112 45158 29124
rect 45649 29121 45661 29124
rect 45695 29121 45707 29155
rect 46109 29155 46167 29161
rect 46109 29152 46121 29155
rect 45649 29115 45707 29121
rect 46032 29124 46121 29152
rect 46032 29096 46060 29124
rect 46109 29121 46121 29124
rect 46155 29121 46167 29155
rect 46109 29115 46167 29121
rect 46198 29112 46204 29164
rect 46256 29152 46262 29164
rect 46293 29155 46351 29161
rect 46293 29152 46305 29155
rect 46256 29124 46305 29152
rect 46256 29112 46262 29124
rect 46293 29121 46305 29124
rect 46339 29121 46351 29155
rect 46293 29115 46351 29121
rect 47486 29112 47492 29164
rect 47544 29152 47550 29164
rect 48225 29155 48283 29161
rect 48225 29152 48237 29155
rect 47544 29124 48237 29152
rect 47544 29112 47550 29124
rect 48225 29121 48237 29124
rect 48271 29121 48283 29155
rect 48225 29115 48283 29121
rect 48498 29112 48504 29164
rect 48556 29112 48562 29164
rect 44177 29087 44235 29093
rect 44177 29053 44189 29087
rect 44223 29053 44235 29087
rect 44358 29084 44364 29096
rect 44177 29047 44235 29053
rect 44284 29056 44364 29084
rect 44284 29016 44312 29056
rect 44358 29044 44364 29056
rect 44416 29084 44422 29096
rect 45741 29087 45799 29093
rect 45741 29084 45753 29087
rect 44416 29056 45753 29084
rect 44416 29044 44422 29056
rect 45741 29053 45753 29056
rect 45787 29084 45799 29087
rect 45830 29084 45836 29096
rect 45787 29056 45836 29084
rect 45787 29053 45799 29056
rect 45741 29047 45799 29053
rect 45830 29044 45836 29056
rect 45888 29044 45894 29096
rect 46014 29044 46020 29096
rect 46072 29044 46078 29096
rect 44100 28988 44312 29016
rect 44453 29019 44511 29025
rect 42852 28976 42858 28988
rect 44453 28985 44465 29019
rect 44499 29016 44511 29019
rect 44542 29016 44548 29028
rect 44499 28988 44548 29016
rect 44499 28985 44511 28988
rect 44453 28979 44511 28985
rect 44542 28976 44548 28988
rect 44600 28976 44606 29028
rect 11977 28951 12035 28957
rect 11977 28917 11989 28951
rect 12023 28948 12035 28951
rect 12250 28948 12256 28960
rect 12023 28920 12256 28948
rect 12023 28917 12035 28920
rect 11977 28911 12035 28917
rect 12250 28908 12256 28920
rect 12308 28908 12314 28960
rect 15473 28951 15531 28957
rect 15473 28917 15485 28951
rect 15519 28948 15531 28951
rect 15654 28948 15660 28960
rect 15519 28920 15660 28948
rect 15519 28917 15531 28920
rect 15473 28911 15531 28917
rect 15654 28908 15660 28920
rect 15712 28908 15718 28960
rect 15930 28908 15936 28960
rect 15988 28948 15994 28960
rect 16761 28951 16819 28957
rect 16761 28948 16773 28951
rect 15988 28920 16773 28948
rect 15988 28908 15994 28920
rect 16761 28917 16773 28920
rect 16807 28917 16819 28951
rect 16761 28911 16819 28917
rect 38378 28908 38384 28960
rect 38436 28948 38442 28960
rect 39485 28951 39543 28957
rect 39485 28948 39497 28951
rect 38436 28920 39497 28948
rect 38436 28908 38442 28920
rect 39485 28917 39497 28920
rect 39531 28917 39543 28951
rect 39485 28911 39543 28917
rect 40126 28908 40132 28960
rect 40184 28948 40190 28960
rect 40497 28951 40555 28957
rect 40497 28948 40509 28951
rect 40184 28920 40509 28948
rect 40184 28908 40190 28920
rect 40497 28917 40509 28920
rect 40543 28917 40555 28951
rect 40497 28911 40555 28917
rect 46474 28908 46480 28960
rect 46532 28908 46538 28960
rect 48314 28908 48320 28960
rect 48372 28908 48378 28960
rect 48593 28951 48651 28957
rect 48593 28917 48605 28951
rect 48639 28948 48651 28951
rect 49234 28948 49240 28960
rect 48639 28920 49240 28948
rect 48639 28917 48651 28920
rect 48593 28911 48651 28917
rect 49234 28908 49240 28920
rect 49292 28908 49298 28960
rect 1104 28858 78844 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 78844 28858
rect 1104 28784 78844 28806
rect 10689 28747 10747 28753
rect 10689 28713 10701 28747
rect 10735 28744 10747 28747
rect 10778 28744 10784 28756
rect 10735 28716 10784 28744
rect 10735 28713 10747 28716
rect 10689 28707 10747 28713
rect 10778 28704 10784 28716
rect 10836 28704 10842 28756
rect 10873 28747 10931 28753
rect 10873 28713 10885 28747
rect 10919 28713 10931 28747
rect 10873 28707 10931 28713
rect 934 28636 940 28688
rect 992 28676 998 28688
rect 1857 28679 1915 28685
rect 1857 28676 1869 28679
rect 992 28648 1869 28676
rect 992 28636 998 28648
rect 1857 28645 1869 28648
rect 1903 28645 1915 28679
rect 1857 28639 1915 28645
rect 10888 28608 10916 28707
rect 11238 28704 11244 28756
rect 11296 28744 11302 28756
rect 11701 28747 11759 28753
rect 11701 28744 11713 28747
rect 11296 28716 11713 28744
rect 11296 28704 11302 28716
rect 11701 28713 11713 28716
rect 11747 28713 11759 28747
rect 11701 28707 11759 28713
rect 14550 28704 14556 28756
rect 14608 28704 14614 28756
rect 15841 28747 15899 28753
rect 15841 28713 15853 28747
rect 15887 28744 15899 28747
rect 16117 28747 16175 28753
rect 16117 28744 16129 28747
rect 15887 28716 16129 28744
rect 15887 28713 15899 28716
rect 15841 28707 15899 28713
rect 16117 28713 16129 28716
rect 16163 28713 16175 28747
rect 20809 28747 20867 28753
rect 20809 28744 20821 28747
rect 16117 28707 16175 28713
rect 20732 28716 20821 28744
rect 11146 28636 11152 28688
rect 11204 28636 11210 28688
rect 13633 28679 13691 28685
rect 13633 28676 13645 28679
rect 12544 28648 13645 28676
rect 11422 28608 11428 28620
rect 10888 28580 11428 28608
rect 11422 28568 11428 28580
rect 11480 28568 11486 28620
rect 2041 28543 2099 28549
rect 2041 28509 2053 28543
rect 2087 28540 2099 28543
rect 2130 28540 2136 28552
rect 2087 28512 2136 28540
rect 2087 28509 2099 28512
rect 2041 28503 2099 28509
rect 2130 28500 2136 28512
rect 2188 28500 2194 28552
rect 9490 28500 9496 28552
rect 9548 28500 9554 28552
rect 12544 28549 12572 28648
rect 13633 28645 13645 28648
rect 13679 28676 13691 28679
rect 19334 28676 19340 28688
rect 13679 28648 15608 28676
rect 13679 28645 13691 28648
rect 13633 28639 13691 28645
rect 13262 28568 13268 28620
rect 13320 28568 13326 28620
rect 15194 28568 15200 28620
rect 15252 28608 15258 28620
rect 15580 28608 15608 28648
rect 15948 28648 19340 28676
rect 15948 28608 15976 28648
rect 19334 28636 19340 28648
rect 19392 28676 19398 28688
rect 20162 28676 20168 28688
rect 19392 28648 20168 28676
rect 19392 28636 19398 28648
rect 20162 28636 20168 28648
rect 20220 28636 20226 28688
rect 20438 28636 20444 28688
rect 20496 28636 20502 28688
rect 20622 28636 20628 28688
rect 20680 28636 20686 28688
rect 16666 28608 16672 28620
rect 15252 28580 15424 28608
rect 15580 28580 15976 28608
rect 16224 28580 16672 28608
rect 15252 28568 15258 28580
rect 11517 28543 11575 28549
rect 11517 28540 11529 28543
rect 10980 28512 11529 28540
rect 9508 28472 9536 28500
rect 10870 28481 10876 28484
rect 10857 28475 10876 28481
rect 9508 28444 10824 28472
rect 10137 28407 10195 28413
rect 10137 28373 10149 28407
rect 10183 28404 10195 28407
rect 10502 28404 10508 28416
rect 10183 28376 10508 28404
rect 10183 28373 10195 28376
rect 10137 28367 10195 28373
rect 10502 28364 10508 28376
rect 10560 28364 10566 28416
rect 10796 28404 10824 28444
rect 10857 28441 10869 28475
rect 10928 28472 10934 28484
rect 10980 28472 11008 28512
rect 11517 28509 11529 28512
rect 11563 28509 11575 28543
rect 11517 28503 11575 28509
rect 12529 28543 12587 28549
rect 12529 28509 12541 28543
rect 12575 28509 12587 28543
rect 12529 28503 12587 28509
rect 13354 28500 13360 28552
rect 13412 28540 13418 28552
rect 14369 28543 14427 28549
rect 14369 28540 14381 28543
rect 13412 28512 14381 28540
rect 13412 28500 13418 28512
rect 14369 28509 14381 28512
rect 14415 28509 14427 28543
rect 14369 28503 14427 28509
rect 14553 28543 14611 28549
rect 14553 28509 14565 28543
rect 14599 28540 14611 28543
rect 14642 28540 14648 28552
rect 14599 28512 14648 28540
rect 14599 28509 14611 28512
rect 14553 28503 14611 28509
rect 14642 28500 14648 28512
rect 14700 28500 14706 28552
rect 15286 28500 15292 28552
rect 15344 28500 15350 28552
rect 15396 28549 15424 28580
rect 15381 28543 15439 28549
rect 15381 28509 15393 28543
rect 15427 28509 15439 28543
rect 15381 28503 15439 28509
rect 15565 28543 15623 28549
rect 15565 28509 15577 28543
rect 15611 28540 15623 28543
rect 15746 28540 15752 28552
rect 15611 28512 15752 28540
rect 15611 28509 15623 28512
rect 15565 28503 15623 28509
rect 15746 28500 15752 28512
rect 15804 28540 15810 28552
rect 16224 28540 16252 28580
rect 16666 28568 16672 28580
rect 16724 28568 16730 28620
rect 20346 28568 20352 28620
rect 20404 28608 20410 28620
rect 20732 28608 20760 28716
rect 20809 28713 20821 28716
rect 20855 28713 20867 28747
rect 20809 28707 20867 28713
rect 38286 28704 38292 28756
rect 38344 28704 38350 28756
rect 39117 28747 39175 28753
rect 39117 28744 39129 28747
rect 38672 28716 39129 28744
rect 20404 28580 20760 28608
rect 20404 28568 20410 28580
rect 35986 28568 35992 28620
rect 36044 28608 36050 28620
rect 36357 28611 36415 28617
rect 36357 28608 36369 28611
rect 36044 28580 36369 28608
rect 36044 28568 36050 28580
rect 36357 28577 36369 28580
rect 36403 28577 36415 28611
rect 36357 28571 36415 28577
rect 15804 28512 16252 28540
rect 15804 28500 15810 28512
rect 17402 28500 17408 28552
rect 17460 28540 17466 28552
rect 17586 28540 17592 28552
rect 17460 28512 17592 28540
rect 17460 28500 17466 28512
rect 17586 28500 17592 28512
rect 17644 28500 17650 28552
rect 19978 28500 19984 28552
rect 20036 28540 20042 28552
rect 20165 28543 20223 28549
rect 20165 28540 20177 28543
rect 20036 28512 20177 28540
rect 20036 28500 20042 28512
rect 20165 28509 20177 28512
rect 20211 28540 20223 28543
rect 20211 28512 20668 28540
rect 20211 28509 20223 28512
rect 20165 28503 20223 28509
rect 10928 28444 11008 28472
rect 11057 28475 11115 28481
rect 10857 28435 10876 28441
rect 10870 28432 10876 28435
rect 10928 28432 10934 28444
rect 11057 28441 11069 28475
rect 11103 28472 11115 28475
rect 11330 28472 11336 28484
rect 11103 28444 11336 28472
rect 11103 28441 11115 28444
rect 11057 28435 11115 28441
rect 11072 28404 11100 28435
rect 11330 28432 11336 28444
rect 11388 28432 11394 28484
rect 15470 28432 15476 28484
rect 15528 28472 15534 28484
rect 15930 28481 15936 28484
rect 15657 28475 15715 28481
rect 15657 28472 15669 28475
rect 15528 28444 15669 28472
rect 15528 28432 15534 28444
rect 15657 28441 15669 28444
rect 15703 28441 15715 28475
rect 15657 28435 15715 28441
rect 15873 28475 15936 28481
rect 15873 28441 15885 28475
rect 15919 28441 15936 28475
rect 15873 28435 15936 28441
rect 15930 28432 15936 28435
rect 15988 28432 15994 28484
rect 16298 28432 16304 28484
rect 16356 28432 16362 28484
rect 16482 28432 16488 28484
rect 16540 28432 16546 28484
rect 20254 28432 20260 28484
rect 20312 28432 20318 28484
rect 20441 28475 20499 28481
rect 20441 28441 20453 28475
rect 20487 28472 20499 28475
rect 20530 28472 20536 28484
rect 20487 28444 20536 28472
rect 20487 28441 20499 28444
rect 20441 28435 20499 28441
rect 20530 28432 20536 28444
rect 20588 28432 20594 28484
rect 20640 28472 20668 28512
rect 36722 28500 36728 28552
rect 36780 28500 36786 28552
rect 38378 28500 38384 28552
rect 38436 28540 38442 28552
rect 38672 28549 38700 28716
rect 39117 28713 39129 28716
rect 39163 28744 39175 28747
rect 43438 28744 43444 28756
rect 39163 28716 43444 28744
rect 39163 28713 39175 28716
rect 39117 28707 39175 28713
rect 43438 28704 43444 28716
rect 43496 28704 43502 28756
rect 38746 28636 38752 28688
rect 38804 28636 38810 28688
rect 42705 28679 42763 28685
rect 42705 28645 42717 28679
rect 42751 28676 42763 28679
rect 42794 28676 42800 28688
rect 42751 28648 42800 28676
rect 42751 28645 42763 28648
rect 42705 28639 42763 28645
rect 42794 28636 42800 28648
rect 42852 28636 42858 28688
rect 46293 28679 46351 28685
rect 46293 28645 46305 28679
rect 46339 28645 46351 28679
rect 46293 28639 46351 28645
rect 38764 28608 38792 28636
rect 39853 28611 39911 28617
rect 39853 28608 39865 28611
rect 38764 28580 39865 28608
rect 39853 28577 39865 28580
rect 39899 28577 39911 28611
rect 39853 28571 39911 28577
rect 40126 28568 40132 28620
rect 40184 28568 40190 28620
rect 40862 28568 40868 28620
rect 40920 28608 40926 28620
rect 41877 28611 41935 28617
rect 41877 28608 41889 28611
rect 40920 28580 41889 28608
rect 40920 28568 40926 28580
rect 41877 28577 41889 28580
rect 41923 28577 41935 28611
rect 45462 28608 45468 28620
rect 41877 28571 41935 28577
rect 42444 28580 45468 28608
rect 38565 28543 38623 28549
rect 38565 28540 38577 28543
rect 38436 28512 38577 28540
rect 38436 28500 38442 28512
rect 38565 28509 38577 28512
rect 38611 28509 38623 28543
rect 38565 28503 38623 28509
rect 38657 28543 38715 28549
rect 38657 28509 38669 28543
rect 38703 28509 38715 28543
rect 38657 28503 38715 28509
rect 38749 28543 38807 28549
rect 38749 28509 38761 28543
rect 38795 28509 38807 28543
rect 38749 28503 38807 28509
rect 38933 28543 38991 28549
rect 38933 28509 38945 28543
rect 38979 28540 38991 28543
rect 39022 28540 39028 28552
rect 38979 28512 39028 28540
rect 38979 28509 38991 28512
rect 38933 28503 38991 28509
rect 20777 28475 20835 28481
rect 20777 28472 20789 28475
rect 20640 28444 20789 28472
rect 20777 28441 20789 28444
rect 20823 28441 20835 28475
rect 20777 28435 20835 28441
rect 20993 28475 21051 28481
rect 20993 28441 21005 28475
rect 21039 28441 21051 28475
rect 20993 28435 21051 28441
rect 10796 28376 11100 28404
rect 11422 28364 11428 28416
rect 11480 28364 11486 28416
rect 14737 28407 14795 28413
rect 14737 28373 14749 28407
rect 14783 28404 14795 28407
rect 15102 28404 15108 28416
rect 14783 28376 15108 28404
rect 14783 28373 14795 28376
rect 14737 28367 14795 28373
rect 15102 28364 15108 28376
rect 15160 28364 15166 28416
rect 16022 28364 16028 28416
rect 16080 28364 16086 28416
rect 16114 28364 16120 28416
rect 16172 28404 16178 28416
rect 16761 28407 16819 28413
rect 16761 28404 16773 28407
rect 16172 28376 16773 28404
rect 16172 28364 16178 28376
rect 16761 28373 16773 28376
rect 16807 28373 16819 28407
rect 16761 28367 16819 28373
rect 19978 28364 19984 28416
rect 20036 28404 20042 28416
rect 20272 28404 20300 28432
rect 21008 28404 21036 28435
rect 37090 28432 37096 28484
rect 37148 28432 37154 28484
rect 20036 28376 21036 28404
rect 20036 28364 20042 28376
rect 37918 28364 37924 28416
rect 37976 28404 37982 28416
rect 38151 28407 38209 28413
rect 38151 28404 38163 28407
rect 37976 28376 38163 28404
rect 37976 28364 37982 28376
rect 38151 28373 38163 28376
rect 38197 28373 38209 28407
rect 38764 28404 38792 28503
rect 39022 28500 39028 28512
rect 39080 28500 39086 28552
rect 42444 28549 42472 28580
rect 45462 28568 45468 28580
rect 45520 28568 45526 28620
rect 42429 28543 42487 28549
rect 42429 28509 42441 28543
rect 42475 28509 42487 28543
rect 42429 28503 42487 28509
rect 42797 28543 42855 28549
rect 42797 28509 42809 28543
rect 42843 28509 42855 28543
rect 42797 28503 42855 28509
rect 42889 28543 42947 28549
rect 42889 28509 42901 28543
rect 42935 28540 42947 28543
rect 43349 28543 43407 28549
rect 43349 28540 43361 28543
rect 42935 28512 43361 28540
rect 42935 28509 42947 28512
rect 42889 28503 42947 28509
rect 43349 28509 43361 28512
rect 43395 28509 43407 28543
rect 43349 28503 43407 28509
rect 43441 28543 43499 28549
rect 43441 28509 43453 28543
rect 43487 28540 43499 28543
rect 43530 28540 43536 28552
rect 43487 28512 43536 28540
rect 43487 28509 43499 28512
rect 43441 28503 43499 28509
rect 42812 28472 42840 28503
rect 43530 28500 43536 28512
rect 43588 28540 43594 28552
rect 45094 28540 45100 28552
rect 43588 28512 45100 28540
rect 43588 28500 43594 28512
rect 45094 28500 45100 28512
rect 45152 28500 45158 28552
rect 46014 28500 46020 28552
rect 46072 28500 46078 28552
rect 46308 28540 46336 28639
rect 46566 28636 46572 28688
rect 46624 28676 46630 28688
rect 46661 28679 46719 28685
rect 46661 28676 46673 28679
rect 46624 28648 46673 28676
rect 46624 28636 46630 28648
rect 46661 28645 46673 28648
rect 46707 28645 46719 28679
rect 46661 28639 46719 28645
rect 47486 28568 47492 28620
rect 47544 28568 47550 28620
rect 49234 28568 49240 28620
rect 49292 28568 49298 28620
rect 46385 28543 46443 28549
rect 46385 28540 46397 28543
rect 46308 28512 46397 28540
rect 46385 28509 46397 28512
rect 46431 28509 46443 28543
rect 46385 28503 46443 28509
rect 46474 28500 46480 28552
rect 46532 28500 46538 28552
rect 49510 28500 49516 28552
rect 49568 28500 49574 28552
rect 40512 28444 40618 28472
rect 42812 28444 42932 28472
rect 40218 28404 40224 28416
rect 38764 28376 40224 28404
rect 38151 28367 38209 28373
rect 40218 28364 40224 28376
rect 40276 28404 40282 28416
rect 40512 28404 40540 28444
rect 42904 28416 42932 28444
rect 43990 28432 43996 28484
rect 44048 28472 44054 28484
rect 46109 28475 46167 28481
rect 46109 28472 46121 28475
rect 44048 28444 46121 28472
rect 44048 28432 44054 28444
rect 46109 28441 46121 28444
rect 46155 28472 46167 28475
rect 46198 28472 46204 28484
rect 46155 28444 46204 28472
rect 46155 28441 46167 28444
rect 46109 28435 46167 28441
rect 46198 28432 46204 28444
rect 46256 28432 46262 28484
rect 46293 28475 46351 28481
rect 46293 28441 46305 28475
rect 46339 28441 46351 28475
rect 46293 28435 46351 28441
rect 40276 28376 40540 28404
rect 40276 28364 40282 28376
rect 41414 28364 41420 28416
rect 41472 28404 41478 28416
rect 42521 28407 42579 28413
rect 42521 28404 42533 28407
rect 41472 28376 42533 28404
rect 41472 28364 41478 28376
rect 42521 28373 42533 28376
rect 42567 28373 42579 28407
rect 42521 28367 42579 28373
rect 42886 28364 42892 28416
rect 42944 28364 42950 28416
rect 43162 28364 43168 28416
rect 43220 28364 43226 28416
rect 45278 28364 45284 28416
rect 45336 28404 45342 28416
rect 45462 28404 45468 28416
rect 45336 28376 45468 28404
rect 45336 28364 45342 28376
rect 45462 28364 45468 28376
rect 45520 28404 45526 28416
rect 46308 28404 46336 28435
rect 46658 28432 46664 28484
rect 46716 28432 46722 28484
rect 48806 28444 49740 28472
rect 45520 28376 46336 28404
rect 45520 28364 45526 28376
rect 48222 28364 48228 28416
rect 48280 28404 48286 28416
rect 48884 28404 48912 28444
rect 49712 28413 49740 28444
rect 48280 28376 48912 28404
rect 49697 28407 49755 28413
rect 48280 28364 48286 28376
rect 49697 28373 49709 28407
rect 49743 28404 49755 28407
rect 55950 28404 55956 28416
rect 49743 28376 55956 28404
rect 49743 28373 49755 28376
rect 49697 28367 49755 28373
rect 55950 28364 55956 28376
rect 56008 28364 56014 28416
rect 1104 28314 78844 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 66314 28314
rect 66366 28262 66378 28314
rect 66430 28262 66442 28314
rect 66494 28262 66506 28314
rect 66558 28262 66570 28314
rect 66622 28262 78844 28314
rect 1104 28240 78844 28262
rect 8389 28203 8447 28209
rect 8389 28169 8401 28203
rect 8435 28200 8447 28203
rect 9490 28200 9496 28212
rect 8435 28172 9496 28200
rect 8435 28169 8447 28172
rect 8389 28163 8447 28169
rect 9490 28160 9496 28172
rect 9548 28160 9554 28212
rect 10686 28200 10692 28212
rect 9784 28172 10692 28200
rect 9784 28132 9812 28172
rect 10686 28160 10692 28172
rect 10744 28160 10750 28212
rect 14734 28200 14740 28212
rect 13280 28172 14740 28200
rect 13280 28144 13308 28172
rect 14734 28160 14740 28172
rect 14792 28160 14798 28212
rect 17954 28160 17960 28212
rect 18012 28200 18018 28212
rect 18417 28203 18475 28209
rect 18417 28200 18429 28203
rect 18012 28172 18429 28200
rect 18012 28160 18018 28172
rect 18417 28169 18429 28172
rect 18463 28169 18475 28203
rect 18417 28163 18475 28169
rect 20257 28203 20315 28209
rect 20257 28169 20269 28203
rect 20303 28200 20315 28203
rect 20346 28200 20352 28212
rect 20303 28172 20352 28200
rect 20303 28169 20315 28172
rect 20257 28163 20315 28169
rect 20346 28160 20352 28172
rect 20404 28160 20410 28212
rect 20530 28160 20536 28212
rect 20588 28200 20594 28212
rect 20625 28203 20683 28209
rect 20625 28200 20637 28203
rect 20588 28172 20637 28200
rect 20588 28160 20594 28172
rect 20625 28169 20637 28172
rect 20671 28169 20683 28203
rect 41969 28203 42027 28209
rect 20625 28163 20683 28169
rect 34900 28172 36308 28200
rect 9430 28104 9812 28132
rect 9861 28135 9919 28141
rect 9861 28101 9873 28135
rect 9907 28132 9919 28135
rect 10229 28135 10287 28141
rect 10229 28132 10241 28135
rect 9907 28104 10241 28132
rect 9907 28101 9919 28104
rect 9861 28095 9919 28101
rect 10229 28101 10241 28104
rect 10275 28101 10287 28135
rect 11057 28135 11115 28141
rect 11057 28132 11069 28135
rect 10229 28095 10287 28101
rect 10704 28104 11069 28132
rect 2041 28067 2099 28073
rect 2041 28033 2053 28067
rect 2087 28064 2099 28067
rect 2133 28067 2191 28073
rect 2133 28064 2145 28067
rect 2087 28036 2145 28064
rect 2087 28033 2099 28036
rect 2041 28027 2099 28033
rect 2133 28033 2145 28036
rect 2179 28033 2191 28067
rect 2133 28027 2191 28033
rect 10502 28024 10508 28076
rect 10560 28024 10566 28076
rect 10594 28024 10600 28076
rect 10652 28024 10658 28076
rect 10704 28073 10732 28104
rect 11057 28101 11069 28104
rect 11103 28101 11115 28135
rect 13262 28132 13268 28144
rect 11057 28095 11115 28101
rect 13096 28104 13268 28132
rect 10689 28067 10747 28073
rect 10689 28033 10701 28067
rect 10735 28033 10747 28067
rect 10689 28027 10747 28033
rect 10778 28024 10784 28076
rect 10836 28064 10842 28076
rect 10873 28067 10931 28073
rect 10873 28064 10885 28067
rect 10836 28036 10885 28064
rect 10836 28024 10842 28036
rect 10873 28033 10885 28036
rect 10919 28033 10931 28067
rect 10873 28027 10931 28033
rect 10962 28024 10968 28076
rect 11020 28024 11026 28076
rect 13096 28073 13124 28104
rect 13262 28092 13268 28104
rect 13320 28092 13326 28144
rect 14921 28135 14979 28141
rect 14921 28132 14933 28135
rect 14582 28104 14933 28132
rect 14921 28101 14933 28104
rect 14967 28132 14979 28135
rect 15010 28132 15016 28144
rect 14967 28104 15016 28132
rect 14967 28101 14979 28104
rect 14921 28095 14979 28101
rect 15010 28092 15016 28104
rect 15068 28092 15074 28144
rect 16022 28092 16028 28144
rect 16080 28132 16086 28144
rect 16945 28135 17003 28141
rect 16945 28132 16957 28135
rect 16080 28104 16957 28132
rect 16080 28092 16086 28104
rect 16945 28101 16957 28104
rect 16991 28101 17003 28135
rect 18598 28132 18604 28144
rect 18170 28104 18604 28132
rect 16945 28095 17003 28101
rect 18598 28092 18604 28104
rect 18656 28092 18662 28144
rect 19978 28092 19984 28144
rect 20036 28092 20042 28144
rect 20070 28092 20076 28144
rect 20128 28132 20134 28144
rect 20364 28132 20392 28160
rect 34900 28132 34928 28172
rect 36280 28132 36308 28172
rect 41969 28169 41981 28203
rect 42015 28200 42027 28203
rect 42794 28200 42800 28212
rect 42015 28172 42800 28200
rect 42015 28169 42027 28172
rect 41969 28163 42027 28169
rect 42794 28160 42800 28172
rect 42852 28160 42858 28212
rect 45833 28203 45891 28209
rect 45833 28169 45845 28203
rect 45879 28200 45891 28203
rect 45922 28200 45928 28212
rect 45879 28172 45928 28200
rect 45879 28169 45891 28172
rect 45833 28163 45891 28169
rect 45922 28160 45928 28172
rect 45980 28160 45986 28212
rect 47486 28200 47492 28212
rect 46032 28172 47492 28200
rect 37090 28132 37096 28144
rect 20128 28104 20300 28132
rect 20364 28104 21220 28132
rect 34270 28104 34928 28132
rect 36202 28104 37096 28132
rect 20128 28092 20134 28104
rect 13081 28067 13139 28073
rect 13081 28033 13093 28067
rect 13127 28033 13139 28067
rect 13081 28027 13139 28033
rect 15470 28024 15476 28076
rect 15528 28024 15534 28076
rect 15654 28024 15660 28076
rect 15712 28024 15718 28076
rect 15746 28024 15752 28076
rect 15804 28024 15810 28076
rect 15841 28067 15899 28073
rect 15841 28033 15853 28067
rect 15887 28064 15899 28067
rect 16114 28064 16120 28076
rect 15887 28036 16120 28064
rect 15887 28033 15899 28036
rect 15841 28027 15899 28033
rect 16114 28024 16120 28036
rect 16172 28024 16178 28076
rect 20162 28024 20168 28076
rect 20220 28024 20226 28076
rect 20272 28064 20300 28104
rect 21192 28073 21220 28104
rect 37090 28092 37096 28104
rect 37148 28092 37154 28144
rect 42886 28092 42892 28144
rect 42944 28132 42950 28144
rect 45462 28132 45468 28144
rect 42944 28104 45468 28132
rect 42944 28092 42950 28104
rect 20349 28067 20407 28073
rect 20349 28064 20361 28067
rect 20272 28036 20361 28064
rect 20349 28033 20361 28036
rect 20395 28033 20407 28067
rect 20349 28027 20407 28033
rect 21177 28067 21235 28073
rect 21177 28033 21189 28067
rect 21223 28033 21235 28067
rect 21177 28027 21235 28033
rect 32876 28036 33364 28064
rect 10137 27999 10195 28005
rect 10137 27965 10149 27999
rect 10183 27996 10195 27999
rect 10226 27996 10232 28008
rect 10183 27968 10232 27996
rect 10183 27965 10195 27968
rect 10137 27959 10195 27965
rect 10226 27956 10232 27968
rect 10284 27956 10290 28008
rect 13354 27956 13360 28008
rect 13412 27956 13418 28008
rect 14734 27956 14740 28008
rect 14792 27996 14798 28008
rect 16669 27999 16727 28005
rect 16669 27996 16681 27999
rect 14792 27968 16681 27996
rect 14792 27956 14798 27968
rect 16669 27965 16681 27968
rect 16715 27965 16727 27999
rect 16669 27959 16727 27965
rect 32030 27956 32036 28008
rect 32088 27996 32094 28008
rect 32876 28005 32904 28036
rect 32861 27999 32919 28005
rect 32861 27996 32873 27999
rect 32088 27968 32873 27996
rect 32088 27956 32094 27968
rect 32861 27965 32873 27968
rect 32907 27965 32919 27999
rect 32861 27959 32919 27965
rect 33226 27956 33232 28008
rect 33284 27956 33290 28008
rect 33336 27996 33364 28036
rect 40862 28024 40868 28076
rect 40920 28064 40926 28076
rect 41141 28067 41199 28073
rect 41141 28064 41153 28067
rect 40920 28036 41153 28064
rect 40920 28024 40926 28036
rect 41141 28033 41153 28036
rect 41187 28064 41199 28067
rect 42794 28064 42800 28076
rect 41187 28036 42800 28064
rect 41187 28033 41199 28036
rect 41141 28027 41199 28033
rect 42794 28024 42800 28036
rect 42852 28024 42858 28076
rect 34793 27999 34851 28005
rect 34793 27996 34805 27999
rect 33336 27968 34805 27996
rect 34793 27965 34805 27968
rect 34839 27965 34851 27999
rect 34793 27959 34851 27965
rect 35161 27999 35219 28005
rect 35161 27965 35173 27999
rect 35207 27996 35219 27999
rect 35342 27996 35348 28008
rect 35207 27968 35348 27996
rect 35207 27965 35219 27968
rect 35161 27959 35219 27965
rect 35342 27956 35348 27968
rect 35400 27956 35406 28008
rect 41230 27956 41236 28008
rect 41288 27956 41294 28008
rect 42978 27956 42984 28008
rect 43036 27996 43042 28008
rect 43180 28005 43208 28104
rect 45462 28092 45468 28104
rect 45520 28132 45526 28144
rect 46032 28132 46060 28172
rect 47486 28160 47492 28172
rect 47544 28160 47550 28212
rect 48317 28203 48375 28209
rect 48317 28169 48329 28203
rect 48363 28200 48375 28203
rect 48498 28200 48504 28212
rect 48363 28172 48504 28200
rect 48363 28169 48375 28172
rect 48317 28163 48375 28169
rect 48498 28160 48504 28172
rect 48556 28160 48562 28212
rect 45520 28104 46060 28132
rect 46385 28135 46443 28141
rect 45520 28092 45526 28104
rect 46385 28101 46397 28135
rect 46431 28132 46443 28135
rect 46658 28132 46664 28144
rect 46431 28104 46664 28132
rect 46431 28101 46443 28104
rect 46385 28095 46443 28101
rect 46658 28092 46664 28104
rect 46716 28092 46722 28144
rect 43257 28067 43315 28073
rect 43257 28033 43269 28067
rect 43303 28064 43315 28067
rect 43530 28064 43536 28076
rect 43303 28036 43536 28064
rect 43303 28033 43315 28036
rect 43257 28027 43315 28033
rect 43530 28024 43536 28036
rect 43588 28024 43594 28076
rect 43714 28024 43720 28076
rect 43772 28064 43778 28076
rect 44085 28067 44143 28073
rect 44085 28064 44097 28067
rect 43772 28036 44097 28064
rect 43772 28024 43778 28036
rect 44085 28033 44097 28036
rect 44131 28033 44143 28067
rect 44085 28027 44143 28033
rect 44174 28024 44180 28076
rect 44232 28064 44238 28076
rect 44232 28036 44277 28064
rect 44232 28024 44238 28036
rect 44726 28024 44732 28076
rect 44784 28064 44790 28076
rect 45094 28064 45100 28076
rect 44784 28036 45100 28064
rect 44784 28024 44790 28036
rect 45094 28024 45100 28036
rect 45152 28064 45158 28076
rect 45925 28067 45983 28073
rect 45925 28064 45937 28067
rect 45152 28036 45937 28064
rect 45152 28024 45158 28036
rect 45925 28033 45937 28036
rect 45971 28033 45983 28067
rect 45925 28027 45983 28033
rect 46566 28024 46572 28076
rect 46624 28064 46630 28076
rect 47857 28067 47915 28073
rect 47857 28064 47869 28067
rect 46624 28036 47869 28064
rect 46624 28024 46630 28036
rect 47857 28033 47869 28036
rect 47903 28033 47915 28067
rect 47857 28027 47915 28033
rect 47949 28067 48007 28073
rect 47949 28033 47961 28067
rect 47995 28064 48007 28067
rect 48314 28064 48320 28076
rect 47995 28036 48320 28064
rect 47995 28033 48007 28036
rect 47949 28027 48007 28033
rect 48314 28024 48320 28036
rect 48372 28024 48378 28076
rect 43073 27999 43131 28005
rect 43073 27996 43085 27999
rect 43036 27968 43085 27996
rect 43036 27956 43042 27968
rect 43073 27965 43085 27968
rect 43119 27965 43131 27999
rect 43073 27959 43131 27965
rect 43165 27999 43223 28005
rect 43165 27965 43177 27999
rect 43211 27965 43223 27999
rect 43165 27959 43223 27965
rect 44453 27999 44511 28005
rect 44453 27965 44465 27999
rect 44499 27996 44511 27999
rect 46106 27996 46112 28008
rect 44499 27968 46112 27996
rect 44499 27965 44511 27968
rect 44453 27959 44511 27965
rect 934 27888 940 27940
rect 992 27928 998 27940
rect 1857 27931 1915 27937
rect 1857 27928 1869 27931
rect 992 27900 1869 27928
rect 992 27888 998 27900
rect 1857 27897 1869 27900
rect 1903 27897 1915 27931
rect 1857 27891 1915 27897
rect 14642 27820 14648 27872
rect 14700 27860 14706 27872
rect 14829 27863 14887 27869
rect 14829 27860 14841 27863
rect 14700 27832 14841 27860
rect 14700 27820 14706 27832
rect 14829 27829 14841 27832
rect 14875 27829 14887 27863
rect 14829 27823 14887 27829
rect 16114 27820 16120 27872
rect 16172 27820 16178 27872
rect 18598 27820 18604 27872
rect 18656 27820 18662 27872
rect 19426 27820 19432 27872
rect 19484 27860 19490 27872
rect 20533 27863 20591 27869
rect 20533 27860 20545 27863
rect 19484 27832 20545 27860
rect 19484 27820 19490 27832
rect 20533 27829 20545 27832
rect 20579 27829 20591 27863
rect 20533 27823 20591 27829
rect 34514 27820 34520 27872
rect 34572 27860 34578 27872
rect 34655 27863 34713 27869
rect 34655 27860 34667 27863
rect 34572 27832 34667 27860
rect 34572 27820 34578 27832
rect 34655 27829 34667 27832
rect 34701 27829 34713 27863
rect 34655 27823 34713 27829
rect 36538 27820 36544 27872
rect 36596 27869 36602 27872
rect 36596 27863 36645 27869
rect 36596 27829 36599 27863
rect 36633 27829 36645 27863
rect 36596 27823 36645 27829
rect 36596 27820 36602 27823
rect 42978 27820 42984 27872
rect 43036 27860 43042 27872
rect 43180 27860 43208 27959
rect 46106 27956 46112 27968
rect 46164 27956 46170 28008
rect 47673 27999 47731 28005
rect 47673 27965 47685 27999
rect 47719 27965 47731 27999
rect 47673 27959 47731 27965
rect 44726 27888 44732 27940
rect 44784 27928 44790 27940
rect 45097 27931 45155 27937
rect 45097 27928 45109 27931
rect 44784 27900 45109 27928
rect 44784 27888 44790 27900
rect 45097 27897 45109 27900
rect 45143 27897 45155 27931
rect 45097 27891 45155 27897
rect 45649 27931 45707 27937
rect 45649 27897 45661 27931
rect 45695 27928 45707 27931
rect 46201 27931 46259 27937
rect 46201 27928 46213 27931
rect 45695 27900 46213 27928
rect 45695 27897 45707 27900
rect 45649 27891 45707 27897
rect 46201 27897 46213 27900
rect 46247 27897 46259 27931
rect 46201 27891 46259 27897
rect 47688 27872 47716 27959
rect 43036 27832 43208 27860
rect 43441 27863 43499 27869
rect 43036 27820 43042 27832
rect 43441 27829 43453 27863
rect 43487 27860 43499 27863
rect 43622 27860 43628 27872
rect 43487 27832 43628 27860
rect 43487 27829 43499 27832
rect 43441 27823 43499 27829
rect 43622 27820 43628 27832
rect 43680 27820 43686 27872
rect 45465 27863 45523 27869
rect 45465 27829 45477 27863
rect 45511 27860 45523 27863
rect 45830 27860 45836 27872
rect 45511 27832 45836 27860
rect 45511 27829 45523 27832
rect 45465 27823 45523 27829
rect 45830 27820 45836 27832
rect 45888 27820 45894 27872
rect 46014 27820 46020 27872
rect 46072 27820 46078 27872
rect 46106 27820 46112 27872
rect 46164 27820 46170 27872
rect 47397 27863 47455 27869
rect 47397 27829 47409 27863
rect 47443 27860 47455 27863
rect 47670 27860 47676 27872
rect 47443 27832 47676 27860
rect 47443 27829 47455 27832
rect 47397 27823 47455 27829
rect 47670 27820 47676 27832
rect 47728 27820 47734 27872
rect 1104 27770 78844 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 78844 27770
rect 1104 27696 78844 27718
rect 10594 27616 10600 27668
rect 10652 27656 10658 27668
rect 16114 27665 16120 27668
rect 10781 27659 10839 27665
rect 10781 27656 10793 27659
rect 10652 27628 10793 27656
rect 10652 27616 10658 27628
rect 10781 27625 10793 27628
rect 10827 27625 10839 27659
rect 10781 27619 10839 27625
rect 16104 27659 16120 27665
rect 16104 27625 16116 27659
rect 16104 27619 16120 27625
rect 16114 27616 16120 27619
rect 16172 27616 16178 27668
rect 17586 27616 17592 27668
rect 17644 27616 17650 27668
rect 33226 27616 33232 27668
rect 33284 27656 33290 27668
rect 33873 27659 33931 27665
rect 33873 27656 33885 27659
rect 33284 27628 33885 27656
rect 33284 27616 33290 27628
rect 33873 27625 33885 27628
rect 33919 27625 33931 27659
rect 33873 27619 33931 27625
rect 35161 27659 35219 27665
rect 35161 27625 35173 27659
rect 35207 27656 35219 27659
rect 35342 27656 35348 27668
rect 35207 27628 35348 27656
rect 35207 27625 35219 27628
rect 35161 27619 35219 27625
rect 35342 27616 35348 27628
rect 35400 27616 35406 27668
rect 36633 27659 36691 27665
rect 36633 27625 36645 27659
rect 36679 27656 36691 27659
rect 36722 27656 36728 27668
rect 36679 27628 36728 27656
rect 36679 27625 36691 27628
rect 36633 27619 36691 27625
rect 36722 27616 36728 27628
rect 36780 27616 36786 27668
rect 42702 27616 42708 27668
rect 42760 27656 42766 27668
rect 43073 27659 43131 27665
rect 42760 27628 43024 27656
rect 42760 27616 42766 27628
rect 12897 27591 12955 27597
rect 12897 27557 12909 27591
rect 12943 27588 12955 27591
rect 13354 27588 13360 27600
rect 12943 27560 13360 27588
rect 12943 27557 12955 27560
rect 12897 27551 12955 27557
rect 13354 27548 13360 27560
rect 13412 27548 13418 27600
rect 34422 27548 34428 27600
rect 34480 27588 34486 27600
rect 35621 27591 35679 27597
rect 35621 27588 35633 27591
rect 34480 27560 35633 27588
rect 34480 27548 34486 27560
rect 35621 27557 35633 27560
rect 35667 27557 35679 27591
rect 42886 27588 42892 27600
rect 35621 27551 35679 27557
rect 42628 27560 42892 27588
rect 12434 27480 12440 27532
rect 12492 27480 12498 27532
rect 14734 27480 14740 27532
rect 14792 27520 14798 27532
rect 15841 27523 15899 27529
rect 15841 27520 15853 27523
rect 14792 27492 15853 27520
rect 14792 27480 14798 27492
rect 15841 27489 15853 27492
rect 15887 27489 15899 27523
rect 15841 27483 15899 27489
rect 20162 27480 20168 27532
rect 20220 27520 20226 27532
rect 20533 27523 20591 27529
rect 20533 27520 20545 27523
rect 20220 27492 20545 27520
rect 20220 27480 20226 27492
rect 20533 27489 20545 27492
rect 20579 27489 20591 27523
rect 20533 27483 20591 27489
rect 31662 27480 31668 27532
rect 31720 27520 31726 27532
rect 34333 27523 34391 27529
rect 34333 27520 34345 27523
rect 31720 27492 34345 27520
rect 31720 27480 31726 27492
rect 34333 27489 34345 27492
rect 34379 27489 34391 27523
rect 34333 27483 34391 27489
rect 37093 27523 37151 27529
rect 37093 27489 37105 27523
rect 37139 27489 37151 27523
rect 37093 27483 37151 27489
rect 2041 27455 2099 27461
rect 2041 27421 2053 27455
rect 2087 27452 2099 27455
rect 2133 27455 2191 27461
rect 2133 27452 2145 27455
rect 2087 27424 2145 27452
rect 2087 27421 2099 27424
rect 2041 27415 2099 27421
rect 2133 27421 2145 27424
rect 2179 27421 2191 27455
rect 2133 27415 2191 27421
rect 10962 27412 10968 27464
rect 11020 27412 11026 27464
rect 11149 27455 11207 27461
rect 11149 27421 11161 27455
rect 11195 27452 11207 27455
rect 11330 27452 11336 27464
rect 11195 27424 11336 27452
rect 11195 27421 11207 27424
rect 11149 27415 11207 27421
rect 11330 27412 11336 27424
rect 11388 27412 11394 27464
rect 12529 27455 12587 27461
rect 12529 27421 12541 27455
rect 12575 27452 12587 27455
rect 14093 27455 14151 27461
rect 14093 27452 14105 27455
rect 12575 27424 14105 27452
rect 12575 27421 12587 27424
rect 12529 27415 12587 27421
rect 14093 27421 14105 27424
rect 14139 27421 14151 27455
rect 14093 27415 14151 27421
rect 14642 27412 14648 27464
rect 14700 27412 14706 27464
rect 19426 27412 19432 27464
rect 19484 27412 19490 27464
rect 19705 27455 19763 27461
rect 19705 27421 19717 27455
rect 19751 27421 19763 27455
rect 19705 27415 19763 27421
rect 19889 27455 19947 27461
rect 19889 27421 19901 27455
rect 19935 27452 19947 27455
rect 19981 27455 20039 27461
rect 19981 27452 19993 27455
rect 19935 27424 19993 27452
rect 19935 27421 19947 27424
rect 19889 27415 19947 27421
rect 19981 27421 19993 27424
rect 20027 27421 20039 27455
rect 19981 27415 20039 27421
rect 22465 27455 22523 27461
rect 22465 27421 22477 27455
rect 22511 27452 22523 27455
rect 23566 27452 23572 27464
rect 22511 27424 23572 27452
rect 22511 27421 22523 27424
rect 22465 27415 22523 27421
rect 15010 27344 15016 27396
rect 15068 27384 15074 27396
rect 19720 27384 19748 27415
rect 23566 27412 23572 27424
rect 23624 27412 23630 27464
rect 34054 27412 34060 27464
rect 34112 27412 34118 27464
rect 34146 27412 34152 27464
rect 34204 27412 34210 27464
rect 34425 27455 34483 27461
rect 34425 27421 34437 27455
rect 34471 27452 34483 27455
rect 34514 27452 34520 27464
rect 34471 27424 34520 27452
rect 34471 27421 34483 27424
rect 34425 27415 34483 27421
rect 34514 27412 34520 27424
rect 34572 27412 34578 27464
rect 35345 27455 35403 27461
rect 35345 27421 35357 27455
rect 35391 27421 35403 27455
rect 35345 27415 35403 27421
rect 20622 27384 20628 27396
rect 15068 27356 16606 27384
rect 19720 27356 20628 27384
rect 15068 27344 15074 27356
rect 934 27276 940 27328
rect 992 27316 998 27328
rect 1857 27319 1915 27325
rect 1857 27316 1869 27319
rect 992 27288 1869 27316
rect 992 27276 998 27288
rect 1857 27285 1869 27288
rect 1903 27285 1915 27319
rect 16546 27316 16574 27356
rect 20622 27344 20628 27356
rect 20680 27344 20686 27396
rect 21758 27356 21864 27384
rect 17681 27319 17739 27325
rect 17681 27316 17693 27319
rect 16546 27288 17693 27316
rect 1857 27279 1915 27285
rect 17681 27285 17693 27288
rect 17727 27316 17739 27319
rect 17954 27316 17960 27328
rect 17727 27288 17960 27316
rect 17727 27285 17739 27288
rect 17681 27279 17739 27285
rect 17954 27276 17960 27288
rect 18012 27276 18018 27328
rect 18506 27276 18512 27328
rect 18564 27316 18570 27328
rect 19245 27319 19303 27325
rect 19245 27316 19257 27319
rect 18564 27288 19257 27316
rect 18564 27276 18570 27288
rect 19245 27285 19257 27288
rect 19291 27285 19303 27319
rect 19245 27279 19303 27285
rect 20346 27276 20352 27328
rect 20404 27316 20410 27328
rect 20717 27319 20775 27325
rect 20717 27316 20729 27319
rect 20404 27288 20729 27316
rect 20404 27276 20410 27288
rect 20717 27285 20729 27288
rect 20763 27285 20775 27319
rect 21836 27316 21864 27356
rect 21910 27344 21916 27396
rect 21968 27384 21974 27396
rect 22189 27387 22247 27393
rect 22189 27384 22201 27387
rect 21968 27356 22201 27384
rect 21968 27344 21974 27356
rect 22189 27353 22201 27356
rect 22235 27353 22247 27387
rect 22189 27347 22247 27353
rect 32582 27344 32588 27396
rect 32640 27384 32646 27396
rect 35360 27384 35388 27415
rect 35434 27412 35440 27464
rect 35492 27412 35498 27464
rect 35713 27455 35771 27461
rect 35713 27421 35725 27455
rect 35759 27452 35771 27455
rect 36538 27452 36544 27464
rect 35759 27424 36544 27452
rect 35759 27421 35771 27424
rect 35713 27415 35771 27421
rect 36538 27412 36544 27424
rect 36596 27412 36602 27464
rect 36817 27455 36875 27461
rect 36817 27421 36829 27455
rect 36863 27421 36875 27455
rect 36817 27415 36875 27421
rect 36832 27384 36860 27415
rect 36906 27412 36912 27464
rect 36964 27412 36970 27464
rect 32640 27356 36860 27384
rect 32640 27344 32646 27356
rect 22649 27319 22707 27325
rect 22649 27316 22661 27319
rect 21836 27288 22661 27316
rect 20717 27279 20775 27285
rect 22649 27285 22661 27288
rect 22695 27316 22707 27319
rect 22830 27316 22836 27328
rect 22695 27288 22836 27316
rect 22695 27285 22707 27288
rect 22649 27279 22707 27285
rect 22830 27276 22836 27288
rect 22888 27276 22894 27328
rect 36354 27276 36360 27328
rect 36412 27316 36418 27328
rect 36449 27319 36507 27325
rect 36449 27316 36461 27319
rect 36412 27288 36461 27316
rect 36412 27276 36418 27288
rect 36449 27285 36461 27288
rect 36495 27316 36507 27319
rect 37108 27316 37136 27483
rect 37826 27480 37832 27532
rect 37884 27520 37890 27532
rect 38746 27520 38752 27532
rect 37884 27492 38752 27520
rect 37884 27480 37890 27492
rect 38746 27480 38752 27492
rect 38804 27480 38810 27532
rect 42628 27529 42656 27560
rect 42886 27548 42892 27560
rect 42944 27548 42950 27600
rect 42996 27588 43024 27628
rect 43073 27625 43085 27659
rect 43119 27656 43131 27659
rect 43530 27656 43536 27668
rect 43119 27628 43536 27656
rect 43119 27625 43131 27628
rect 43073 27619 43131 27625
rect 43530 27616 43536 27628
rect 43588 27616 43594 27668
rect 43993 27591 44051 27597
rect 43993 27588 44005 27591
rect 42996 27560 44005 27588
rect 43993 27557 44005 27560
rect 44039 27557 44051 27591
rect 43993 27551 44051 27557
rect 42613 27523 42671 27529
rect 42613 27489 42625 27523
rect 42659 27489 42671 27523
rect 44174 27520 44180 27532
rect 42613 27483 42671 27489
rect 42720 27492 44180 27520
rect 37185 27455 37243 27461
rect 37185 27421 37197 27455
rect 37231 27452 37243 27455
rect 37918 27452 37924 27464
rect 37231 27424 37924 27452
rect 37231 27421 37243 27424
rect 37185 27415 37243 27421
rect 37918 27412 37924 27424
rect 37976 27412 37982 27464
rect 38102 27412 38108 27464
rect 38160 27452 38166 27464
rect 42720 27461 42748 27492
rect 44174 27480 44180 27492
rect 44232 27480 44238 27532
rect 38197 27455 38255 27461
rect 38197 27452 38209 27455
rect 38160 27424 38209 27452
rect 38160 27412 38166 27424
rect 38197 27421 38209 27424
rect 38243 27421 38255 27455
rect 38197 27415 38255 27421
rect 42705 27455 42763 27461
rect 42705 27421 42717 27455
rect 42751 27421 42763 27455
rect 42705 27415 42763 27421
rect 39206 27344 39212 27396
rect 39264 27344 39270 27396
rect 41230 27344 41236 27396
rect 41288 27384 41294 27396
rect 42720 27384 42748 27415
rect 42978 27412 42984 27464
rect 43036 27452 43042 27464
rect 43073 27455 43131 27461
rect 43073 27452 43085 27455
rect 43036 27424 43085 27452
rect 43036 27412 43042 27424
rect 43073 27421 43085 27424
rect 43119 27421 43131 27455
rect 43073 27415 43131 27421
rect 43346 27412 43352 27464
rect 43404 27412 43410 27464
rect 43533 27455 43591 27461
rect 43533 27421 43545 27455
rect 43579 27421 43591 27455
rect 43533 27415 43591 27421
rect 43548 27384 43576 27415
rect 43622 27412 43628 27464
rect 43680 27412 43686 27464
rect 43714 27412 43720 27464
rect 43772 27452 43778 27464
rect 43772 27424 43817 27452
rect 43772 27412 43778 27424
rect 45830 27412 45836 27464
rect 45888 27412 45894 27464
rect 41288 27356 42748 27384
rect 43272 27356 43576 27384
rect 41288 27344 41294 27356
rect 43272 27328 43300 27356
rect 36495 27288 37136 27316
rect 36495 27285 36507 27288
rect 36449 27279 36507 27285
rect 38654 27276 38660 27328
rect 38712 27316 38718 27328
rect 39623 27319 39681 27325
rect 39623 27316 39635 27319
rect 38712 27288 39635 27316
rect 38712 27276 38718 27288
rect 39623 27285 39635 27288
rect 39669 27285 39681 27319
rect 39623 27279 39681 27285
rect 43254 27276 43260 27328
rect 43312 27276 43318 27328
rect 45922 27276 45928 27328
rect 45980 27276 45986 27328
rect 49326 27276 49332 27328
rect 49384 27316 49390 27328
rect 51258 27316 51264 27328
rect 49384 27288 51264 27316
rect 49384 27276 49390 27288
rect 51258 27276 51264 27288
rect 51316 27276 51322 27328
rect 1104 27226 78844 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 66314 27226
rect 66366 27174 66378 27226
rect 66430 27174 66442 27226
rect 66494 27174 66506 27226
rect 66558 27174 66570 27226
rect 66622 27174 78844 27226
rect 1104 27152 78844 27174
rect 10305 27115 10363 27121
rect 10305 27081 10317 27115
rect 10351 27112 10363 27115
rect 10689 27115 10747 27121
rect 10689 27112 10701 27115
rect 10351 27084 10701 27112
rect 10351 27081 10363 27084
rect 10305 27075 10363 27081
rect 10689 27081 10701 27084
rect 10735 27081 10747 27115
rect 10689 27075 10747 27081
rect 10778 27072 10784 27124
rect 10836 27072 10842 27124
rect 12066 27072 12072 27124
rect 12124 27112 12130 27124
rect 12124 27084 12572 27112
rect 12124 27072 12130 27084
rect 10042 27004 10048 27056
rect 10100 27044 10106 27056
rect 10505 27047 10563 27053
rect 10505 27044 10517 27047
rect 10100 27016 10517 27044
rect 10100 27004 10106 27016
rect 10505 27013 10517 27016
rect 10551 27044 10563 27047
rect 10796 27044 10824 27072
rect 10551 27016 12296 27044
rect 10551 27013 10563 27016
rect 10505 27007 10563 27013
rect 10594 26936 10600 26988
rect 10652 26976 10658 26988
rect 10781 26979 10839 26985
rect 10781 26976 10793 26979
rect 10652 26948 10793 26976
rect 10652 26936 10658 26948
rect 10781 26945 10793 26948
rect 10827 26945 10839 26979
rect 10781 26939 10839 26945
rect 11330 26936 11336 26988
rect 11388 26976 11394 26988
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11388 26948 11713 26976
rect 11388 26936 11394 26948
rect 11701 26945 11713 26948
rect 11747 26976 11759 26979
rect 12066 26976 12072 26988
rect 11747 26948 12072 26976
rect 11747 26945 11759 26948
rect 11701 26939 11759 26945
rect 12066 26936 12072 26948
rect 12124 26936 12130 26988
rect 12268 26985 12296 27016
rect 12253 26979 12311 26985
rect 12253 26945 12265 26979
rect 12299 26945 12311 26979
rect 12253 26939 12311 26945
rect 12434 26936 12440 26988
rect 12492 26936 12498 26988
rect 12544 26985 12572 27084
rect 18138 27072 18144 27124
rect 18196 27112 18202 27124
rect 18598 27112 18604 27124
rect 18196 27084 18604 27112
rect 18196 27072 18202 27084
rect 18598 27072 18604 27084
rect 18656 27072 18662 27124
rect 19981 27115 20039 27121
rect 19981 27081 19993 27115
rect 20027 27112 20039 27115
rect 20162 27112 20168 27124
rect 20027 27084 20168 27112
rect 20027 27081 20039 27084
rect 19981 27075 20039 27081
rect 20162 27072 20168 27084
rect 20220 27072 20226 27124
rect 20533 27115 20591 27121
rect 20533 27081 20545 27115
rect 20579 27112 20591 27115
rect 21910 27112 21916 27124
rect 20579 27084 21916 27112
rect 20579 27081 20591 27084
rect 20533 27075 20591 27081
rect 21910 27072 21916 27084
rect 21968 27072 21974 27124
rect 31386 27072 31392 27124
rect 31444 27112 31450 27124
rect 31941 27115 31999 27121
rect 31941 27112 31953 27115
rect 31444 27084 31953 27112
rect 31444 27072 31450 27084
rect 31941 27081 31953 27084
rect 31987 27112 31999 27115
rect 35253 27115 35311 27121
rect 31987 27084 32812 27112
rect 31987 27081 31999 27084
rect 31941 27075 31999 27081
rect 18506 27004 18512 27056
rect 18564 27004 18570 27056
rect 18616 27044 18644 27072
rect 32784 27044 32812 27084
rect 35253 27081 35265 27115
rect 35299 27112 35311 27115
rect 35434 27112 35440 27124
rect 35299 27084 35440 27112
rect 35299 27081 35311 27084
rect 35253 27075 35311 27081
rect 35434 27072 35440 27084
rect 35492 27072 35498 27124
rect 36722 27112 36728 27124
rect 35728 27084 36728 27112
rect 18616 27016 18998 27044
rect 32784 27016 32890 27044
rect 34514 27004 34520 27056
rect 34572 27044 34578 27056
rect 34572 27016 35572 27044
rect 34572 27004 34578 27016
rect 35544 26988 35572 27016
rect 12529 26979 12587 26985
rect 12529 26945 12541 26979
rect 12575 26945 12587 26979
rect 12529 26939 12587 26945
rect 12621 26979 12679 26985
rect 12621 26945 12633 26979
rect 12667 26976 12679 26979
rect 12986 26976 12992 26988
rect 12667 26948 12992 26976
rect 12667 26945 12679 26948
rect 12621 26939 12679 26945
rect 12986 26936 12992 26948
rect 13044 26936 13050 26988
rect 13354 26936 13360 26988
rect 13412 26936 13418 26988
rect 14734 26936 14740 26988
rect 14792 26936 14798 26988
rect 20438 26936 20444 26988
rect 20496 26936 20502 26988
rect 20622 26936 20628 26988
rect 20680 26936 20686 26988
rect 35437 26979 35495 26985
rect 35437 26976 35449 26979
rect 35084 26948 35449 26976
rect 2038 26868 2044 26920
rect 2096 26868 2102 26920
rect 11793 26911 11851 26917
rect 11793 26877 11805 26911
rect 11839 26877 11851 26911
rect 11793 26871 11851 26877
rect 11885 26911 11943 26917
rect 11885 26877 11897 26911
rect 11931 26877 11943 26911
rect 11885 26871 11943 26877
rect 11977 26911 12035 26917
rect 11977 26877 11989 26911
rect 12023 26908 12035 26911
rect 12897 26911 12955 26917
rect 12023 26880 12434 26908
rect 12023 26877 12035 26880
rect 11977 26871 12035 26877
rect 11517 26843 11575 26849
rect 11517 26840 11529 26843
rect 10336 26812 11529 26840
rect 10134 26732 10140 26784
rect 10192 26732 10198 26784
rect 10336 26781 10364 26812
rect 11517 26809 11529 26812
rect 11563 26809 11575 26843
rect 11517 26803 11575 26809
rect 10321 26775 10379 26781
rect 10321 26741 10333 26775
rect 10367 26741 10379 26775
rect 11808 26772 11836 26871
rect 11900 26840 11928 26871
rect 12158 26840 12164 26852
rect 11900 26812 12164 26840
rect 12158 26800 12164 26812
rect 12216 26800 12222 26852
rect 12406 26840 12434 26880
rect 12897 26877 12909 26911
rect 12943 26908 12955 26911
rect 14461 26911 14519 26917
rect 14461 26908 14473 26911
rect 12943 26880 14473 26908
rect 12943 26877 12955 26880
rect 12897 26871 12955 26877
rect 14461 26877 14473 26880
rect 14507 26877 14519 26911
rect 14461 26871 14519 26877
rect 18230 26868 18236 26920
rect 18288 26868 18294 26920
rect 32030 26868 32036 26920
rect 32088 26908 32094 26920
rect 32125 26911 32183 26917
rect 32125 26908 32137 26911
rect 32088 26880 32137 26908
rect 32088 26868 32094 26880
rect 32125 26877 32137 26880
rect 32171 26877 32183 26911
rect 32125 26871 32183 26877
rect 32490 26868 32496 26920
rect 32548 26868 32554 26920
rect 12526 26840 12532 26852
rect 12406 26812 12532 26840
rect 12526 26800 12532 26812
rect 12584 26800 12590 26852
rect 12912 26812 13492 26840
rect 11974 26772 11980 26784
rect 11808 26744 11980 26772
rect 10321 26735 10379 26741
rect 11974 26732 11980 26744
rect 12032 26772 12038 26784
rect 12912 26772 12940 26812
rect 12032 26744 12940 26772
rect 12032 26732 12038 26744
rect 12986 26732 12992 26784
rect 13044 26732 13050 26784
rect 13464 26772 13492 26812
rect 14642 26772 14648 26784
rect 13464 26744 14648 26772
rect 14642 26732 14648 26744
rect 14700 26732 14706 26784
rect 18138 26732 18144 26784
rect 18196 26732 18202 26784
rect 33962 26781 33968 26784
rect 33919 26775 33968 26781
rect 33919 26741 33931 26775
rect 33965 26741 33968 26775
rect 33919 26735 33968 26741
rect 33962 26732 33968 26735
rect 34020 26732 34026 26784
rect 34606 26732 34612 26784
rect 34664 26772 34670 26784
rect 35084 26781 35112 26948
rect 35437 26945 35449 26948
rect 35483 26945 35495 26979
rect 35437 26939 35495 26945
rect 35452 26908 35480 26939
rect 35526 26936 35532 26988
rect 35584 26936 35590 26988
rect 35618 26936 35624 26988
rect 35676 26936 35682 26988
rect 35728 26908 35756 27084
rect 36722 27072 36728 27084
rect 36780 27072 36786 27124
rect 36906 27072 36912 27124
rect 36964 27072 36970 27124
rect 38102 27072 38108 27124
rect 38160 27072 38166 27124
rect 43714 27112 43720 27124
rect 42904 27084 43720 27112
rect 36265 27047 36323 27053
rect 36265 27013 36277 27047
rect 36311 27044 36323 27047
rect 36541 27047 36599 27053
rect 36541 27044 36553 27047
rect 36311 27016 36553 27044
rect 36311 27013 36323 27016
rect 36265 27007 36323 27013
rect 36541 27013 36553 27016
rect 36587 27044 36599 27047
rect 36998 27044 37004 27056
rect 36587 27016 37004 27044
rect 36587 27013 36599 27016
rect 36541 27007 36599 27013
rect 36998 27004 37004 27016
rect 37056 27004 37062 27056
rect 39206 27004 39212 27056
rect 39264 27044 39270 27056
rect 39264 27016 40434 27044
rect 39264 27004 39270 27016
rect 35805 26979 35863 26985
rect 35805 26945 35817 26979
rect 35851 26976 35863 26979
rect 36357 26979 36415 26985
rect 35851 26948 36308 26976
rect 35851 26945 35863 26948
rect 35805 26939 35863 26945
rect 35989 26911 36047 26917
rect 35989 26908 36001 26911
rect 35452 26880 36001 26908
rect 35989 26877 36001 26880
rect 36035 26877 36047 26911
rect 35989 26871 36047 26877
rect 35069 26775 35127 26781
rect 35069 26772 35081 26775
rect 34664 26744 35081 26772
rect 34664 26732 34670 26744
rect 35069 26741 35081 26744
rect 35115 26741 35127 26775
rect 36280 26772 36308 26948
rect 36357 26945 36369 26979
rect 36403 26945 36415 26979
rect 36357 26939 36415 26945
rect 36633 26979 36691 26985
rect 36633 26945 36645 26979
rect 36679 26945 36691 26979
rect 36633 26939 36691 26945
rect 36372 26840 36400 26939
rect 36538 26868 36544 26920
rect 36596 26908 36602 26920
rect 36648 26908 36676 26939
rect 36722 26936 36728 26988
rect 36780 26976 36786 26988
rect 37274 26976 37280 26988
rect 36780 26948 37280 26976
rect 36780 26936 36786 26948
rect 37274 26936 37280 26948
rect 37332 26936 37338 26988
rect 37366 26936 37372 26988
rect 37424 26976 37430 26988
rect 38289 26979 38347 26985
rect 38289 26976 38301 26979
rect 37424 26948 38301 26976
rect 37424 26936 37430 26948
rect 38289 26945 38301 26948
rect 38335 26945 38347 26979
rect 38289 26939 38347 26945
rect 38378 26936 38384 26988
rect 38436 26936 38442 26988
rect 38654 26936 38660 26988
rect 38712 26936 38718 26988
rect 38746 26936 38752 26988
rect 38804 26976 38810 26988
rect 39669 26979 39727 26985
rect 39669 26976 39681 26979
rect 38804 26948 39681 26976
rect 38804 26936 38810 26948
rect 39669 26945 39681 26948
rect 39715 26945 39727 26979
rect 39669 26939 39727 26945
rect 42429 26979 42487 26985
rect 42429 26945 42441 26979
rect 42475 26976 42487 26979
rect 42794 26976 42800 26988
rect 42475 26948 42800 26976
rect 42475 26945 42487 26948
rect 42429 26939 42487 26945
rect 42794 26936 42800 26948
rect 42852 26976 42858 26988
rect 42904 26985 42932 27084
rect 43714 27072 43720 27084
rect 43772 27072 43778 27124
rect 46014 27072 46020 27124
rect 46072 27072 46078 27124
rect 48406 27072 48412 27124
rect 48464 27112 48470 27124
rect 48464 27084 50108 27112
rect 48464 27072 48470 27084
rect 42981 27047 43039 27053
rect 42981 27013 42993 27047
rect 43027 27044 43039 27047
rect 46032 27044 46060 27072
rect 50080 27044 50108 27084
rect 53926 27044 53932 27056
rect 43027 27016 43668 27044
rect 43027 27013 43039 27016
rect 42981 27007 43039 27013
rect 42889 26979 42947 26985
rect 42889 26976 42901 26979
rect 42852 26948 42901 26976
rect 42852 26936 42858 26948
rect 42889 26945 42901 26948
rect 42935 26945 42947 26979
rect 42889 26939 42947 26945
rect 43073 26979 43131 26985
rect 43073 26945 43085 26979
rect 43119 26976 43131 26979
rect 43530 26976 43536 26988
rect 43119 26948 43536 26976
rect 43119 26945 43131 26948
rect 43073 26939 43131 26945
rect 43530 26936 43536 26948
rect 43588 26936 43594 26988
rect 43640 26985 43668 27016
rect 44100 27016 46060 27044
rect 50002 27016 51106 27044
rect 53774 27016 53932 27044
rect 43625 26979 43683 26985
rect 43625 26945 43637 26979
rect 43671 26945 43683 26979
rect 43625 26939 43683 26945
rect 38672 26908 38700 26936
rect 36596 26880 36676 26908
rect 37200 26880 38700 26908
rect 39945 26911 40003 26917
rect 36596 26868 36602 26880
rect 37200 26852 37228 26880
rect 39945 26877 39957 26911
rect 39991 26908 40003 26911
rect 40402 26908 40408 26920
rect 39991 26880 40408 26908
rect 39991 26877 40003 26880
rect 39945 26871 40003 26877
rect 40402 26868 40408 26880
rect 40460 26868 40466 26920
rect 41230 26868 41236 26920
rect 41288 26908 41294 26920
rect 41693 26911 41751 26917
rect 41693 26908 41705 26911
rect 41288 26880 41705 26908
rect 41288 26868 41294 26880
rect 41693 26877 41705 26880
rect 41739 26877 41751 26911
rect 41693 26871 41751 26877
rect 42705 26911 42763 26917
rect 42705 26877 42717 26911
rect 42751 26908 42763 26911
rect 43254 26908 43260 26920
rect 42751 26880 43260 26908
rect 42751 26877 42763 26880
rect 42705 26871 42763 26877
rect 43254 26868 43260 26880
rect 43312 26868 43318 26920
rect 43346 26868 43352 26920
rect 43404 26908 43410 26920
rect 44100 26908 44128 27016
rect 53926 27004 53932 27016
rect 53984 27004 53990 27056
rect 44177 26979 44235 26985
rect 44177 26945 44189 26979
rect 44223 26976 44235 26979
rect 44223 26948 45048 26976
rect 44223 26945 44235 26948
rect 44177 26939 44235 26945
rect 43404 26880 44128 26908
rect 43404 26868 43410 26880
rect 44266 26868 44272 26920
rect 44324 26908 44330 26920
rect 44545 26911 44603 26917
rect 44545 26908 44557 26911
rect 44324 26880 44557 26908
rect 44324 26868 44330 26880
rect 44545 26877 44557 26880
rect 44591 26877 44603 26911
rect 44545 26871 44603 26877
rect 44637 26911 44695 26917
rect 44637 26877 44649 26911
rect 44683 26877 44695 26911
rect 44637 26871 44695 26877
rect 44729 26911 44787 26917
rect 44729 26877 44741 26911
rect 44775 26877 44787 26911
rect 44729 26871 44787 26877
rect 37182 26840 37188 26852
rect 36372 26812 37188 26840
rect 37182 26800 37188 26812
rect 37240 26800 37246 26852
rect 42521 26843 42579 26849
rect 42521 26809 42533 26843
rect 42567 26840 42579 26843
rect 43622 26840 43628 26852
rect 42567 26812 43628 26840
rect 42567 26809 42579 26812
rect 42521 26803 42579 26809
rect 43622 26800 43628 26812
rect 43680 26800 43686 26852
rect 44174 26800 44180 26852
rect 44232 26800 44238 26852
rect 38102 26772 38108 26784
rect 36280 26744 38108 26772
rect 35069 26735 35127 26741
rect 38102 26732 38108 26744
rect 38160 26732 38166 26784
rect 38565 26775 38623 26781
rect 38565 26741 38577 26775
rect 38611 26772 38623 26775
rect 38930 26772 38936 26784
rect 38611 26744 38936 26772
rect 38611 26741 38623 26744
rect 38565 26735 38623 26741
rect 38930 26732 38936 26744
rect 38988 26732 38994 26784
rect 42613 26775 42671 26781
rect 42613 26741 42625 26775
rect 42659 26772 42671 26775
rect 42702 26772 42708 26784
rect 42659 26744 42708 26772
rect 42659 26741 42671 26744
rect 42613 26735 42671 26741
rect 42702 26732 42708 26744
rect 42760 26732 42766 26784
rect 43714 26732 43720 26784
rect 43772 26772 43778 26784
rect 44652 26772 44680 26871
rect 44744 26840 44772 26871
rect 44818 26868 44824 26920
rect 44876 26868 44882 26920
rect 45020 26917 45048 26948
rect 45278 26936 45284 26988
rect 45336 26976 45342 26988
rect 45925 26979 45983 26985
rect 45925 26976 45937 26979
rect 45336 26948 45937 26976
rect 45336 26936 45342 26948
rect 45925 26945 45937 26948
rect 45971 26945 45983 26979
rect 45925 26939 45983 26945
rect 45005 26911 45063 26917
rect 45005 26877 45017 26911
rect 45051 26877 45063 26911
rect 45005 26871 45063 26877
rect 48498 26868 48504 26920
rect 48556 26868 48562 26920
rect 48777 26911 48835 26917
rect 48777 26877 48789 26911
rect 48823 26908 48835 26911
rect 49142 26908 49148 26920
rect 48823 26880 49148 26908
rect 48823 26877 48835 26880
rect 48777 26871 48835 26877
rect 49142 26868 49148 26880
rect 49200 26868 49206 26920
rect 50341 26911 50399 26917
rect 50341 26877 50353 26911
rect 50387 26877 50399 26911
rect 50341 26871 50399 26877
rect 50617 26911 50675 26917
rect 50617 26877 50629 26911
rect 50663 26908 50675 26911
rect 51166 26908 51172 26920
rect 50663 26880 51172 26908
rect 50663 26877 50675 26880
rect 50617 26871 50675 26877
rect 45922 26840 45928 26852
rect 44744 26812 45928 26840
rect 45922 26800 45928 26812
rect 45980 26800 45986 26852
rect 43772 26744 44680 26772
rect 43772 26732 43778 26744
rect 49970 26732 49976 26784
rect 50028 26772 50034 26784
rect 50249 26775 50307 26781
rect 50249 26772 50261 26775
rect 50028 26744 50261 26772
rect 50028 26732 50034 26744
rect 50249 26741 50261 26744
rect 50295 26741 50307 26775
rect 50356 26772 50384 26871
rect 51166 26868 51172 26880
rect 51224 26868 51230 26920
rect 51258 26868 51264 26920
rect 51316 26908 51322 26920
rect 52362 26908 52368 26920
rect 51316 26880 52368 26908
rect 51316 26868 51322 26880
rect 52362 26868 52368 26880
rect 52420 26868 52426 26920
rect 54202 26868 54208 26920
rect 54260 26868 54266 26920
rect 54478 26868 54484 26920
rect 54536 26868 54542 26920
rect 51074 26772 51080 26784
rect 50356 26744 51080 26772
rect 50249 26735 50307 26741
rect 51074 26732 51080 26744
rect 51132 26732 51138 26784
rect 52086 26732 52092 26784
rect 52144 26732 52150 26784
rect 52730 26732 52736 26784
rect 52788 26732 52794 26784
rect 1104 26682 78844 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 78844 26682
rect 1104 26608 78844 26630
rect 1302 26528 1308 26580
rect 1360 26568 1366 26580
rect 1857 26571 1915 26577
rect 1857 26568 1869 26571
rect 1360 26540 1869 26568
rect 1360 26528 1366 26540
rect 1857 26537 1869 26540
rect 1903 26537 1915 26571
rect 1857 26531 1915 26537
rect 10962 26528 10968 26580
rect 11020 26568 11026 26580
rect 11793 26571 11851 26577
rect 11793 26568 11805 26571
rect 11020 26540 11805 26568
rect 11020 26528 11026 26540
rect 11793 26537 11805 26540
rect 11839 26537 11851 26571
rect 11793 26531 11851 26537
rect 11974 26528 11980 26580
rect 12032 26528 12038 26580
rect 12345 26571 12403 26577
rect 12345 26537 12357 26571
rect 12391 26568 12403 26571
rect 12434 26568 12440 26580
rect 12391 26540 12440 26568
rect 12391 26537 12403 26540
rect 12345 26531 12403 26537
rect 12434 26528 12440 26540
rect 12492 26528 12498 26580
rect 20346 26528 20352 26580
rect 20404 26528 20410 26580
rect 31021 26571 31079 26577
rect 31021 26537 31033 26571
rect 31067 26568 31079 26571
rect 31110 26568 31116 26580
rect 31067 26540 31116 26568
rect 31067 26537 31079 26540
rect 31021 26531 31079 26537
rect 31110 26528 31116 26540
rect 31168 26568 31174 26580
rect 31662 26568 31668 26580
rect 31168 26540 31668 26568
rect 31168 26528 31174 26540
rect 31662 26528 31668 26540
rect 31720 26568 31726 26580
rect 32217 26571 32275 26577
rect 32217 26568 32229 26571
rect 31720 26540 32229 26568
rect 31720 26528 31726 26540
rect 32217 26537 32229 26540
rect 32263 26537 32275 26571
rect 32217 26531 32275 26537
rect 32490 26528 32496 26580
rect 32548 26568 32554 26580
rect 32677 26571 32735 26577
rect 32677 26568 32689 26571
rect 32548 26540 32689 26568
rect 32548 26528 32554 26540
rect 32677 26537 32689 26540
rect 32723 26537 32735 26571
rect 32677 26531 32735 26537
rect 34146 26528 34152 26580
rect 34204 26568 34210 26580
rect 34701 26571 34759 26577
rect 34701 26568 34713 26571
rect 34204 26540 34713 26568
rect 34204 26528 34210 26540
rect 34701 26537 34713 26540
rect 34747 26537 34759 26571
rect 34701 26531 34759 26537
rect 40402 26528 40408 26580
rect 40460 26528 40466 26580
rect 41138 26528 41144 26580
rect 41196 26568 41202 26580
rect 41233 26571 41291 26577
rect 41233 26568 41245 26571
rect 41196 26540 41245 26568
rect 41196 26528 41202 26540
rect 41233 26537 41245 26540
rect 41279 26537 41291 26571
rect 41233 26531 41291 26537
rect 42794 26528 42800 26580
rect 42852 26568 42858 26580
rect 45833 26571 45891 26577
rect 45833 26568 45845 26571
rect 42852 26540 45845 26568
rect 42852 26528 42858 26540
rect 45833 26537 45845 26540
rect 45879 26537 45891 26571
rect 45833 26531 45891 26537
rect 49142 26528 49148 26580
rect 49200 26528 49206 26580
rect 49605 26571 49663 26577
rect 49605 26537 49617 26571
rect 49651 26568 49663 26571
rect 51534 26568 51540 26580
rect 49651 26540 51540 26568
rect 49651 26537 49663 26540
rect 49605 26531 49663 26537
rect 51534 26528 51540 26540
rect 51592 26568 51598 26580
rect 53561 26571 53619 26577
rect 53561 26568 53573 26571
rect 51592 26540 53573 26568
rect 51592 26528 51598 26540
rect 53561 26537 53573 26540
rect 53607 26537 53619 26571
rect 53561 26531 53619 26537
rect 54021 26571 54079 26577
rect 54021 26537 54033 26571
rect 54067 26568 54079 26571
rect 54202 26568 54208 26580
rect 54067 26540 54208 26568
rect 54067 26537 54079 26540
rect 54021 26531 54079 26537
rect 54202 26528 54208 26540
rect 54260 26528 54266 26580
rect 13354 26500 13360 26512
rect 11256 26472 13360 26500
rect 9953 26435 10011 26441
rect 9953 26401 9965 26435
rect 9999 26432 10011 26435
rect 10226 26432 10232 26444
rect 9999 26404 10232 26432
rect 9999 26401 10011 26404
rect 9953 26395 10011 26401
rect 10226 26392 10232 26404
rect 10284 26392 10290 26444
rect 10686 26392 10692 26444
rect 10744 26432 10750 26444
rect 11256 26432 11284 26472
rect 13354 26460 13360 26472
rect 13412 26460 13418 26512
rect 10744 26404 11284 26432
rect 11701 26435 11759 26441
rect 10744 26392 10750 26404
rect 11701 26401 11713 26435
rect 11747 26432 11759 26435
rect 12526 26432 12532 26444
rect 11747 26404 12532 26432
rect 11747 26401 11759 26404
rect 11701 26395 11759 26401
rect 2038 26324 2044 26376
rect 2096 26324 2102 26376
rect 10134 26256 10140 26308
rect 10192 26296 10198 26308
rect 10229 26299 10287 26305
rect 10229 26296 10241 26299
rect 10192 26268 10241 26296
rect 10192 26256 10198 26268
rect 10229 26265 10241 26268
rect 10275 26265 10287 26299
rect 10229 26259 10287 26265
rect 10318 26256 10324 26308
rect 10376 26296 10382 26308
rect 10686 26296 10692 26308
rect 10376 26268 10692 26296
rect 10376 26256 10382 26268
rect 10686 26256 10692 26268
rect 10744 26256 10750 26308
rect 11992 26305 12020 26404
rect 12526 26392 12532 26404
rect 12584 26432 12590 26444
rect 12894 26432 12900 26444
rect 12584 26404 12900 26432
rect 12584 26392 12590 26404
rect 12894 26392 12900 26404
rect 12952 26392 12958 26444
rect 20257 26435 20315 26441
rect 20257 26401 20269 26435
rect 20303 26432 20315 26435
rect 20622 26432 20628 26444
rect 20303 26404 20628 26432
rect 20303 26401 20315 26404
rect 20257 26395 20315 26401
rect 20622 26392 20628 26404
rect 20680 26392 20686 26444
rect 35345 26435 35403 26441
rect 35345 26432 35357 26435
rect 30760 26404 32536 26432
rect 12066 26324 12072 26376
rect 12124 26364 12130 26376
rect 12253 26367 12311 26373
rect 12253 26364 12265 26367
rect 12124 26336 12265 26364
rect 12124 26324 12130 26336
rect 12253 26333 12265 26336
rect 12299 26333 12311 26367
rect 12434 26364 12440 26376
rect 12253 26327 12311 26333
rect 12406 26324 12440 26364
rect 12492 26364 12498 26376
rect 12986 26364 12992 26376
rect 12492 26336 12992 26364
rect 12492 26324 12498 26336
rect 12986 26324 12992 26336
rect 13044 26324 13050 26376
rect 20073 26367 20131 26373
rect 20073 26333 20085 26367
rect 20119 26364 20131 26367
rect 20162 26364 20168 26376
rect 20119 26336 20168 26364
rect 20119 26333 20131 26336
rect 20073 26327 20131 26333
rect 20162 26324 20168 26336
rect 20220 26324 20226 26376
rect 21913 26367 21971 26373
rect 21913 26333 21925 26367
rect 21959 26333 21971 26367
rect 21913 26327 21971 26333
rect 11961 26299 12020 26305
rect 11961 26265 11973 26299
rect 12007 26268 12020 26299
rect 12007 26265 12019 26268
rect 11961 26259 12019 26265
rect 12158 26256 12164 26308
rect 12216 26296 12222 26308
rect 12406 26296 12434 26324
rect 12216 26268 12434 26296
rect 20349 26299 20407 26305
rect 12216 26256 12222 26268
rect 20349 26265 20361 26299
rect 20395 26296 20407 26299
rect 20714 26296 20720 26308
rect 20395 26268 20720 26296
rect 20395 26265 20407 26268
rect 20349 26259 20407 26265
rect 20714 26256 20720 26268
rect 20772 26296 20778 26308
rect 21928 26296 21956 26327
rect 30374 26324 30380 26376
rect 30432 26364 30438 26376
rect 30760 26373 30788 26404
rect 30745 26367 30803 26373
rect 30745 26364 30757 26367
rect 30432 26336 30757 26364
rect 30432 26324 30438 26336
rect 30745 26333 30757 26336
rect 30791 26333 30803 26367
rect 30745 26327 30803 26333
rect 30834 26324 30840 26376
rect 30892 26324 30898 26376
rect 31113 26367 31171 26373
rect 31113 26333 31125 26367
rect 31159 26364 31171 26367
rect 31570 26364 31576 26376
rect 31159 26336 31576 26364
rect 31159 26333 31171 26336
rect 31113 26327 31171 26333
rect 31570 26324 31576 26336
rect 31628 26324 31634 26376
rect 32122 26373 32128 26376
rect 32113 26367 32128 26373
rect 32113 26333 32125 26367
rect 32113 26327 32128 26333
rect 32122 26324 32128 26327
rect 32180 26324 32186 26376
rect 32398 26324 32404 26376
rect 32456 26324 32462 26376
rect 32508 26373 32536 26404
rect 34900 26404 35357 26432
rect 32493 26367 32551 26373
rect 32493 26333 32505 26367
rect 32539 26364 32551 26367
rect 32582 26364 32588 26376
rect 32539 26336 32588 26364
rect 32539 26333 32551 26336
rect 32493 26327 32551 26333
rect 32582 26324 32588 26336
rect 32640 26324 32646 26376
rect 34606 26324 34612 26376
rect 34664 26364 34670 26376
rect 34900 26373 34928 26404
rect 35345 26401 35357 26404
rect 35391 26401 35403 26435
rect 35345 26395 35403 26401
rect 41049 26435 41107 26441
rect 41049 26401 41061 26435
rect 41095 26432 41107 26435
rect 41156 26432 41184 26528
rect 44082 26460 44088 26512
rect 44140 26500 44146 26512
rect 45005 26503 45063 26509
rect 45005 26500 45017 26503
rect 44140 26472 45017 26500
rect 44140 26460 44146 26472
rect 45005 26469 45017 26472
rect 45051 26469 45063 26503
rect 45005 26463 45063 26469
rect 45465 26503 45523 26509
rect 45465 26469 45477 26503
rect 45511 26500 45523 26503
rect 46014 26500 46020 26512
rect 45511 26472 46020 26500
rect 45511 26469 45523 26472
rect 45465 26463 45523 26469
rect 46014 26460 46020 26472
rect 46072 26460 46078 26512
rect 49510 26500 49516 26512
rect 48792 26472 49516 26500
rect 45830 26432 45836 26444
rect 41095 26404 41184 26432
rect 44284 26404 45416 26432
rect 41095 26401 41107 26404
rect 41049 26395 41107 26401
rect 34885 26367 34943 26373
rect 34885 26364 34897 26367
rect 34664 26336 34897 26364
rect 34664 26324 34670 26336
rect 34885 26333 34897 26336
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 35253 26367 35311 26373
rect 35253 26333 35265 26367
rect 35299 26364 35311 26367
rect 36538 26364 36544 26376
rect 35299 26336 36544 26364
rect 35299 26333 35311 26336
rect 35253 26327 35311 26333
rect 36538 26324 36544 26336
rect 36596 26324 36602 26376
rect 40773 26367 40831 26373
rect 40773 26333 40785 26367
rect 40819 26364 40831 26367
rect 41230 26364 41236 26376
rect 40819 26336 41236 26364
rect 40819 26333 40831 26336
rect 40773 26327 40831 26333
rect 41230 26324 41236 26336
rect 41288 26324 41294 26376
rect 43622 26324 43628 26376
rect 43680 26364 43686 26376
rect 44284 26373 44312 26404
rect 44085 26367 44143 26373
rect 44085 26364 44097 26367
rect 43680 26336 44097 26364
rect 43680 26324 43686 26336
rect 44085 26333 44097 26336
rect 44131 26333 44143 26367
rect 44085 26327 44143 26333
rect 44269 26367 44327 26373
rect 44269 26333 44281 26367
rect 44315 26333 44327 26367
rect 44269 26327 44327 26333
rect 44637 26367 44695 26373
rect 44637 26333 44649 26367
rect 44683 26364 44695 26367
rect 44726 26364 44732 26376
rect 44683 26336 44732 26364
rect 44683 26333 44695 26336
rect 44637 26327 44695 26333
rect 44726 26324 44732 26336
rect 44784 26324 44790 26376
rect 44821 26367 44879 26373
rect 44821 26333 44833 26367
rect 44867 26364 44879 26367
rect 45002 26364 45008 26376
rect 44867 26336 45008 26364
rect 44867 26333 44879 26336
rect 44821 26327 44879 26333
rect 45002 26324 45008 26336
rect 45060 26324 45066 26376
rect 45388 26373 45416 26404
rect 45756 26404 45836 26432
rect 45281 26367 45339 26373
rect 45281 26333 45293 26367
rect 45327 26333 45339 26367
rect 45281 26327 45339 26333
rect 45373 26367 45431 26373
rect 45373 26333 45385 26367
rect 45419 26333 45431 26367
rect 45373 26327 45431 26333
rect 20772 26268 21956 26296
rect 20772 26256 20778 26268
rect 34514 26256 34520 26308
rect 34572 26296 34578 26308
rect 34977 26299 35035 26305
rect 34977 26296 34989 26299
rect 34572 26268 34989 26296
rect 34572 26256 34578 26268
rect 34977 26265 34989 26268
rect 35023 26265 35035 26299
rect 34977 26259 35035 26265
rect 35066 26256 35072 26308
rect 35124 26296 35130 26308
rect 35618 26296 35624 26308
rect 35124 26268 35624 26296
rect 35124 26256 35130 26268
rect 35618 26256 35624 26268
rect 35676 26256 35682 26308
rect 44450 26256 44456 26308
rect 44508 26256 44514 26308
rect 45296 26296 45324 26327
rect 44836 26268 45324 26296
rect 45388 26296 45416 26327
rect 45462 26324 45468 26376
rect 45520 26364 45526 26376
rect 45756 26373 45784 26404
rect 45830 26392 45836 26404
rect 45888 26432 45894 26444
rect 46385 26435 46443 26441
rect 46385 26432 46397 26435
rect 45888 26404 46397 26432
rect 45888 26392 45894 26404
rect 46385 26401 46397 26404
rect 46431 26401 46443 26435
rect 46385 26395 46443 26401
rect 48498 26392 48504 26444
rect 48556 26432 48562 26444
rect 48792 26441 48820 26472
rect 49510 26460 49516 26472
rect 49568 26500 49574 26512
rect 51074 26500 51080 26512
rect 49568 26472 51080 26500
rect 49568 26460 49574 26472
rect 51074 26460 51080 26472
rect 51132 26500 51138 26512
rect 54478 26500 54484 26512
rect 51132 26472 54484 26500
rect 51132 26460 51138 26472
rect 48777 26435 48835 26441
rect 48777 26432 48789 26435
rect 48556 26404 48789 26432
rect 48556 26392 48562 26404
rect 48777 26401 48789 26404
rect 48823 26401 48835 26435
rect 48777 26395 48835 26401
rect 49970 26392 49976 26444
rect 50028 26432 50034 26444
rect 50709 26435 50767 26441
rect 50709 26432 50721 26435
rect 50028 26404 50721 26432
rect 50028 26392 50034 26404
rect 50709 26401 50721 26404
rect 50755 26401 50767 26435
rect 52270 26432 52276 26444
rect 50709 26395 50767 26401
rect 51092 26404 52276 26432
rect 45557 26367 45615 26373
rect 45557 26364 45569 26367
rect 45520 26336 45569 26364
rect 45520 26324 45526 26336
rect 45557 26333 45569 26336
rect 45603 26333 45615 26367
rect 45557 26327 45615 26333
rect 45741 26367 45799 26373
rect 45741 26333 45753 26367
rect 45787 26333 45799 26367
rect 45741 26327 45799 26333
rect 45958 26367 46016 26373
rect 45958 26333 45970 26367
rect 46004 26364 46016 26367
rect 46004 26336 46244 26364
rect 46004 26333 46016 26336
rect 45958 26327 46016 26333
rect 46106 26305 46112 26308
rect 46083 26299 46112 26305
rect 46083 26296 46095 26299
rect 45388 26268 46095 26296
rect 44836 26240 44864 26268
rect 46083 26265 46095 26268
rect 46083 26259 46112 26265
rect 46106 26256 46112 26259
rect 46164 26256 46170 26308
rect 19426 26188 19432 26240
rect 19484 26228 19490 26240
rect 19889 26231 19947 26237
rect 19889 26228 19901 26231
rect 19484 26200 19901 26228
rect 19484 26188 19490 26200
rect 19889 26197 19901 26200
rect 19935 26197 19947 26231
rect 19889 26191 19947 26197
rect 21358 26188 21364 26240
rect 21416 26188 21422 26240
rect 30558 26188 30564 26240
rect 30616 26188 30622 26240
rect 40862 26188 40868 26240
rect 40920 26188 40926 26240
rect 44729 26231 44787 26237
rect 44729 26197 44741 26231
rect 44775 26228 44787 26231
rect 44818 26228 44824 26240
rect 44775 26200 44824 26228
rect 44775 26197 44787 26200
rect 44729 26191 44787 26197
rect 44818 26188 44824 26200
rect 44876 26188 44882 26240
rect 45278 26188 45284 26240
rect 45336 26228 45342 26240
rect 46216 26228 46244 26336
rect 46474 26324 46480 26376
rect 46532 26324 46538 26376
rect 49326 26324 49332 26376
rect 49384 26324 49390 26376
rect 49421 26367 49479 26373
rect 49421 26333 49433 26367
rect 49467 26333 49479 26367
rect 49421 26327 49479 26333
rect 49697 26367 49755 26373
rect 49697 26333 49709 26367
rect 49743 26364 49755 26367
rect 50157 26367 50215 26373
rect 50157 26364 50169 26367
rect 49743 26336 50169 26364
rect 49743 26333 49755 26336
rect 49697 26327 49755 26333
rect 50157 26333 50169 26336
rect 50203 26333 50215 26367
rect 50724 26364 50752 26395
rect 51092 26373 51120 26404
rect 52270 26392 52276 26404
rect 52328 26392 52334 26444
rect 52380 26441 52408 26472
rect 54478 26460 54484 26472
rect 54536 26460 54542 26512
rect 52365 26435 52423 26441
rect 52365 26401 52377 26435
rect 52411 26401 52423 26435
rect 52365 26395 52423 26401
rect 52454 26392 52460 26444
rect 52512 26432 52518 26444
rect 52512 26404 53880 26432
rect 52512 26392 52518 26404
rect 50893 26367 50951 26373
rect 50893 26364 50905 26367
rect 50724 26336 50905 26364
rect 50157 26327 50215 26333
rect 50893 26333 50905 26336
rect 50939 26333 50951 26367
rect 50893 26327 50951 26333
rect 51077 26367 51135 26373
rect 51077 26333 51089 26367
rect 51123 26333 51135 26367
rect 51077 26327 51135 26333
rect 51261 26367 51319 26373
rect 51261 26333 51273 26367
rect 51307 26364 51319 26367
rect 51350 26364 51356 26376
rect 51307 26336 51356 26364
rect 51307 26333 51319 26336
rect 51261 26327 51319 26333
rect 46750 26256 46756 26308
rect 46808 26256 46814 26308
rect 48406 26296 48412 26308
rect 48070 26268 48412 26296
rect 48406 26256 48412 26268
rect 48464 26256 48470 26308
rect 48498 26256 48504 26308
rect 48556 26256 48562 26308
rect 49436 26296 49464 26327
rect 51350 26324 51356 26336
rect 51408 26324 51414 26376
rect 52730 26364 52736 26376
rect 51552 26336 52736 26364
rect 49878 26296 49884 26308
rect 49436 26268 49884 26296
rect 49878 26256 49884 26268
rect 49936 26256 49942 26308
rect 50798 26256 50804 26308
rect 50856 26296 50862 26308
rect 51169 26299 51227 26305
rect 51169 26296 51181 26299
rect 50856 26268 51181 26296
rect 50856 26256 50862 26268
rect 51169 26265 51181 26268
rect 51215 26296 51227 26299
rect 51552 26296 51580 26336
rect 52730 26324 52736 26336
rect 52788 26324 52794 26376
rect 53377 26367 53435 26373
rect 53377 26333 53389 26367
rect 53423 26364 53435 26367
rect 53469 26367 53527 26373
rect 53469 26364 53481 26367
rect 53423 26336 53481 26364
rect 53423 26333 53435 26336
rect 53377 26327 53435 26333
rect 53469 26333 53481 26336
rect 53515 26333 53527 26367
rect 53469 26327 53527 26333
rect 53742 26324 53748 26376
rect 53800 26324 53806 26376
rect 53852 26373 53880 26404
rect 53837 26367 53895 26373
rect 53837 26333 53849 26367
rect 53883 26333 53895 26367
rect 53837 26327 53895 26333
rect 51215 26268 51580 26296
rect 51629 26299 51687 26305
rect 51215 26265 51227 26268
rect 51169 26259 51227 26265
rect 51629 26265 51641 26299
rect 51675 26296 51687 26299
rect 51810 26296 51816 26308
rect 51675 26268 51816 26296
rect 51675 26265 51687 26268
rect 51629 26259 51687 26265
rect 51810 26256 51816 26268
rect 51868 26256 51874 26308
rect 52454 26256 52460 26308
rect 52512 26296 52518 26308
rect 53006 26296 53012 26308
rect 52512 26268 53012 26296
rect 52512 26256 52518 26268
rect 53006 26256 53012 26268
rect 53064 26256 53070 26308
rect 45336 26200 46244 26228
rect 45336 26188 45342 26200
rect 51442 26188 51448 26240
rect 51500 26188 51506 26240
rect 1104 26138 78844 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 66314 26138
rect 66366 26086 66378 26138
rect 66430 26086 66442 26138
rect 66494 26086 66506 26138
rect 66558 26086 66570 26138
rect 66622 26086 78844 26138
rect 1104 26064 78844 26086
rect 934 25984 940 26036
rect 992 26024 998 26036
rect 1857 26027 1915 26033
rect 1857 26024 1869 26027
rect 992 25996 1869 26024
rect 992 25984 998 25996
rect 1857 25993 1869 25996
rect 1903 25993 1915 26027
rect 1857 25987 1915 25993
rect 10042 25984 10048 26036
rect 10100 26024 10106 26036
rect 12986 26024 12992 26036
rect 10100 25996 12992 26024
rect 10100 25984 10106 25996
rect 12986 25984 12992 25996
rect 13044 26024 13050 26036
rect 15470 26024 15476 26036
rect 13044 25996 15476 26024
rect 13044 25984 13050 25996
rect 15470 25984 15476 25996
rect 15528 26024 15534 26036
rect 15749 26027 15807 26033
rect 15749 26024 15761 26027
rect 15528 25996 15761 26024
rect 15528 25984 15534 25996
rect 15749 25993 15761 25996
rect 15795 25993 15807 26027
rect 15749 25987 15807 25993
rect 16942 25984 16948 26036
rect 17000 26024 17006 26036
rect 17865 26027 17923 26033
rect 17865 26024 17877 26027
rect 17000 25996 17877 26024
rect 17000 25984 17006 25996
rect 17865 25993 17877 25996
rect 17911 26024 17923 26027
rect 17954 26024 17960 26036
rect 17911 25996 17960 26024
rect 17911 25993 17923 25996
rect 17865 25987 17923 25993
rect 17954 25984 17960 25996
rect 18012 25984 18018 26036
rect 29178 25984 29184 26036
rect 29236 26024 29242 26036
rect 31386 26024 31392 26036
rect 29236 25996 31392 26024
rect 29236 25984 29242 25996
rect 15102 25916 15108 25968
rect 15160 25916 15166 25968
rect 19426 25956 19432 25968
rect 17328 25928 19432 25956
rect 2041 25891 2099 25897
rect 2041 25857 2053 25891
rect 2087 25888 2099 25891
rect 2133 25891 2191 25897
rect 2133 25888 2145 25891
rect 2087 25860 2145 25888
rect 2087 25857 2099 25860
rect 2041 25851 2099 25857
rect 2133 25857 2145 25860
rect 2179 25857 2191 25891
rect 17328 25888 17356 25928
rect 19426 25916 19432 25928
rect 19484 25916 19490 25968
rect 19705 25959 19763 25965
rect 19705 25925 19717 25959
rect 19751 25956 19763 25959
rect 21358 25956 21364 25968
rect 19751 25928 21364 25956
rect 19751 25925 19763 25928
rect 19705 25919 19763 25925
rect 2133 25851 2191 25857
rect 15488 25860 17356 25888
rect 17405 25891 17463 25897
rect 15488 25829 15516 25860
rect 17405 25857 17417 25891
rect 17451 25888 17463 25891
rect 17586 25888 17592 25900
rect 17451 25860 17592 25888
rect 17451 25857 17463 25860
rect 17405 25851 17463 25857
rect 17586 25848 17592 25860
rect 17644 25848 17650 25900
rect 17681 25891 17739 25897
rect 17681 25857 17693 25891
rect 17727 25888 17739 25891
rect 17954 25888 17960 25900
rect 17727 25860 17960 25888
rect 17727 25857 17739 25860
rect 17681 25851 17739 25857
rect 17954 25848 17960 25860
rect 18012 25848 18018 25900
rect 19518 25848 19524 25900
rect 19576 25888 19582 25900
rect 19613 25891 19671 25897
rect 19613 25888 19625 25891
rect 19576 25860 19625 25888
rect 19576 25848 19582 25860
rect 19613 25857 19625 25860
rect 19659 25857 19671 25891
rect 19613 25851 19671 25857
rect 19889 25891 19947 25897
rect 19889 25857 19901 25891
rect 19935 25888 19947 25891
rect 20349 25891 20407 25897
rect 20349 25888 20361 25891
rect 19935 25860 20361 25888
rect 19935 25857 19947 25860
rect 19889 25851 19947 25857
rect 20349 25857 20361 25860
rect 20395 25857 20407 25891
rect 20349 25851 20407 25857
rect 15473 25823 15531 25829
rect 15473 25789 15485 25823
rect 15519 25789 15531 25823
rect 15473 25783 15531 25789
rect 17310 25780 17316 25832
rect 17368 25820 17374 25832
rect 17497 25823 17555 25829
rect 17497 25820 17509 25823
rect 17368 25792 17509 25820
rect 17368 25780 17374 25792
rect 17497 25789 17509 25792
rect 17543 25789 17555 25823
rect 19628 25820 19656 25851
rect 20622 25848 20628 25900
rect 20680 25888 20686 25900
rect 21284 25897 21312 25928
rect 21358 25916 21364 25928
rect 21416 25916 21422 25968
rect 22830 25916 22836 25968
rect 22888 25956 22894 25968
rect 30392 25956 30420 25996
rect 31386 25984 31392 25996
rect 31444 26024 31450 26036
rect 31757 26027 31815 26033
rect 31757 26024 31769 26027
rect 31444 25996 31769 26024
rect 31444 25984 31450 25996
rect 31757 25993 31769 25996
rect 31803 25993 31815 26027
rect 31757 25987 31815 25993
rect 32398 25984 32404 26036
rect 32456 25984 32462 26036
rect 37274 25984 37280 26036
rect 37332 26024 37338 26036
rect 37734 26024 37740 26036
rect 37332 25996 37740 26024
rect 37332 25984 37338 25996
rect 37734 25984 37740 25996
rect 37792 26024 37798 26036
rect 37829 26027 37887 26033
rect 37829 26024 37841 26027
rect 37792 25996 37841 26024
rect 37792 25984 37798 25996
rect 37829 25993 37841 25996
rect 37875 25993 37887 26027
rect 37829 25987 37887 25993
rect 38378 25984 38384 26036
rect 38436 26024 38442 26036
rect 38565 26027 38623 26033
rect 38565 26024 38577 26027
rect 38436 25996 38577 26024
rect 38436 25984 38442 25996
rect 38565 25993 38577 25996
rect 38611 25993 38623 26027
rect 38565 25987 38623 25993
rect 40862 25984 40868 26036
rect 40920 25984 40926 26036
rect 42889 26027 42947 26033
rect 42889 25993 42901 26027
rect 42935 26024 42947 26027
rect 43070 26024 43076 26036
rect 42935 25996 43076 26024
rect 42935 25993 42947 25996
rect 42889 25987 42947 25993
rect 43070 25984 43076 25996
rect 43128 25984 43134 26036
rect 46474 25984 46480 26036
rect 46532 26024 46538 26036
rect 46569 26027 46627 26033
rect 46569 26024 46581 26027
rect 46532 25996 46581 26024
rect 46532 25984 46538 25996
rect 46569 25993 46581 25996
rect 46615 25993 46627 26027
rect 46569 25987 46627 25993
rect 46750 25984 46756 26036
rect 46808 26024 46814 26036
rect 47949 26027 48007 26033
rect 47949 26024 47961 26027
rect 46808 25996 47961 26024
rect 46808 25984 46814 25996
rect 47949 25993 47961 25996
rect 47995 25993 48007 26027
rect 47949 25987 48007 25993
rect 48317 26027 48375 26033
rect 48317 25993 48329 26027
rect 48363 26024 48375 26027
rect 48498 26024 48504 26036
rect 48363 25996 48504 26024
rect 48363 25993 48375 25996
rect 48317 25987 48375 25993
rect 48498 25984 48504 25996
rect 48556 25984 48562 26036
rect 49878 25984 49884 26036
rect 49936 25984 49942 26036
rect 51074 25984 51080 26036
rect 51132 25984 51138 26036
rect 51350 25984 51356 26036
rect 51408 25984 51414 26036
rect 53285 26027 53343 26033
rect 53285 25993 53297 26027
rect 53331 26024 53343 26027
rect 53742 26024 53748 26036
rect 53331 25996 53748 26024
rect 53331 25993 53343 25996
rect 53285 25987 53343 25993
rect 53742 25984 53748 25996
rect 53800 25984 53806 26036
rect 31570 25965 31576 25968
rect 31527 25959 31576 25965
rect 31527 25956 31539 25959
rect 22888 25928 23796 25956
rect 30392 25928 30498 25956
rect 31483 25928 31539 25956
rect 22888 25916 22894 25928
rect 20901 25891 20959 25897
rect 20901 25888 20913 25891
rect 20680 25860 20913 25888
rect 20680 25848 20686 25860
rect 20901 25857 20913 25860
rect 20947 25857 20959 25891
rect 20901 25851 20959 25857
rect 21269 25891 21327 25897
rect 21269 25857 21281 25891
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 20070 25820 20076 25832
rect 19628 25792 20076 25820
rect 17497 25783 17555 25789
rect 20070 25780 20076 25792
rect 20128 25820 20134 25832
rect 21177 25823 21235 25829
rect 21177 25820 21189 25823
rect 20128 25792 21189 25820
rect 20128 25780 20134 25792
rect 21177 25789 21189 25792
rect 21223 25789 21235 25823
rect 21177 25783 21235 25789
rect 21637 25823 21695 25829
rect 21637 25789 21649 25823
rect 21683 25820 21695 25823
rect 23293 25823 23351 25829
rect 23293 25820 23305 25823
rect 21683 25792 23305 25820
rect 21683 25789 21695 25792
rect 21637 25783 21695 25789
rect 23293 25789 23305 25792
rect 23339 25789 23351 25823
rect 23293 25783 23351 25789
rect 23566 25780 23572 25832
rect 23624 25780 23630 25832
rect 15381 25755 15439 25761
rect 15381 25721 15393 25755
rect 15427 25752 15439 25755
rect 17221 25755 17279 25761
rect 17221 25752 17233 25755
rect 15427 25724 17233 25752
rect 15427 25721 15439 25724
rect 15381 25715 15439 25721
rect 17221 25721 17233 25724
rect 17267 25721 17279 25755
rect 17221 25715 17279 25721
rect 20714 25712 20720 25764
rect 20772 25752 20778 25764
rect 23768 25761 23796 25928
rect 31527 25925 31539 25928
rect 31573 25925 31576 25959
rect 31527 25919 31576 25925
rect 31570 25916 31576 25919
rect 31628 25956 31634 25968
rect 32677 25959 32735 25965
rect 32677 25956 32689 25959
rect 31628 25928 32689 25956
rect 31628 25916 31634 25928
rect 32677 25925 32689 25928
rect 32723 25925 32735 25959
rect 34790 25956 34796 25968
rect 32677 25919 32735 25925
rect 32784 25928 34796 25956
rect 32582 25848 32588 25900
rect 32640 25848 32646 25900
rect 32784 25897 32812 25928
rect 34790 25916 34796 25928
rect 34848 25956 34854 25968
rect 35066 25956 35072 25968
rect 34848 25928 35072 25956
rect 34848 25916 34854 25928
rect 35066 25916 35072 25928
rect 35124 25916 35130 25968
rect 38197 25959 38255 25965
rect 38197 25956 38209 25959
rect 37568 25928 38209 25956
rect 32769 25891 32827 25897
rect 32769 25857 32781 25891
rect 32815 25857 32827 25891
rect 32769 25851 32827 25857
rect 32953 25891 33011 25897
rect 32953 25857 32965 25891
rect 32999 25888 33011 25891
rect 32999 25860 34008 25888
rect 32999 25857 33011 25860
rect 32953 25851 33011 25857
rect 28442 25780 28448 25832
rect 28500 25820 28506 25832
rect 29733 25823 29791 25829
rect 29733 25820 29745 25823
rect 28500 25792 29745 25820
rect 28500 25780 28506 25792
rect 29733 25789 29745 25792
rect 29779 25789 29791 25823
rect 29733 25783 29791 25789
rect 30101 25823 30159 25829
rect 30101 25789 30113 25823
rect 30147 25820 30159 25823
rect 30558 25820 30564 25832
rect 30147 25792 30564 25820
rect 30147 25789 30159 25792
rect 30101 25783 30159 25789
rect 30558 25780 30564 25792
rect 30616 25780 30622 25832
rect 31386 25780 31392 25832
rect 31444 25820 31450 25832
rect 32784 25820 32812 25851
rect 31444 25792 32812 25820
rect 31444 25780 31450 25792
rect 21821 25755 21879 25761
rect 21821 25752 21833 25755
rect 20772 25724 21833 25752
rect 20772 25712 20778 25724
rect 21821 25721 21833 25724
rect 21867 25721 21879 25755
rect 21821 25715 21879 25721
rect 23753 25755 23811 25761
rect 23753 25721 23765 25755
rect 23799 25752 23811 25755
rect 29178 25752 29184 25764
rect 23799 25724 29184 25752
rect 23799 25721 23811 25724
rect 23753 25715 23811 25721
rect 29178 25712 29184 25724
rect 29236 25712 29242 25764
rect 14550 25644 14556 25696
rect 14608 25684 14614 25696
rect 15243 25687 15301 25693
rect 15243 25684 15255 25687
rect 14608 25656 15255 25684
rect 14608 25644 14614 25656
rect 15243 25653 15255 25656
rect 15289 25653 15301 25687
rect 15243 25647 15301 25653
rect 17678 25644 17684 25696
rect 17736 25644 17742 25696
rect 19058 25644 19064 25696
rect 19116 25684 19122 25696
rect 19889 25687 19947 25693
rect 19889 25684 19901 25687
rect 19116 25656 19901 25684
rect 19116 25644 19122 25656
rect 19889 25653 19901 25656
rect 19935 25653 19947 25687
rect 33980 25684 34008 25860
rect 34054 25848 34060 25900
rect 34112 25888 34118 25900
rect 34517 25891 34575 25897
rect 34517 25888 34529 25891
rect 34112 25860 34529 25888
rect 34112 25848 34118 25860
rect 34517 25857 34529 25860
rect 34563 25888 34575 25891
rect 36630 25888 36636 25900
rect 34563 25860 36636 25888
rect 34563 25857 34575 25860
rect 34517 25851 34575 25857
rect 36630 25848 36636 25860
rect 36688 25888 36694 25900
rect 37366 25888 37372 25900
rect 36688 25860 37372 25888
rect 36688 25848 36694 25860
rect 37366 25848 37372 25860
rect 37424 25848 37430 25900
rect 37461 25891 37519 25897
rect 37461 25857 37473 25891
rect 37507 25888 37519 25891
rect 37568 25888 37596 25928
rect 38197 25925 38209 25928
rect 38243 25925 38255 25959
rect 43162 25956 43168 25968
rect 38197 25919 38255 25925
rect 42628 25928 43168 25956
rect 37507 25860 37596 25888
rect 37507 25857 37519 25860
rect 37461 25851 37519 25857
rect 34238 25780 34244 25832
rect 34296 25780 34302 25832
rect 37568 25752 37596 25860
rect 37645 25891 37703 25897
rect 37645 25857 37657 25891
rect 37691 25857 37703 25891
rect 37645 25851 37703 25857
rect 37660 25820 37688 25851
rect 37734 25848 37740 25900
rect 37792 25848 37798 25900
rect 38013 25891 38071 25897
rect 38013 25888 38025 25891
rect 37844 25860 38025 25888
rect 37844 25820 37872 25860
rect 38013 25857 38025 25860
rect 38059 25857 38071 25891
rect 38013 25851 38071 25857
rect 38102 25848 38108 25900
rect 38160 25888 38166 25900
rect 42628 25897 42656 25928
rect 43162 25916 43168 25928
rect 43220 25916 43226 25968
rect 45002 25956 45008 25968
rect 44652 25928 45008 25956
rect 38289 25891 38347 25897
rect 38289 25888 38301 25891
rect 38160 25860 38301 25888
rect 38160 25848 38166 25860
rect 38289 25857 38301 25860
rect 38335 25857 38347 25891
rect 38289 25851 38347 25857
rect 38381 25891 38439 25897
rect 38381 25857 38393 25891
rect 38427 25857 38439 25891
rect 38381 25851 38439 25857
rect 40773 25891 40831 25897
rect 40773 25857 40785 25891
rect 40819 25888 40831 25891
rect 42613 25891 42671 25897
rect 40819 25860 41276 25888
rect 40819 25857 40831 25860
rect 40773 25851 40831 25857
rect 37660 25792 37872 25820
rect 37642 25752 37648 25764
rect 37568 25724 37648 25752
rect 37642 25712 37648 25724
rect 37700 25712 37706 25764
rect 37844 25752 37872 25792
rect 37918 25780 37924 25832
rect 37976 25820 37982 25832
rect 38396 25820 38424 25851
rect 41248 25832 41276 25860
rect 42613 25857 42625 25891
rect 42659 25857 42671 25891
rect 42613 25851 42671 25857
rect 42705 25891 42763 25897
rect 42705 25857 42717 25891
rect 42751 25888 42763 25891
rect 42794 25888 42800 25900
rect 42751 25860 42800 25888
rect 42751 25857 42763 25860
rect 42705 25851 42763 25857
rect 42794 25848 42800 25860
rect 42852 25848 42858 25900
rect 44542 25848 44548 25900
rect 44600 25848 44606 25900
rect 44652 25897 44680 25928
rect 45002 25916 45008 25928
rect 45060 25956 45066 25968
rect 45462 25956 45468 25968
rect 45060 25928 45468 25956
rect 45060 25916 45066 25928
rect 45462 25916 45468 25928
rect 45520 25956 45526 25968
rect 46109 25959 46167 25965
rect 46109 25956 46121 25959
rect 45520 25928 46121 25956
rect 45520 25916 45526 25928
rect 46109 25925 46121 25928
rect 46155 25925 46167 25959
rect 51368 25956 51396 25984
rect 46109 25919 46167 25925
rect 51046 25928 51396 25956
rect 44637 25891 44695 25897
rect 44637 25857 44649 25891
rect 44683 25857 44695 25891
rect 44637 25851 44695 25857
rect 44818 25848 44824 25900
rect 44876 25848 44882 25900
rect 44913 25891 44971 25897
rect 44913 25857 44925 25891
rect 44959 25888 44971 25891
rect 45278 25888 45284 25900
rect 44959 25860 45284 25888
rect 44959 25857 44971 25860
rect 44913 25851 44971 25857
rect 45278 25848 45284 25860
rect 45336 25848 45342 25900
rect 49142 25848 49148 25900
rect 49200 25888 49206 25900
rect 49329 25891 49387 25897
rect 49329 25888 49341 25891
rect 49200 25860 49341 25888
rect 49200 25848 49206 25860
rect 49329 25857 49341 25860
rect 49375 25857 49387 25891
rect 49329 25851 49387 25857
rect 49418 25848 49424 25900
rect 49476 25888 49482 25900
rect 49513 25891 49571 25897
rect 49513 25888 49525 25891
rect 49476 25860 49525 25888
rect 49476 25848 49482 25860
rect 49513 25857 49525 25860
rect 49559 25857 49571 25891
rect 49513 25851 49571 25857
rect 49605 25891 49663 25897
rect 49605 25857 49617 25891
rect 49651 25857 49663 25891
rect 49605 25851 49663 25857
rect 49697 25891 49755 25897
rect 49697 25857 49709 25891
rect 49743 25888 49755 25891
rect 51046 25888 51074 25928
rect 52546 25916 52552 25968
rect 52604 25956 52610 25968
rect 53009 25959 53067 25965
rect 53009 25956 53021 25959
rect 52604 25928 53021 25956
rect 52604 25916 52610 25928
rect 53009 25925 53021 25928
rect 53055 25925 53067 25959
rect 53009 25919 53067 25925
rect 49743 25860 51074 25888
rect 49743 25857 49755 25860
rect 49697 25851 49755 25857
rect 37976 25792 38424 25820
rect 37976 25780 37982 25792
rect 41230 25780 41236 25832
rect 41288 25820 41294 25832
rect 47397 25823 47455 25829
rect 41288 25792 41414 25820
rect 41288 25780 41294 25792
rect 38746 25752 38752 25764
rect 37844 25724 38752 25752
rect 38746 25712 38752 25724
rect 38804 25712 38810 25764
rect 41386 25752 41414 25792
rect 47397 25789 47409 25823
rect 47443 25820 47455 25823
rect 47670 25820 47676 25832
rect 47443 25792 47676 25820
rect 47443 25789 47455 25792
rect 47397 25783 47455 25789
rect 47670 25780 47676 25792
rect 47728 25780 47734 25832
rect 47857 25823 47915 25829
rect 47857 25789 47869 25823
rect 47903 25820 47915 25823
rect 47946 25820 47952 25832
rect 47903 25792 47952 25820
rect 47903 25789 47915 25792
rect 47857 25783 47915 25789
rect 47946 25780 47952 25792
rect 48004 25780 48010 25832
rect 49620 25820 49648 25851
rect 51166 25848 51172 25900
rect 51224 25888 51230 25900
rect 51261 25891 51319 25897
rect 51261 25888 51273 25891
rect 51224 25860 51273 25888
rect 51224 25848 51230 25860
rect 51261 25857 51273 25860
rect 51307 25857 51319 25891
rect 51261 25851 51319 25857
rect 51353 25891 51411 25897
rect 51353 25857 51365 25891
rect 51399 25888 51411 25891
rect 51442 25888 51448 25900
rect 51399 25860 51448 25888
rect 51399 25857 51411 25860
rect 51353 25851 51411 25857
rect 51442 25848 51448 25860
rect 51500 25848 51506 25900
rect 51629 25891 51687 25897
rect 51629 25857 51641 25891
rect 51675 25888 51687 25891
rect 52086 25888 52092 25900
rect 51675 25860 52092 25888
rect 51675 25857 51687 25860
rect 51629 25851 51687 25857
rect 49620 25792 51212 25820
rect 51184 25764 51212 25792
rect 51534 25780 51540 25832
rect 51592 25780 51598 25832
rect 44174 25752 44180 25764
rect 41386 25724 44180 25752
rect 44174 25712 44180 25724
rect 44232 25712 44238 25764
rect 44726 25712 44732 25764
rect 44784 25752 44790 25764
rect 46477 25755 46535 25761
rect 46477 25752 46489 25755
rect 44784 25724 46489 25752
rect 44784 25712 44790 25724
rect 46477 25721 46489 25724
rect 46523 25752 46535 25755
rect 46750 25752 46756 25764
rect 46523 25724 46756 25752
rect 46523 25721 46535 25724
rect 46477 25715 46535 25721
rect 46750 25712 46756 25724
rect 46808 25712 46814 25764
rect 51166 25712 51172 25764
rect 51224 25752 51230 25764
rect 51644 25752 51672 25851
rect 52086 25848 52092 25860
rect 52144 25888 52150 25900
rect 52733 25891 52791 25897
rect 52733 25888 52745 25891
rect 52144 25860 52745 25888
rect 52144 25848 52150 25860
rect 52733 25857 52745 25860
rect 52779 25857 52791 25891
rect 52733 25851 52791 25857
rect 52917 25891 52975 25897
rect 52917 25857 52929 25891
rect 52963 25857 52975 25891
rect 52917 25851 52975 25857
rect 53101 25891 53159 25897
rect 53101 25857 53113 25891
rect 53147 25857 53159 25891
rect 53101 25851 53159 25857
rect 52932 25820 52960 25851
rect 53006 25820 53012 25832
rect 52932 25792 53012 25820
rect 53006 25780 53012 25792
rect 53064 25780 53070 25832
rect 53116 25752 53144 25851
rect 53377 25755 53435 25761
rect 53377 25752 53389 25755
rect 51224 25724 51672 25752
rect 51736 25724 53389 25752
rect 51224 25712 51230 25724
rect 34698 25684 34704 25696
rect 33980 25656 34704 25684
rect 19889 25647 19947 25653
rect 34698 25644 34704 25656
rect 34756 25644 34762 25696
rect 37274 25644 37280 25696
rect 37332 25644 37338 25696
rect 44358 25644 44364 25696
rect 44416 25644 44422 25696
rect 50522 25644 50528 25696
rect 50580 25684 50586 25696
rect 51736 25684 51764 25724
rect 53377 25721 53389 25724
rect 53423 25721 53435 25755
rect 53377 25715 53435 25721
rect 50580 25656 51764 25684
rect 50580 25644 50586 25656
rect 51810 25644 51816 25696
rect 51868 25644 51874 25696
rect 1104 25594 78844 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 78844 25594
rect 1104 25520 78844 25542
rect 13265 25483 13323 25489
rect 13265 25449 13277 25483
rect 13311 25480 13323 25483
rect 13814 25480 13820 25492
rect 13311 25452 13820 25480
rect 13311 25449 13323 25452
rect 13265 25443 13323 25449
rect 13814 25440 13820 25452
rect 13872 25440 13878 25492
rect 14277 25483 14335 25489
rect 14277 25449 14289 25483
rect 14323 25449 14335 25483
rect 14277 25443 14335 25449
rect 13449 25415 13507 25421
rect 13449 25381 13461 25415
rect 13495 25412 13507 25415
rect 13495 25384 14228 25412
rect 13495 25381 13507 25384
rect 13449 25375 13507 25381
rect 12434 25304 12440 25356
rect 12492 25344 12498 25356
rect 14200 25353 14228 25384
rect 12805 25347 12863 25353
rect 12805 25344 12817 25347
rect 12492 25316 12817 25344
rect 12492 25304 12498 25316
rect 12805 25313 12817 25316
rect 12851 25313 12863 25347
rect 12805 25307 12863 25313
rect 14185 25347 14243 25353
rect 14185 25313 14197 25347
rect 14231 25313 14243 25347
rect 14185 25307 14243 25313
rect 2041 25279 2099 25285
rect 2041 25245 2053 25279
rect 2087 25276 2099 25279
rect 2133 25279 2191 25285
rect 2133 25276 2145 25279
rect 2087 25248 2145 25276
rect 2087 25245 2099 25248
rect 2041 25239 2099 25245
rect 2133 25245 2145 25248
rect 2179 25245 2191 25279
rect 2133 25239 2191 25245
rect 12894 25236 12900 25288
rect 12952 25236 12958 25288
rect 13265 25279 13323 25285
rect 13265 25245 13277 25279
rect 13311 25276 13323 25279
rect 13446 25276 13452 25288
rect 13311 25248 13452 25276
rect 13311 25245 13323 25248
rect 13265 25239 13323 25245
rect 13446 25236 13452 25248
rect 13504 25236 13510 25288
rect 13722 25236 13728 25288
rect 13780 25276 13786 25288
rect 14292 25276 14320 25443
rect 14550 25440 14556 25492
rect 14608 25440 14614 25492
rect 20622 25440 20628 25492
rect 20680 25480 20686 25492
rect 20993 25483 21051 25489
rect 20993 25480 21005 25483
rect 20680 25452 21005 25480
rect 20680 25440 20686 25452
rect 20993 25449 21005 25452
rect 21039 25449 21051 25483
rect 20993 25443 21051 25449
rect 26973 25483 27031 25489
rect 26973 25449 26985 25483
rect 27019 25480 27031 25483
rect 27706 25480 27712 25492
rect 27019 25452 27712 25480
rect 27019 25449 27031 25452
rect 26973 25443 27031 25449
rect 17678 25372 17684 25424
rect 17736 25412 17742 25424
rect 18693 25415 18751 25421
rect 18693 25412 18705 25415
rect 17736 25384 18705 25412
rect 17736 25372 17742 25384
rect 18693 25381 18705 25384
rect 18739 25381 18751 25415
rect 18693 25375 18751 25381
rect 15565 25347 15623 25353
rect 15565 25313 15577 25347
rect 15611 25344 15623 25347
rect 16574 25344 16580 25356
rect 15611 25316 16580 25344
rect 15611 25313 15623 25316
rect 15565 25307 15623 25313
rect 16574 25304 16580 25316
rect 16632 25344 16638 25356
rect 18230 25344 18236 25356
rect 16632 25316 18236 25344
rect 16632 25304 16638 25316
rect 18230 25304 18236 25316
rect 18288 25344 18294 25356
rect 19245 25347 19303 25353
rect 19245 25344 19257 25347
rect 18288 25316 19257 25344
rect 18288 25304 18294 25316
rect 19245 25313 19257 25316
rect 19291 25313 19303 25347
rect 19245 25307 19303 25313
rect 23566 25304 23572 25356
rect 23624 25344 23630 25356
rect 23624 25316 26234 25344
rect 23624 25304 23630 25316
rect 13780 25248 14320 25276
rect 13780 25236 13786 25248
rect 14366 25236 14372 25288
rect 14424 25236 14430 25288
rect 14458 25236 14464 25288
rect 14516 25276 14522 25288
rect 14645 25279 14703 25285
rect 14645 25276 14657 25279
rect 14516 25248 14657 25276
rect 14516 25236 14522 25248
rect 14645 25245 14657 25248
rect 14691 25245 14703 25279
rect 14645 25239 14703 25245
rect 14829 25279 14887 25285
rect 14829 25245 14841 25279
rect 14875 25276 14887 25279
rect 15010 25276 15016 25288
rect 14875 25248 15016 25276
rect 14875 25245 14887 25248
rect 14829 25239 14887 25245
rect 15010 25236 15016 25248
rect 15068 25236 15074 25288
rect 16942 25236 16948 25288
rect 17000 25236 17006 25288
rect 17589 25279 17647 25285
rect 17589 25245 17601 25279
rect 17635 25245 17647 25279
rect 17589 25239 17647 25245
rect 13170 25168 13176 25220
rect 13228 25208 13234 25220
rect 14093 25211 14151 25217
rect 14093 25208 14105 25211
rect 13228 25180 14105 25208
rect 13228 25168 13234 25180
rect 14093 25177 14105 25180
rect 14139 25177 14151 25211
rect 14093 25171 14151 25177
rect 15841 25211 15899 25217
rect 15841 25177 15853 25211
rect 15887 25177 15899 25211
rect 17604 25208 17632 25239
rect 17678 25236 17684 25288
rect 17736 25236 17742 25288
rect 17954 25236 17960 25288
rect 18012 25236 18018 25288
rect 18049 25279 18107 25285
rect 18049 25245 18061 25279
rect 18095 25276 18107 25279
rect 18322 25276 18328 25288
rect 18095 25248 18328 25276
rect 18095 25245 18107 25248
rect 18049 25239 18107 25245
rect 18322 25236 18328 25248
rect 18380 25276 18386 25288
rect 18877 25279 18935 25285
rect 18877 25276 18889 25279
rect 18380 25248 18889 25276
rect 18380 25236 18386 25248
rect 18877 25245 18889 25248
rect 18923 25245 18935 25279
rect 18877 25239 18935 25245
rect 19058 25236 19064 25288
rect 19116 25236 19122 25288
rect 17862 25208 17868 25220
rect 17604 25180 17868 25208
rect 15841 25171 15899 25177
rect 934 25100 940 25152
rect 992 25140 998 25152
rect 1857 25143 1915 25149
rect 1857 25140 1869 25143
rect 992 25112 1869 25140
rect 992 25100 998 25112
rect 1857 25109 1869 25112
rect 1903 25109 1915 25143
rect 1857 25103 1915 25109
rect 14734 25100 14740 25152
rect 14792 25100 14798 25152
rect 15856 25140 15884 25171
rect 17862 25168 17868 25180
rect 17920 25208 17926 25220
rect 18417 25211 18475 25217
rect 18417 25208 18429 25211
rect 17920 25180 18429 25208
rect 17920 25168 17926 25180
rect 18417 25177 18429 25180
rect 18463 25177 18475 25211
rect 18417 25171 18475 25177
rect 18969 25211 19027 25217
rect 18969 25177 18981 25211
rect 19015 25208 19027 25211
rect 19521 25211 19579 25217
rect 19521 25208 19533 25211
rect 19015 25180 19533 25208
rect 19015 25177 19027 25180
rect 18969 25171 19027 25177
rect 19521 25177 19533 25180
rect 19567 25177 19579 25211
rect 26206 25208 26234 25316
rect 27080 25285 27108 25452
rect 27706 25440 27712 25452
rect 27764 25480 27770 25492
rect 29362 25480 29368 25492
rect 27764 25452 29368 25480
rect 27764 25440 27770 25452
rect 29362 25440 29368 25452
rect 29420 25440 29426 25492
rect 30834 25440 30840 25492
rect 30892 25480 30898 25492
rect 31021 25483 31079 25489
rect 31021 25480 31033 25483
rect 30892 25452 31033 25480
rect 30892 25440 30898 25452
rect 31021 25449 31033 25452
rect 31067 25449 31079 25483
rect 31021 25443 31079 25449
rect 42061 25483 42119 25489
rect 42061 25449 42073 25483
rect 42107 25480 42119 25483
rect 42426 25480 42432 25492
rect 42107 25452 42432 25480
rect 42107 25449 42119 25452
rect 42061 25443 42119 25449
rect 42426 25440 42432 25452
rect 42484 25440 42490 25492
rect 51534 25440 51540 25492
rect 51592 25480 51598 25492
rect 51902 25480 51908 25492
rect 51592 25452 51908 25480
rect 51592 25440 51598 25452
rect 51902 25440 51908 25452
rect 51960 25440 51966 25492
rect 53650 25440 53656 25492
rect 53708 25440 53714 25492
rect 42337 25415 42395 25421
rect 42337 25412 42349 25415
rect 40788 25384 42349 25412
rect 31294 25344 31300 25356
rect 31220 25316 31300 25344
rect 31220 25285 31248 25316
rect 31294 25304 31300 25316
rect 31352 25344 31358 25356
rect 32582 25344 32588 25356
rect 31352 25316 32588 25344
rect 31352 25304 31358 25316
rect 32582 25304 32588 25316
rect 32640 25304 32646 25356
rect 34422 25304 34428 25356
rect 34480 25304 34486 25356
rect 34790 25304 34796 25356
rect 34848 25344 34854 25356
rect 34848 25316 35112 25344
rect 34848 25304 34854 25316
rect 27065 25279 27123 25285
rect 27065 25245 27077 25279
rect 27111 25245 27123 25279
rect 27065 25239 27123 25245
rect 31205 25279 31263 25285
rect 31205 25245 31217 25279
rect 31251 25245 31263 25279
rect 31205 25239 31263 25245
rect 31386 25236 31392 25288
rect 31444 25236 31450 25288
rect 31573 25279 31631 25285
rect 31573 25245 31585 25279
rect 31619 25276 31631 25279
rect 32122 25276 32128 25288
rect 31619 25248 32128 25276
rect 31619 25245 31631 25248
rect 31573 25239 31631 25245
rect 32122 25236 32128 25248
rect 32180 25276 32186 25288
rect 33962 25276 33968 25288
rect 32180 25248 33968 25276
rect 32180 25236 32186 25248
rect 33962 25236 33968 25248
rect 34020 25236 34026 25288
rect 34054 25236 34060 25288
rect 34112 25276 34118 25288
rect 34149 25279 34207 25285
rect 34149 25276 34161 25279
rect 34112 25248 34161 25276
rect 34112 25236 34118 25248
rect 34149 25245 34161 25248
rect 34195 25245 34207 25279
rect 34149 25239 34207 25245
rect 34241 25279 34299 25285
rect 34241 25245 34253 25279
rect 34287 25245 34299 25279
rect 34241 25239 34299 25245
rect 27801 25211 27859 25217
rect 27801 25208 27813 25211
rect 19521 25171 19579 25177
rect 19628 25180 20010 25208
rect 26206 25180 27813 25208
rect 16850 25140 16856 25152
rect 15856 25112 16856 25140
rect 16850 25100 16856 25112
rect 16908 25100 16914 25152
rect 17310 25100 17316 25152
rect 17368 25100 17374 25152
rect 17402 25100 17408 25152
rect 17460 25100 17466 25152
rect 17770 25100 17776 25152
rect 17828 25100 17834 25152
rect 18138 25100 18144 25152
rect 18196 25100 18202 25152
rect 18322 25100 18328 25152
rect 18380 25100 18386 25152
rect 18506 25100 18512 25152
rect 18564 25100 18570 25152
rect 18598 25100 18604 25152
rect 18656 25140 18662 25152
rect 19628 25140 19656 25180
rect 18656 25112 19656 25140
rect 19904 25140 19932 25180
rect 27801 25177 27813 25180
rect 27847 25208 27859 25211
rect 28442 25208 28448 25220
rect 27847 25180 28448 25208
rect 27847 25177 27859 25180
rect 27801 25171 27859 25177
rect 28442 25168 28448 25180
rect 28500 25168 28506 25220
rect 30926 25168 30932 25220
rect 30984 25208 30990 25220
rect 31297 25211 31355 25217
rect 31297 25208 31309 25211
rect 30984 25180 31309 25208
rect 30984 25168 30990 25180
rect 31297 25177 31309 25180
rect 31343 25177 31355 25211
rect 34256 25208 34284 25239
rect 34514 25236 34520 25288
rect 34572 25236 34578 25288
rect 34882 25236 34888 25288
rect 34940 25236 34946 25288
rect 35084 25285 35112 25316
rect 37826 25304 37832 25356
rect 37884 25304 37890 25356
rect 35069 25279 35127 25285
rect 35069 25245 35081 25279
rect 35115 25245 35127 25279
rect 35069 25239 35127 25245
rect 35253 25279 35311 25285
rect 35253 25245 35265 25279
rect 35299 25276 35311 25279
rect 35434 25276 35440 25288
rect 35299 25248 35440 25276
rect 35299 25245 35311 25248
rect 35253 25239 35311 25245
rect 35434 25236 35440 25248
rect 35492 25236 35498 25288
rect 35713 25279 35771 25285
rect 35713 25276 35725 25279
rect 35544 25248 35725 25276
rect 34256 25180 34744 25208
rect 31297 25171 31355 25177
rect 21085 25143 21143 25149
rect 21085 25140 21097 25143
rect 19904 25112 21097 25140
rect 18656 25100 18662 25112
rect 21085 25109 21097 25112
rect 21131 25109 21143 25143
rect 21085 25103 21143 25109
rect 33778 25100 33784 25152
rect 33836 25140 33842 25152
rect 34716 25149 34744 25180
rect 34790 25168 34796 25220
rect 34848 25208 34854 25220
rect 34977 25211 35035 25217
rect 34977 25208 34989 25211
rect 34848 25180 34989 25208
rect 34848 25168 34854 25180
rect 34977 25177 34989 25180
rect 35023 25177 35035 25211
rect 34977 25171 35035 25177
rect 33965 25143 34023 25149
rect 33965 25140 33977 25143
rect 33836 25112 33977 25140
rect 33836 25100 33842 25112
rect 33965 25109 33977 25112
rect 34011 25109 34023 25143
rect 33965 25103 34023 25109
rect 34701 25143 34759 25149
rect 34701 25109 34713 25143
rect 34747 25109 34759 25143
rect 34701 25103 34759 25109
rect 34882 25100 34888 25152
rect 34940 25140 34946 25152
rect 35544 25140 35572 25248
rect 35713 25245 35725 25248
rect 35759 25245 35771 25279
rect 35713 25239 35771 25245
rect 36078 25236 36084 25288
rect 36136 25236 36142 25288
rect 38194 25236 38200 25288
rect 38252 25236 38258 25288
rect 40788 25276 40816 25384
rect 42337 25381 42349 25384
rect 42383 25412 42395 25415
rect 42518 25412 42524 25424
rect 42383 25384 42524 25412
rect 42383 25381 42395 25384
rect 42337 25375 42395 25381
rect 42518 25372 42524 25384
rect 42576 25372 42582 25424
rect 42794 25372 42800 25424
rect 42852 25412 42858 25424
rect 42852 25384 43300 25412
rect 42852 25372 42858 25384
rect 40862 25304 40868 25356
rect 40920 25344 40926 25356
rect 41049 25347 41107 25353
rect 41049 25344 41061 25347
rect 40920 25316 41061 25344
rect 40920 25304 40926 25316
rect 41049 25313 41061 25316
rect 41095 25313 41107 25347
rect 41049 25307 41107 25313
rect 41141 25347 41199 25353
rect 41141 25313 41153 25347
rect 41187 25344 41199 25347
rect 43162 25344 43168 25356
rect 41187 25316 42932 25344
rect 41187 25313 41199 25316
rect 41141 25307 41199 25313
rect 40957 25279 41015 25285
rect 40957 25276 40969 25279
rect 40788 25248 40969 25276
rect 40957 25245 40969 25248
rect 41003 25245 41015 25279
rect 40957 25239 41015 25245
rect 41414 25236 41420 25288
rect 41472 25236 41478 25288
rect 41509 25279 41567 25285
rect 41509 25245 41521 25279
rect 41555 25245 41567 25279
rect 41509 25239 41567 25245
rect 41877 25279 41935 25285
rect 41877 25245 41889 25279
rect 41923 25276 41935 25279
rect 42150 25276 42156 25288
rect 41923 25248 42156 25276
rect 41923 25245 41935 25248
rect 41877 25239 41935 25245
rect 37090 25168 37096 25220
rect 37148 25168 37154 25220
rect 39206 25168 39212 25220
rect 39264 25168 39270 25220
rect 41325 25211 41383 25217
rect 41325 25177 41337 25211
rect 41371 25208 41383 25211
rect 41524 25208 41552 25239
rect 42150 25236 42156 25248
rect 42208 25236 42214 25288
rect 42429 25279 42487 25285
rect 42429 25245 42441 25279
rect 42475 25276 42487 25279
rect 42610 25276 42616 25288
rect 42475 25248 42616 25276
rect 42475 25245 42487 25248
rect 42429 25239 42487 25245
rect 42610 25236 42616 25248
rect 42668 25236 42674 25288
rect 41371 25180 41552 25208
rect 41371 25177 41383 25180
rect 41325 25171 41383 25177
rect 41690 25168 41696 25220
rect 41748 25168 41754 25220
rect 41785 25211 41843 25217
rect 41785 25177 41797 25211
rect 41831 25177 41843 25211
rect 41785 25171 41843 25177
rect 37550 25149 37556 25152
rect 34940 25112 35572 25140
rect 37507 25143 37556 25149
rect 34940 25100 34946 25112
rect 37507 25109 37519 25143
rect 37553 25109 37556 25143
rect 37507 25103 37556 25109
rect 37550 25100 37556 25103
rect 37608 25100 37614 25152
rect 39623 25143 39681 25149
rect 39623 25109 39635 25143
rect 39669 25140 39681 25143
rect 39758 25140 39764 25152
rect 39669 25112 39764 25140
rect 39669 25109 39681 25112
rect 39623 25103 39681 25109
rect 39758 25100 39764 25112
rect 39816 25100 39822 25152
rect 41230 25100 41236 25152
rect 41288 25140 41294 25152
rect 41800 25140 41828 25171
rect 41288 25112 41828 25140
rect 42904 25140 42932 25316
rect 42996 25316 43168 25344
rect 42996 25285 43024 25316
rect 43162 25304 43168 25316
rect 43220 25304 43226 25356
rect 43272 25353 43300 25384
rect 52362 25372 52368 25424
rect 52420 25412 52426 25424
rect 54478 25412 54484 25424
rect 52420 25384 54484 25412
rect 52420 25372 52426 25384
rect 54478 25372 54484 25384
rect 54536 25412 54542 25424
rect 54536 25384 55214 25412
rect 54536 25372 54542 25384
rect 43257 25347 43315 25353
rect 43257 25313 43269 25347
rect 43303 25313 43315 25347
rect 55186 25344 55214 25384
rect 55309 25347 55367 25353
rect 55309 25344 55321 25347
rect 55186 25316 55321 25344
rect 43257 25307 43315 25313
rect 55309 25313 55321 25316
rect 55355 25313 55367 25347
rect 55309 25307 55367 25313
rect 42981 25279 43039 25285
rect 42981 25245 42993 25279
rect 43027 25245 43039 25279
rect 42981 25239 43039 25245
rect 43625 25279 43683 25285
rect 43625 25245 43637 25279
rect 43671 25276 43683 25279
rect 46566 25276 46572 25288
rect 43671 25248 46572 25276
rect 43671 25245 43683 25248
rect 43625 25239 43683 25245
rect 46566 25236 46572 25248
rect 46624 25236 46630 25288
rect 51258 25236 51264 25288
rect 51316 25276 51322 25288
rect 51629 25279 51687 25285
rect 51629 25276 51641 25279
rect 51316 25248 51641 25276
rect 51316 25236 51322 25248
rect 51629 25245 51641 25248
rect 51675 25245 51687 25279
rect 51629 25239 51687 25245
rect 43346 25168 43352 25220
rect 43404 25208 43410 25220
rect 43441 25211 43499 25217
rect 43441 25208 43453 25211
rect 43404 25180 43453 25208
rect 43404 25168 43410 25180
rect 43441 25177 43453 25180
rect 43487 25177 43499 25211
rect 51644 25208 51672 25239
rect 51718 25236 51724 25288
rect 51776 25236 51782 25288
rect 51994 25236 52000 25288
rect 52052 25236 52058 25288
rect 53101 25279 53159 25285
rect 53101 25245 53113 25279
rect 53147 25276 53159 25279
rect 53374 25276 53380 25288
rect 53147 25248 53380 25276
rect 53147 25245 53159 25248
rect 53101 25239 53159 25245
rect 53374 25236 53380 25248
rect 53432 25236 53438 25288
rect 53466 25236 53472 25288
rect 53524 25236 53530 25288
rect 53558 25236 53564 25288
rect 53616 25276 53622 25288
rect 53699 25279 53757 25285
rect 53699 25276 53711 25279
rect 53616 25248 53711 25276
rect 53616 25236 53622 25248
rect 53699 25245 53711 25248
rect 53745 25245 53757 25279
rect 53699 25239 53757 25245
rect 52270 25208 52276 25220
rect 51644 25180 52276 25208
rect 43441 25171 43499 25177
rect 52270 25168 52276 25180
rect 52328 25168 52334 25220
rect 55582 25168 55588 25220
rect 55640 25168 55646 25220
rect 55692 25180 56074 25208
rect 43714 25140 43720 25152
rect 42904 25112 43720 25140
rect 41288 25100 41294 25112
rect 43714 25100 43720 25112
rect 43772 25100 43778 25152
rect 51074 25100 51080 25152
rect 51132 25140 51138 25152
rect 51445 25143 51503 25149
rect 51445 25140 51457 25143
rect 51132 25112 51457 25140
rect 51132 25100 51138 25112
rect 51445 25109 51457 25112
rect 51491 25109 51503 25143
rect 51445 25103 51503 25109
rect 53190 25100 53196 25152
rect 53248 25100 53254 25152
rect 53926 25100 53932 25152
rect 53984 25140 53990 25152
rect 54478 25140 54484 25152
rect 53984 25112 54484 25140
rect 53984 25100 53990 25112
rect 54478 25100 54484 25112
rect 54536 25140 54542 25152
rect 55692 25140 55720 25180
rect 54536 25112 55720 25140
rect 54536 25100 54542 25112
rect 55766 25100 55772 25152
rect 55824 25140 55830 25152
rect 57057 25143 57115 25149
rect 57057 25140 57069 25143
rect 55824 25112 57069 25140
rect 55824 25100 55830 25112
rect 57057 25109 57069 25112
rect 57103 25109 57115 25143
rect 57057 25103 57115 25109
rect 1104 25050 78844 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 66314 25050
rect 66366 24998 66378 25050
rect 66430 24998 66442 25050
rect 66494 24998 66506 25050
rect 66558 24998 66570 25050
rect 66622 24998 78844 25050
rect 1104 24976 78844 24998
rect 12894 24896 12900 24948
rect 12952 24936 12958 24948
rect 13173 24939 13231 24945
rect 13173 24936 13185 24939
rect 12952 24908 13185 24936
rect 12952 24896 12958 24908
rect 13173 24905 13185 24908
rect 13219 24936 13231 24939
rect 13722 24936 13728 24948
rect 13219 24908 13728 24936
rect 13219 24905 13231 24908
rect 13173 24899 13231 24905
rect 13722 24896 13728 24908
rect 13780 24896 13786 24948
rect 14366 24896 14372 24948
rect 14424 24936 14430 24948
rect 14424 24908 15700 24936
rect 14424 24896 14430 24908
rect 12989 24871 13047 24877
rect 12989 24837 13001 24871
rect 13035 24868 13047 24871
rect 13814 24868 13820 24880
rect 13035 24840 13820 24868
rect 13035 24837 13047 24840
rect 12989 24831 13047 24837
rect 13814 24828 13820 24840
rect 13872 24868 13878 24880
rect 15672 24877 15700 24908
rect 17402 24896 17408 24948
rect 17460 24936 17466 24948
rect 17589 24939 17647 24945
rect 17589 24936 17601 24939
rect 17460 24908 17601 24936
rect 17460 24896 17466 24908
rect 17589 24905 17601 24908
rect 17635 24905 17647 24939
rect 17589 24899 17647 24905
rect 17773 24939 17831 24945
rect 17773 24905 17785 24939
rect 17819 24936 17831 24939
rect 17862 24936 17868 24948
rect 17819 24908 17868 24936
rect 17819 24905 17831 24908
rect 17773 24899 17831 24905
rect 17862 24896 17868 24908
rect 17920 24896 17926 24948
rect 18046 24896 18052 24948
rect 18104 24936 18110 24948
rect 18598 24936 18604 24948
rect 18104 24908 18604 24936
rect 18104 24896 18110 24908
rect 18598 24896 18604 24908
rect 18656 24896 18662 24948
rect 20070 24945 20076 24948
rect 20057 24939 20076 24945
rect 20057 24905 20069 24939
rect 20057 24899 20076 24905
rect 20070 24896 20076 24899
rect 20128 24896 20134 24948
rect 30834 24936 30840 24948
rect 29104 24908 30840 24936
rect 15457 24871 15515 24877
rect 13872 24840 15148 24868
rect 13872 24828 13878 24840
rect 15120 24812 15148 24840
rect 15457 24837 15469 24871
rect 15503 24868 15515 24871
rect 15657 24871 15715 24877
rect 15503 24837 15516 24868
rect 15457 24831 15516 24837
rect 15657 24837 15669 24871
rect 15703 24837 15715 24871
rect 15657 24831 15715 24837
rect 20257 24871 20315 24877
rect 20257 24837 20269 24871
rect 20303 24868 20315 24871
rect 20622 24868 20628 24880
rect 20303 24840 20628 24868
rect 20303 24837 20315 24840
rect 20257 24831 20315 24837
rect 2041 24803 2099 24809
rect 2041 24769 2053 24803
rect 2087 24800 2099 24803
rect 2133 24803 2191 24809
rect 2133 24800 2145 24803
rect 2087 24772 2145 24800
rect 2087 24769 2099 24772
rect 2041 24763 2099 24769
rect 2133 24769 2145 24772
rect 2179 24769 2191 24803
rect 10321 24803 10379 24809
rect 10321 24800 10333 24803
rect 9154 24772 10333 24800
rect 2133 24763 2191 24769
rect 10321 24769 10333 24772
rect 10367 24769 10379 24803
rect 10321 24763 10379 24769
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24800 10839 24803
rect 10870 24800 10876 24812
rect 10827 24772 10876 24800
rect 10827 24769 10839 24772
rect 10781 24763 10839 24769
rect 7742 24692 7748 24744
rect 7800 24692 7806 24744
rect 8021 24735 8079 24741
rect 8021 24701 8033 24735
rect 8067 24732 8079 24735
rect 9030 24732 9036 24744
rect 8067 24704 9036 24732
rect 8067 24701 8079 24704
rect 8021 24695 8079 24701
rect 9030 24692 9036 24704
rect 9088 24692 9094 24744
rect 9493 24735 9551 24741
rect 9493 24701 9505 24735
rect 9539 24732 9551 24735
rect 10137 24735 10195 24741
rect 10137 24732 10149 24735
rect 9539 24704 10149 24732
rect 9539 24701 9551 24704
rect 9493 24695 9551 24701
rect 10137 24701 10149 24704
rect 10183 24701 10195 24735
rect 10336 24732 10364 24763
rect 10870 24760 10876 24772
rect 10928 24760 10934 24812
rect 12345 24803 12403 24809
rect 12345 24769 12357 24803
rect 12391 24769 12403 24803
rect 12345 24763 12403 24769
rect 10336 24704 11008 24732
rect 10137 24695 10195 24701
rect 10152 24664 10180 24695
rect 10410 24664 10416 24676
rect 10152 24636 10416 24664
rect 10410 24624 10416 24636
rect 10468 24664 10474 24676
rect 10980 24664 11008 24704
rect 11054 24692 11060 24744
rect 11112 24692 11118 24744
rect 11146 24692 11152 24744
rect 11204 24732 11210 24744
rect 12360 24732 12388 24763
rect 12526 24760 12532 24812
rect 12584 24760 12590 24812
rect 13081 24803 13139 24809
rect 13081 24769 13093 24803
rect 13127 24769 13139 24803
rect 13081 24763 13139 24769
rect 12805 24735 12863 24741
rect 12805 24732 12817 24735
rect 11204 24704 12817 24732
rect 11204 24692 11210 24704
rect 12805 24701 12817 24704
rect 12851 24701 12863 24735
rect 13096 24732 13124 24763
rect 13722 24760 13728 24812
rect 13780 24800 13786 24812
rect 14185 24803 14243 24809
rect 14185 24800 14197 24803
rect 13780 24772 14197 24800
rect 13780 24760 13786 24772
rect 14185 24769 14197 24772
rect 14231 24769 14243 24803
rect 14185 24763 14243 24769
rect 13446 24732 13452 24744
rect 13096 24704 13452 24732
rect 12805 24695 12863 24701
rect 13446 24692 13452 24704
rect 13504 24692 13510 24744
rect 14200 24732 14228 24763
rect 14274 24760 14280 24812
rect 14332 24760 14338 24812
rect 14461 24803 14519 24809
rect 14461 24769 14473 24803
rect 14507 24800 14519 24803
rect 14553 24803 14611 24809
rect 14553 24800 14565 24803
rect 14507 24772 14565 24800
rect 14507 24769 14519 24772
rect 14461 24763 14519 24769
rect 14553 24769 14565 24772
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 15102 24760 15108 24812
rect 15160 24800 15166 24812
rect 15197 24803 15255 24809
rect 15197 24800 15209 24803
rect 15160 24772 15209 24800
rect 15160 24760 15166 24772
rect 15197 24769 15209 24772
rect 15243 24800 15255 24803
rect 15488 24800 15516 24831
rect 20622 24828 20628 24840
rect 20680 24828 20686 24880
rect 29104 24868 29132 24908
rect 30834 24896 30840 24908
rect 30892 24936 30898 24948
rect 31021 24939 31079 24945
rect 31021 24936 31033 24939
rect 30892 24908 31033 24936
rect 30892 24896 30898 24908
rect 31021 24905 31033 24908
rect 31067 24905 31079 24939
rect 31021 24899 31079 24905
rect 34514 24896 34520 24948
rect 34572 24936 34578 24948
rect 35207 24939 35265 24945
rect 35207 24936 35219 24939
rect 34572 24908 35219 24936
rect 34572 24896 34578 24908
rect 35207 24905 35219 24908
rect 35253 24936 35265 24939
rect 35342 24936 35348 24948
rect 35253 24908 35348 24936
rect 35253 24905 35265 24908
rect 35207 24899 35265 24905
rect 35342 24896 35348 24908
rect 35400 24896 35406 24948
rect 36078 24896 36084 24948
rect 36136 24936 36142 24948
rect 36449 24939 36507 24945
rect 36449 24936 36461 24939
rect 36136 24908 36461 24936
rect 36136 24896 36142 24908
rect 36449 24905 36461 24908
rect 36495 24905 36507 24939
rect 37090 24936 37096 24948
rect 36449 24899 36507 24905
rect 36556 24908 37096 24936
rect 29178 24868 29184 24880
rect 29104 24840 29184 24868
rect 29178 24828 29184 24840
rect 29236 24828 29242 24880
rect 36170 24868 36176 24880
rect 34822 24840 36176 24868
rect 15243 24772 15516 24800
rect 15243 24769 15255 24772
rect 15197 24763 15255 24769
rect 16850 24760 16856 24812
rect 16908 24800 16914 24812
rect 16945 24803 17003 24809
rect 16945 24800 16957 24803
rect 16908 24772 16957 24800
rect 16908 24760 16914 24772
rect 16945 24769 16957 24772
rect 16991 24769 17003 24803
rect 16945 24763 17003 24769
rect 17310 24760 17316 24812
rect 17368 24800 17374 24812
rect 17681 24803 17739 24809
rect 17681 24800 17693 24803
rect 17368 24772 17693 24800
rect 17368 24760 17374 24772
rect 17681 24769 17693 24772
rect 17727 24769 17739 24803
rect 17681 24763 17739 24769
rect 17770 24760 17776 24812
rect 17828 24800 17834 24812
rect 18506 24800 18512 24812
rect 17828 24772 18512 24800
rect 17828 24760 17834 24772
rect 18506 24760 18512 24772
rect 18564 24760 18570 24812
rect 28442 24760 28448 24812
rect 28500 24760 28506 24812
rect 30466 24760 30472 24812
rect 30524 24800 30530 24812
rect 30561 24803 30619 24809
rect 30561 24800 30573 24803
rect 30524 24772 30573 24800
rect 30524 24760 30530 24772
rect 30561 24769 30573 24772
rect 30607 24769 30619 24803
rect 30561 24763 30619 24769
rect 30650 24760 30656 24812
rect 30708 24760 30714 24812
rect 30926 24760 30932 24812
rect 30984 24760 30990 24812
rect 33778 24760 33784 24812
rect 33836 24760 33842 24812
rect 17129 24735 17187 24741
rect 14200 24704 15516 24732
rect 11238 24664 11244 24676
rect 10468 24636 10916 24664
rect 10980 24636 11244 24664
rect 10468 24624 10474 24636
rect 934 24556 940 24608
rect 992 24596 998 24608
rect 1857 24599 1915 24605
rect 1857 24596 1869 24599
rect 992 24568 1869 24596
rect 992 24556 998 24568
rect 1857 24565 1869 24568
rect 1903 24565 1915 24599
rect 1857 24559 1915 24565
rect 9582 24556 9588 24608
rect 9640 24556 9646 24608
rect 10888 24605 10916 24636
rect 11238 24624 11244 24636
rect 11296 24624 11302 24676
rect 11333 24667 11391 24673
rect 11333 24633 11345 24667
rect 11379 24664 11391 24667
rect 13170 24664 13176 24676
rect 11379 24636 13176 24664
rect 11379 24633 11391 24636
rect 11333 24627 11391 24633
rect 13170 24624 13176 24636
rect 13228 24624 13234 24676
rect 13357 24667 13415 24673
rect 13357 24633 13369 24667
rect 13403 24664 13415 24667
rect 14366 24664 14372 24676
rect 13403 24636 14372 24664
rect 13403 24633 13415 24636
rect 13357 24627 13415 24633
rect 14366 24624 14372 24636
rect 14424 24624 14430 24676
rect 14458 24624 14464 24676
rect 14516 24624 14522 24676
rect 10873 24599 10931 24605
rect 10873 24565 10885 24599
rect 10919 24565 10931 24599
rect 10873 24559 10931 24565
rect 11882 24556 11888 24608
rect 11940 24596 11946 24608
rect 12529 24599 12587 24605
rect 12529 24596 12541 24599
rect 11940 24568 12541 24596
rect 11940 24556 11946 24568
rect 12529 24565 12541 24568
rect 12575 24565 12587 24599
rect 12529 24559 12587 24565
rect 13630 24556 13636 24608
rect 13688 24596 13694 24608
rect 14093 24599 14151 24605
rect 14093 24596 14105 24599
rect 13688 24568 14105 24596
rect 13688 24556 13694 24568
rect 14093 24565 14105 24568
rect 14139 24565 14151 24599
rect 14093 24559 14151 24565
rect 15010 24556 15016 24608
rect 15068 24596 15074 24608
rect 15488 24605 15516 24704
rect 17129 24701 17141 24735
rect 17175 24701 17187 24735
rect 17129 24695 17187 24701
rect 17221 24735 17279 24741
rect 17221 24701 17233 24735
rect 17267 24732 17279 24735
rect 17862 24732 17868 24744
rect 17267 24704 17868 24732
rect 17267 24701 17279 24704
rect 17221 24695 17279 24701
rect 17144 24664 17172 24695
rect 17862 24692 17868 24704
rect 17920 24692 17926 24744
rect 28813 24735 28871 24741
rect 28813 24701 28825 24735
rect 28859 24732 28871 24735
rect 30377 24735 30435 24741
rect 30377 24732 30389 24735
rect 28859 24704 30389 24732
rect 28859 24701 28871 24704
rect 28813 24695 28871 24701
rect 30377 24701 30389 24704
rect 30423 24701 30435 24735
rect 30377 24695 30435 24701
rect 30837 24735 30895 24741
rect 30837 24701 30849 24735
rect 30883 24732 30895 24735
rect 31110 24732 31116 24744
rect 30883 24704 31116 24732
rect 30883 24701 30895 24704
rect 30837 24695 30895 24701
rect 31110 24692 31116 24704
rect 31168 24692 31174 24744
rect 33410 24692 33416 24744
rect 33468 24732 33474 24744
rect 34882 24732 34888 24744
rect 33468 24704 34888 24732
rect 33468 24692 33474 24704
rect 34882 24692 34888 24704
rect 34940 24692 34946 24744
rect 18138 24664 18144 24676
rect 17144 24636 18144 24664
rect 18138 24624 18144 24636
rect 18196 24624 18202 24676
rect 30239 24667 30297 24673
rect 30239 24633 30251 24667
rect 30285 24664 30297 24667
rect 30926 24664 30932 24676
rect 30285 24636 30932 24664
rect 30285 24633 30297 24636
rect 30239 24627 30297 24633
rect 30926 24624 30932 24636
rect 30984 24624 30990 24676
rect 15289 24599 15347 24605
rect 15289 24596 15301 24599
rect 15068 24568 15301 24596
rect 15068 24556 15074 24568
rect 15289 24565 15301 24568
rect 15335 24565 15347 24599
rect 15289 24559 15347 24565
rect 15473 24599 15531 24605
rect 15473 24565 15485 24599
rect 15519 24565 15531 24599
rect 15473 24559 15531 24565
rect 18322 24556 18328 24608
rect 18380 24596 18386 24608
rect 19242 24596 19248 24608
rect 18380 24568 19248 24596
rect 18380 24556 18386 24568
rect 19242 24556 19248 24568
rect 19300 24596 19306 24608
rect 19889 24599 19947 24605
rect 19889 24596 19901 24599
rect 19300 24568 19901 24596
rect 19300 24556 19306 24568
rect 19889 24565 19901 24568
rect 19935 24565 19947 24599
rect 19889 24559 19947 24565
rect 20073 24599 20131 24605
rect 20073 24565 20085 24599
rect 20119 24596 20131 24599
rect 20714 24596 20720 24608
rect 20119 24568 20720 24596
rect 20119 24565 20131 24568
rect 20073 24559 20131 24565
rect 20714 24556 20720 24568
rect 20772 24556 20778 24608
rect 34146 24556 34152 24608
rect 34204 24596 34210 24608
rect 34992 24596 35020 24840
rect 36170 24828 36176 24840
rect 36228 24868 36234 24880
rect 36556 24868 36584 24908
rect 37090 24896 37096 24908
rect 37148 24896 37154 24948
rect 38194 24896 38200 24948
rect 38252 24896 38258 24948
rect 43070 24896 43076 24948
rect 43128 24936 43134 24948
rect 43441 24939 43499 24945
rect 43441 24936 43453 24939
rect 43128 24908 43453 24936
rect 43128 24896 43134 24908
rect 43441 24905 43453 24908
rect 43487 24905 43499 24939
rect 43441 24899 43499 24905
rect 43533 24939 43591 24945
rect 43533 24905 43545 24939
rect 43579 24936 43591 24939
rect 44069 24939 44127 24945
rect 44069 24936 44081 24939
rect 43579 24908 44081 24936
rect 43579 24905 43591 24908
rect 43533 24899 43591 24905
rect 44069 24905 44081 24908
rect 44115 24936 44127 24939
rect 44358 24936 44364 24948
rect 44115 24908 44364 24936
rect 44115 24905 44127 24908
rect 44069 24899 44127 24905
rect 44358 24896 44364 24908
rect 44416 24896 44422 24948
rect 44729 24939 44787 24945
rect 44729 24905 44741 24939
rect 44775 24936 44787 24939
rect 46382 24936 46388 24948
rect 44775 24908 46388 24936
rect 44775 24905 44787 24908
rect 44729 24899 44787 24905
rect 46382 24896 46388 24908
rect 46440 24896 46446 24948
rect 51353 24939 51411 24945
rect 51353 24905 51365 24939
rect 51399 24936 51411 24939
rect 51718 24936 51724 24948
rect 51399 24908 51724 24936
rect 51399 24905 51411 24908
rect 51353 24899 51411 24905
rect 51718 24896 51724 24908
rect 51776 24896 51782 24948
rect 51905 24939 51963 24945
rect 51905 24905 51917 24939
rect 51951 24936 51963 24939
rect 51994 24936 52000 24948
rect 51951 24908 52000 24936
rect 51951 24905 51963 24908
rect 51905 24899 51963 24905
rect 51994 24896 52000 24908
rect 52052 24896 52058 24948
rect 53558 24936 53564 24948
rect 53116 24908 53564 24936
rect 36228 24840 36584 24868
rect 36648 24840 38424 24868
rect 36228 24828 36234 24840
rect 36648 24812 36676 24840
rect 36630 24760 36636 24812
rect 36688 24760 36694 24812
rect 36725 24803 36783 24809
rect 36725 24769 36737 24803
rect 36771 24769 36783 24803
rect 36725 24763 36783 24769
rect 37001 24803 37059 24809
rect 37001 24769 37013 24803
rect 37047 24800 37059 24803
rect 37550 24800 37556 24812
rect 37047 24772 37556 24800
rect 37047 24769 37059 24772
rect 37001 24763 37059 24769
rect 36740 24732 36768 24763
rect 37550 24760 37556 24772
rect 37608 24760 37614 24812
rect 37642 24760 37648 24812
rect 37700 24800 37706 24812
rect 37737 24803 37795 24809
rect 37737 24800 37749 24803
rect 37700 24772 37749 24800
rect 37700 24760 37706 24772
rect 37737 24769 37749 24772
rect 37783 24769 37795 24803
rect 37737 24763 37795 24769
rect 37829 24803 37887 24809
rect 37829 24769 37841 24803
rect 37875 24769 37887 24803
rect 37829 24763 37887 24769
rect 37274 24732 37280 24744
rect 36740 24704 37280 24732
rect 37274 24692 37280 24704
rect 37332 24692 37338 24744
rect 37182 24624 37188 24676
rect 37240 24664 37246 24676
rect 37844 24664 37872 24763
rect 37918 24760 37924 24812
rect 37976 24760 37982 24812
rect 38396 24809 38424 24840
rect 41690 24828 41696 24880
rect 41748 24868 41754 24880
rect 41877 24871 41935 24877
rect 41877 24868 41889 24871
rect 41748 24840 41889 24868
rect 41748 24828 41754 24840
rect 41877 24837 41889 24840
rect 41923 24837 41935 24871
rect 44269 24871 44327 24877
rect 44269 24868 44281 24871
rect 41877 24831 41935 24837
rect 44192 24840 44281 24868
rect 38381 24803 38439 24809
rect 38381 24769 38393 24803
rect 38427 24769 38439 24803
rect 38381 24763 38439 24769
rect 38473 24803 38531 24809
rect 38473 24769 38485 24803
rect 38519 24769 38531 24803
rect 38473 24763 38531 24769
rect 38488 24732 38516 24763
rect 38746 24760 38752 24812
rect 38804 24800 38810 24812
rect 39758 24800 39764 24812
rect 38804 24772 39764 24800
rect 38804 24760 38810 24772
rect 39758 24760 39764 24772
rect 39816 24760 39822 24812
rect 42061 24803 42119 24809
rect 42061 24769 42073 24803
rect 42107 24769 42119 24803
rect 42061 24763 42119 24769
rect 38120 24704 38516 24732
rect 42076 24732 42104 24763
rect 42610 24760 42616 24812
rect 42668 24800 42674 24812
rect 42705 24803 42763 24809
rect 42705 24800 42717 24803
rect 42668 24772 42717 24800
rect 42668 24760 42674 24772
rect 42705 24769 42717 24772
rect 42751 24769 42763 24803
rect 42705 24763 42763 24769
rect 42794 24760 42800 24812
rect 42852 24760 42858 24812
rect 42886 24760 42892 24812
rect 42944 24760 42950 24812
rect 43073 24803 43131 24809
rect 43073 24769 43085 24803
rect 43119 24800 43131 24803
rect 43162 24800 43168 24812
rect 43119 24772 43168 24800
rect 43119 24769 43131 24772
rect 43073 24763 43131 24769
rect 43162 24760 43168 24772
rect 43220 24760 43226 24812
rect 43625 24803 43683 24809
rect 43625 24769 43637 24803
rect 43671 24800 43683 24803
rect 44082 24800 44088 24812
rect 43671 24772 44088 24800
rect 43671 24769 43683 24772
rect 43625 24763 43683 24769
rect 44082 24760 44088 24772
rect 44140 24760 44146 24812
rect 43898 24732 43904 24744
rect 42076 24704 43904 24732
rect 38120 24673 38148 24704
rect 43898 24692 43904 24704
rect 43956 24692 43962 24744
rect 44192 24732 44220 24840
rect 44269 24837 44281 24840
rect 44315 24837 44327 24871
rect 44269 24831 44327 24837
rect 48406 24828 48412 24880
rect 48464 24828 48470 24880
rect 50890 24828 50896 24880
rect 50948 24868 50954 24880
rect 51077 24871 51135 24877
rect 51077 24868 51089 24871
rect 50948 24840 51089 24868
rect 50948 24828 50954 24840
rect 51077 24837 51089 24840
rect 51123 24868 51135 24871
rect 53116 24868 53144 24908
rect 53558 24896 53564 24908
rect 53616 24936 53622 24948
rect 54754 24936 54760 24948
rect 53616 24908 54760 24936
rect 53616 24896 53622 24908
rect 54754 24896 54760 24908
rect 54812 24896 54818 24948
rect 55582 24896 55588 24948
rect 55640 24936 55646 24948
rect 55677 24939 55735 24945
rect 55677 24936 55689 24939
rect 55640 24908 55689 24936
rect 55640 24896 55646 24908
rect 55677 24905 55689 24908
rect 55723 24905 55735 24939
rect 55677 24899 55735 24905
rect 51123 24840 53144 24868
rect 51123 24837 51135 24840
rect 51077 24831 51135 24837
rect 53190 24828 53196 24880
rect 53248 24868 53254 24880
rect 53285 24871 53343 24877
rect 53285 24868 53297 24871
rect 53248 24840 53297 24868
rect 53248 24828 53254 24840
rect 53285 24837 53297 24840
rect 53331 24837 53343 24871
rect 55766 24868 55772 24880
rect 53285 24831 53343 24837
rect 55324 24840 55772 24868
rect 55324 24812 55352 24840
rect 55766 24828 55772 24840
rect 55824 24828 55830 24880
rect 44450 24760 44456 24812
rect 44508 24800 44514 24812
rect 44637 24803 44695 24809
rect 44637 24800 44649 24803
rect 44508 24772 44649 24800
rect 44508 24760 44514 24772
rect 44637 24769 44649 24772
rect 44683 24769 44695 24803
rect 44637 24763 44695 24769
rect 44818 24760 44824 24812
rect 44876 24800 44882 24812
rect 45005 24803 45063 24809
rect 45005 24800 45017 24803
rect 44876 24772 45017 24800
rect 44876 24760 44882 24772
rect 45005 24769 45017 24772
rect 45051 24769 45063 24803
rect 45005 24763 45063 24769
rect 45189 24803 45247 24809
rect 45189 24769 45201 24803
rect 45235 24800 45247 24803
rect 45278 24800 45284 24812
rect 45235 24772 45284 24800
rect 45235 24769 45247 24772
rect 45189 24763 45247 24769
rect 45278 24760 45284 24772
rect 45336 24760 45342 24812
rect 49418 24760 49424 24812
rect 49476 24800 49482 24812
rect 49476 24772 50752 24800
rect 49476 24760 49482 24772
rect 44100 24704 44220 24732
rect 37240 24636 37872 24664
rect 38105 24667 38163 24673
rect 37240 24624 37246 24636
rect 38105 24633 38117 24667
rect 38151 24633 38163 24667
rect 38105 24627 38163 24633
rect 43346 24624 43352 24676
rect 43404 24664 43410 24676
rect 43809 24667 43867 24673
rect 43809 24664 43821 24667
rect 43404 24636 43821 24664
rect 43404 24624 43410 24636
rect 43809 24633 43821 24636
rect 43855 24664 43867 24667
rect 44100 24664 44128 24704
rect 45462 24692 45468 24744
rect 45520 24732 45526 24744
rect 47673 24735 47731 24741
rect 47673 24732 47685 24735
rect 45520 24704 47685 24732
rect 45520 24692 45526 24704
rect 47673 24701 47685 24704
rect 47719 24701 47731 24735
rect 47673 24695 47731 24701
rect 47949 24735 48007 24741
rect 47949 24701 47961 24735
rect 47995 24732 48007 24735
rect 48406 24732 48412 24744
rect 47995 24704 48412 24732
rect 47995 24701 48007 24704
rect 47949 24695 48007 24701
rect 48406 24692 48412 24704
rect 48464 24692 48470 24744
rect 50065 24735 50123 24741
rect 50065 24732 50077 24735
rect 49436 24704 50077 24732
rect 43855 24636 44128 24664
rect 43855 24633 43867 24636
rect 43809 24627 43867 24633
rect 34204 24568 35020 24596
rect 36909 24599 36967 24605
rect 34204 24556 34210 24568
rect 36909 24565 36921 24599
rect 36955 24596 36967 24599
rect 38657 24599 38715 24605
rect 38657 24596 38669 24599
rect 36955 24568 38669 24596
rect 36955 24565 36967 24568
rect 36909 24559 36967 24565
rect 38657 24565 38669 24568
rect 38703 24596 38715 24599
rect 38930 24596 38936 24608
rect 38703 24568 38936 24596
rect 38703 24565 38715 24568
rect 38657 24559 38715 24565
rect 38930 24556 38936 24568
rect 38988 24556 38994 24608
rect 42150 24556 42156 24608
rect 42208 24596 42214 24608
rect 42429 24599 42487 24605
rect 42429 24596 42441 24599
rect 42208 24568 42441 24596
rect 42208 24556 42214 24568
rect 42429 24565 42441 24568
rect 42475 24565 42487 24599
rect 42429 24559 42487 24565
rect 43257 24599 43315 24605
rect 43257 24565 43269 24599
rect 43303 24596 43315 24599
rect 43438 24596 43444 24608
rect 43303 24568 43444 24596
rect 43303 24565 43315 24568
rect 43257 24559 43315 24565
rect 43438 24556 43444 24568
rect 43496 24556 43502 24608
rect 43714 24556 43720 24608
rect 43772 24596 43778 24608
rect 43901 24599 43959 24605
rect 43901 24596 43913 24599
rect 43772 24568 43913 24596
rect 43772 24556 43778 24568
rect 43901 24565 43913 24568
rect 43947 24565 43959 24599
rect 43901 24559 43959 24565
rect 44082 24556 44088 24608
rect 44140 24556 44146 24608
rect 49142 24556 49148 24608
rect 49200 24596 49206 24608
rect 49436 24605 49464 24704
rect 50065 24701 50077 24704
rect 50111 24701 50123 24735
rect 50724 24732 50752 24772
rect 50798 24760 50804 24812
rect 50856 24760 50862 24812
rect 50985 24803 51043 24809
rect 50985 24769 50997 24803
rect 51031 24769 51043 24803
rect 50985 24763 51043 24769
rect 51169 24803 51227 24809
rect 51169 24769 51181 24803
rect 51215 24800 51227 24803
rect 51350 24800 51356 24812
rect 51215 24772 51356 24800
rect 51215 24769 51227 24772
rect 51169 24763 51227 24769
rect 51000 24732 51028 24763
rect 51350 24760 51356 24772
rect 51408 24800 51414 24812
rect 52086 24800 52092 24812
rect 51408 24772 52092 24800
rect 51408 24760 51414 24772
rect 52086 24760 52092 24772
rect 52144 24760 52150 24812
rect 52362 24760 52368 24812
rect 52420 24800 52426 24812
rect 53009 24803 53067 24809
rect 53009 24800 53021 24803
rect 52420 24772 53021 24800
rect 52420 24760 52426 24772
rect 53009 24769 53021 24772
rect 53055 24769 53067 24803
rect 55125 24803 55183 24809
rect 53009 24763 53067 24769
rect 50724 24704 51028 24732
rect 50065 24695 50123 24701
rect 51000 24664 51028 24704
rect 52546 24692 52552 24744
rect 52604 24692 52610 24744
rect 53374 24692 53380 24744
rect 53432 24732 53438 24744
rect 54404 24732 54432 24786
rect 55125 24769 55137 24803
rect 55171 24800 55183 24803
rect 55306 24800 55312 24812
rect 55171 24772 55312 24800
rect 55171 24769 55183 24772
rect 55125 24763 55183 24769
rect 55306 24760 55312 24772
rect 55364 24760 55370 24812
rect 55398 24760 55404 24812
rect 55456 24760 55462 24812
rect 55493 24803 55551 24809
rect 55493 24769 55505 24803
rect 55539 24769 55551 24803
rect 55493 24763 55551 24769
rect 54478 24732 54484 24744
rect 53432 24704 54340 24732
rect 54404 24704 54484 24732
rect 53432 24692 53438 24704
rect 53006 24664 53012 24676
rect 51000 24636 53012 24664
rect 53006 24624 53012 24636
rect 53064 24624 53070 24676
rect 54312 24664 54340 24704
rect 54478 24692 54484 24704
rect 54536 24692 54542 24744
rect 55033 24735 55091 24741
rect 55033 24701 55045 24735
rect 55079 24732 55091 24735
rect 55508 24732 55536 24763
rect 55079 24704 55536 24732
rect 55079 24701 55091 24704
rect 55033 24695 55091 24701
rect 55048 24664 55076 24695
rect 54312 24636 55076 24664
rect 49421 24599 49479 24605
rect 49421 24596 49433 24599
rect 49200 24568 49433 24596
rect 49200 24556 49206 24568
rect 49421 24565 49433 24568
rect 49467 24565 49479 24599
rect 49421 24559 49479 24565
rect 49510 24556 49516 24608
rect 49568 24556 49574 24608
rect 55214 24556 55220 24608
rect 55272 24556 55278 24608
rect 1104 24506 78844 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 78844 24506
rect 1104 24432 78844 24454
rect 9030 24352 9036 24404
rect 9088 24352 9094 24404
rect 9861 24395 9919 24401
rect 9861 24392 9873 24395
rect 9416 24364 9873 24392
rect 9416 24265 9444 24364
rect 9861 24361 9873 24364
rect 9907 24392 9919 24395
rect 10781 24395 10839 24401
rect 10781 24392 10793 24395
rect 9907 24364 10793 24392
rect 9907 24361 9919 24364
rect 9861 24355 9919 24361
rect 10781 24361 10793 24364
rect 10827 24361 10839 24395
rect 10781 24355 10839 24361
rect 13357 24395 13415 24401
rect 13357 24361 13369 24395
rect 13403 24392 13415 24395
rect 13446 24392 13452 24404
rect 13403 24364 13452 24392
rect 13403 24361 13415 24364
rect 13357 24355 13415 24361
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 13814 24352 13820 24404
rect 13872 24392 13878 24404
rect 14918 24392 14924 24404
rect 13872 24364 14924 24392
rect 13872 24352 13878 24364
rect 14918 24352 14924 24364
rect 14976 24352 14982 24404
rect 15102 24352 15108 24404
rect 15160 24392 15166 24404
rect 16209 24395 16267 24401
rect 16209 24392 16221 24395
rect 15160 24364 16221 24392
rect 15160 24352 15166 24364
rect 16209 24361 16221 24364
rect 16255 24361 16267 24395
rect 16209 24355 16267 24361
rect 30650 24352 30656 24404
rect 30708 24392 30714 24404
rect 31113 24395 31171 24401
rect 31113 24392 31125 24395
rect 30708 24364 31125 24392
rect 30708 24352 30714 24364
rect 31113 24361 31125 24364
rect 31159 24361 31171 24395
rect 31113 24355 31171 24361
rect 39666 24352 39672 24404
rect 39724 24392 39730 24404
rect 43070 24392 43076 24404
rect 39724 24364 43076 24392
rect 39724 24352 39730 24364
rect 43070 24352 43076 24364
rect 43128 24352 43134 24404
rect 43898 24352 43904 24404
rect 43956 24352 43962 24404
rect 48406 24352 48412 24404
rect 48464 24352 48470 24404
rect 49418 24352 49424 24404
rect 49476 24392 49482 24404
rect 49789 24395 49847 24401
rect 49789 24392 49801 24395
rect 49476 24364 49801 24392
rect 49476 24352 49482 24364
rect 49789 24361 49801 24364
rect 49835 24361 49847 24395
rect 53282 24392 53288 24404
rect 49789 24355 49847 24361
rect 49896 24364 53288 24392
rect 10137 24327 10195 24333
rect 10137 24293 10149 24327
rect 10183 24324 10195 24327
rect 11330 24324 11336 24336
rect 10183 24296 11336 24324
rect 10183 24293 10195 24296
rect 10137 24287 10195 24293
rect 11330 24284 11336 24296
rect 11388 24284 11394 24336
rect 34790 24284 34796 24336
rect 34848 24324 34854 24336
rect 37826 24324 37832 24336
rect 34848 24296 37832 24324
rect 34848 24284 34854 24296
rect 37826 24284 37832 24296
rect 37884 24284 37890 24336
rect 38194 24284 38200 24336
rect 38252 24324 38258 24336
rect 42058 24324 42064 24336
rect 38252 24296 42064 24324
rect 38252 24284 38258 24296
rect 42058 24284 42064 24296
rect 42116 24284 42122 24336
rect 42610 24324 42616 24336
rect 42536 24296 42616 24324
rect 9401 24259 9459 24265
rect 9401 24225 9413 24259
rect 9447 24225 9459 24259
rect 11054 24256 11060 24268
rect 9401 24219 9459 24225
rect 10796 24228 11060 24256
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 9582 24188 9588 24200
rect 9355 24160 9588 24188
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 10594 24188 10600 24200
rect 9968 24160 10600 24188
rect 9845 24123 9903 24129
rect 9845 24089 9857 24123
rect 9891 24120 9903 24123
rect 9968 24120 9996 24160
rect 10594 24148 10600 24160
rect 10652 24148 10658 24200
rect 10796 24197 10824 24228
rect 11054 24216 11060 24228
rect 11112 24216 11118 24268
rect 11882 24216 11888 24268
rect 11940 24216 11946 24268
rect 12526 24216 12532 24268
rect 12584 24256 12590 24268
rect 13541 24259 13599 24265
rect 13541 24256 13553 24259
rect 12584 24228 13553 24256
rect 12584 24216 12590 24228
rect 13541 24225 13553 24228
rect 13587 24225 13599 24259
rect 13541 24219 13599 24225
rect 14734 24216 14740 24268
rect 14792 24216 14798 24268
rect 31386 24216 31392 24268
rect 31444 24256 31450 24268
rect 31444 24228 31524 24256
rect 31444 24216 31450 24228
rect 10689 24191 10747 24197
rect 10689 24157 10701 24191
rect 10735 24188 10747 24191
rect 10781 24191 10839 24197
rect 10781 24188 10793 24191
rect 10735 24160 10793 24188
rect 10735 24157 10747 24160
rect 10689 24151 10747 24157
rect 10781 24157 10793 24160
rect 10827 24157 10839 24191
rect 10781 24151 10839 24157
rect 10870 24148 10876 24200
rect 10928 24148 10934 24200
rect 10962 24148 10968 24200
rect 11020 24188 11026 24200
rect 11609 24191 11667 24197
rect 11609 24188 11621 24191
rect 11020 24160 11621 24188
rect 11020 24148 11026 24160
rect 11609 24157 11621 24160
rect 11655 24157 11667 24191
rect 11609 24151 11667 24157
rect 13449 24191 13507 24197
rect 13449 24157 13461 24191
rect 13495 24157 13507 24191
rect 13449 24151 13507 24157
rect 9891 24092 9996 24120
rect 9891 24089 9903 24092
rect 9845 24083 9903 24089
rect 10042 24080 10048 24132
rect 10100 24080 10106 24132
rect 10410 24080 10416 24132
rect 10468 24080 10474 24132
rect 10505 24123 10563 24129
rect 10505 24089 10517 24123
rect 10551 24120 10563 24123
rect 10888 24120 10916 24148
rect 10551 24092 10916 24120
rect 11057 24123 11115 24129
rect 10551 24089 10563 24092
rect 10505 24083 10563 24089
rect 11057 24089 11069 24123
rect 11103 24120 11115 24123
rect 11146 24120 11152 24132
rect 11103 24092 11152 24120
rect 11103 24089 11115 24092
rect 11057 24083 11115 24089
rect 2038 24012 2044 24064
rect 2096 24012 2102 24064
rect 9030 24012 9036 24064
rect 9088 24052 9094 24064
rect 9677 24055 9735 24061
rect 9677 24052 9689 24055
rect 9088 24024 9689 24052
rect 9088 24012 9094 24024
rect 9677 24021 9689 24024
rect 9723 24021 9735 24055
rect 9677 24015 9735 24021
rect 10321 24055 10379 24061
rect 10321 24021 10333 24055
rect 10367 24052 10379 24055
rect 11072 24052 11100 24083
rect 11146 24080 11152 24092
rect 11204 24080 11210 24132
rect 11238 24080 11244 24132
rect 11296 24120 11302 24132
rect 13464 24120 13492 24151
rect 13630 24148 13636 24200
rect 13688 24148 13694 24200
rect 14366 24148 14372 24200
rect 14424 24188 14430 24200
rect 14461 24191 14519 24197
rect 14461 24188 14473 24191
rect 14424 24160 14473 24188
rect 14424 24148 14430 24160
rect 14461 24157 14473 24160
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 17218 24148 17224 24200
rect 17276 24188 17282 24200
rect 17405 24191 17463 24197
rect 17405 24188 17417 24191
rect 17276 24160 17417 24188
rect 17276 24148 17282 24160
rect 17405 24157 17417 24160
rect 17451 24157 17463 24191
rect 17405 24151 17463 24157
rect 17494 24148 17500 24200
rect 17552 24188 17558 24200
rect 17589 24191 17647 24197
rect 17589 24188 17601 24191
rect 17552 24160 17601 24188
rect 17552 24148 17558 24160
rect 17589 24157 17601 24160
rect 17635 24157 17647 24191
rect 17589 24151 17647 24157
rect 18506 24148 18512 24200
rect 18564 24188 18570 24200
rect 21082 24188 21088 24200
rect 18564 24160 21088 24188
rect 18564 24148 18570 24160
rect 21082 24148 21088 24160
rect 21140 24148 21146 24200
rect 31294 24148 31300 24200
rect 31352 24148 31358 24200
rect 31496 24197 31524 24228
rect 37090 24216 37096 24268
rect 37148 24256 37154 24268
rect 37148 24228 42472 24256
rect 37148 24216 37154 24228
rect 31481 24191 31539 24197
rect 31481 24157 31493 24191
rect 31527 24157 31539 24191
rect 31481 24151 31539 24157
rect 31570 24148 31576 24200
rect 31628 24188 31634 24200
rect 31665 24191 31723 24197
rect 31665 24188 31677 24191
rect 31628 24160 31677 24188
rect 31628 24148 31634 24160
rect 31665 24157 31677 24160
rect 31711 24157 31723 24191
rect 31665 24151 31723 24157
rect 33321 24191 33379 24197
rect 33321 24157 33333 24191
rect 33367 24188 33379 24191
rect 34333 24191 34391 24197
rect 34333 24188 34345 24191
rect 33367 24160 34345 24188
rect 33367 24157 33379 24160
rect 33321 24151 33379 24157
rect 34333 24157 34345 24160
rect 34379 24188 34391 24191
rect 38838 24188 38844 24200
rect 34379 24160 38844 24188
rect 34379 24157 34391 24160
rect 34333 24151 34391 24157
rect 38838 24148 38844 24160
rect 38896 24188 38902 24200
rect 42242 24188 42248 24200
rect 38896 24160 42248 24188
rect 38896 24148 38902 24160
rect 42242 24148 42248 24160
rect 42300 24148 42306 24200
rect 15010 24120 15016 24132
rect 11296 24092 12374 24120
rect 13464 24092 15016 24120
rect 11296 24080 11302 24092
rect 10367 24024 11100 24052
rect 12268 24052 12296 24092
rect 15010 24080 15016 24092
rect 15068 24080 15074 24132
rect 31389 24123 31447 24129
rect 15962 24092 16068 24120
rect 13814 24052 13820 24064
rect 12268 24024 13820 24052
rect 10367 24021 10379 24024
rect 10321 24015 10379 24021
rect 13814 24012 13820 24024
rect 13872 24012 13878 24064
rect 14918 24012 14924 24064
rect 14976 24052 14982 24064
rect 16040 24052 16068 24092
rect 31389 24089 31401 24123
rect 31435 24089 31447 24123
rect 31389 24083 31447 24089
rect 16301 24055 16359 24061
rect 16301 24052 16313 24055
rect 14976 24024 16313 24052
rect 14976 24012 14982 24024
rect 16301 24021 16313 24024
rect 16347 24021 16359 24055
rect 16301 24015 16359 24021
rect 17497 24055 17555 24061
rect 17497 24021 17509 24055
rect 17543 24052 17555 24055
rect 17586 24052 17592 24064
rect 17543 24024 17592 24052
rect 17543 24021 17555 24024
rect 17497 24015 17555 24021
rect 17586 24012 17592 24024
rect 17644 24012 17650 24064
rect 19518 24012 19524 24064
rect 19576 24052 19582 24064
rect 20441 24055 20499 24061
rect 20441 24052 20453 24055
rect 19576 24024 20453 24052
rect 19576 24012 19582 24024
rect 20441 24021 20453 24024
rect 20487 24021 20499 24055
rect 20441 24015 20499 24021
rect 31294 24012 31300 24064
rect 31352 24052 31358 24064
rect 31404 24052 31432 24083
rect 32766 24080 32772 24132
rect 32824 24120 32830 24132
rect 33410 24120 33416 24132
rect 32824 24092 33416 24120
rect 32824 24080 32830 24092
rect 33410 24080 33416 24092
rect 33468 24120 33474 24132
rect 34057 24123 34115 24129
rect 34057 24120 34069 24123
rect 33468 24092 34069 24120
rect 33468 24080 33474 24092
rect 34057 24089 34069 24092
rect 34103 24089 34115 24123
rect 34057 24083 34115 24089
rect 35986 24080 35992 24132
rect 36044 24120 36050 24132
rect 36081 24123 36139 24129
rect 36081 24120 36093 24123
rect 36044 24092 36093 24120
rect 36044 24080 36050 24092
rect 36081 24089 36093 24092
rect 36127 24120 36139 24123
rect 37458 24120 37464 24132
rect 36127 24092 37464 24120
rect 36127 24089 36139 24092
rect 36081 24083 36139 24089
rect 37458 24080 37464 24092
rect 37516 24080 37522 24132
rect 40034 24080 40040 24132
rect 40092 24080 40098 24132
rect 40221 24123 40279 24129
rect 40221 24089 40233 24123
rect 40267 24089 40279 24123
rect 40221 24083 40279 24089
rect 31352 24024 31432 24052
rect 31352 24012 31358 24024
rect 35434 24012 35440 24064
rect 35492 24052 35498 24064
rect 36265 24055 36323 24061
rect 36265 24052 36277 24055
rect 35492 24024 36277 24052
rect 35492 24012 35498 24024
rect 36265 24021 36277 24024
rect 36311 24052 36323 24055
rect 36446 24052 36452 24064
rect 36311 24024 36452 24052
rect 36311 24021 36323 24024
rect 36265 24015 36323 24021
rect 36446 24012 36452 24024
rect 36504 24012 36510 24064
rect 36906 24012 36912 24064
rect 36964 24052 36970 24064
rect 38194 24052 38200 24064
rect 36964 24024 38200 24052
rect 36964 24012 36970 24024
rect 38194 24012 38200 24024
rect 38252 24012 38258 24064
rect 39114 24012 39120 24064
rect 39172 24052 39178 24064
rect 39853 24055 39911 24061
rect 39853 24052 39865 24055
rect 39172 24024 39865 24052
rect 39172 24012 39178 24024
rect 39853 24021 39865 24024
rect 39899 24021 39911 24055
rect 40236 24052 40264 24083
rect 40402 24052 40408 24064
rect 40236 24024 40408 24052
rect 39853 24015 39911 24021
rect 40402 24012 40408 24024
rect 40460 24012 40466 24064
rect 42334 24012 42340 24064
rect 42392 24012 42398 24064
rect 42444 24052 42472 24228
rect 42536 24129 42564 24296
rect 42610 24284 42616 24296
rect 42668 24324 42674 24336
rect 45278 24324 45284 24336
rect 42668 24296 45284 24324
rect 42668 24284 42674 24296
rect 45278 24284 45284 24296
rect 45336 24324 45342 24336
rect 48317 24327 48375 24333
rect 45336 24296 45600 24324
rect 45336 24284 45342 24296
rect 43254 24216 43260 24268
rect 43312 24256 43318 24268
rect 45462 24256 45468 24268
rect 43312 24228 45468 24256
rect 43312 24216 43318 24228
rect 45462 24216 45468 24228
rect 45520 24216 45526 24268
rect 45572 24256 45600 24296
rect 48317 24293 48329 24327
rect 48363 24324 48375 24327
rect 49896 24324 49924 24364
rect 53282 24352 53288 24364
rect 53340 24352 53346 24404
rect 53377 24395 53435 24401
rect 53377 24361 53389 24395
rect 53423 24392 53435 24395
rect 53466 24392 53472 24404
rect 53423 24364 53472 24392
rect 53423 24361 53435 24364
rect 53377 24355 53435 24361
rect 53466 24352 53472 24364
rect 53524 24352 53530 24404
rect 55398 24352 55404 24404
rect 55456 24392 55462 24404
rect 55861 24395 55919 24401
rect 55861 24392 55873 24395
rect 55456 24364 55873 24392
rect 55456 24352 55462 24364
rect 55861 24361 55873 24364
rect 55907 24361 55919 24395
rect 55861 24355 55919 24361
rect 48363 24296 49924 24324
rect 48363 24293 48375 24296
rect 48317 24287 48375 24293
rect 47489 24259 47547 24265
rect 47489 24256 47501 24259
rect 45572 24228 47501 24256
rect 47489 24225 47501 24228
rect 47535 24225 47547 24259
rect 47489 24219 47547 24225
rect 48424 24200 48452 24296
rect 52086 24284 52092 24336
rect 52144 24324 52150 24336
rect 52144 24296 53236 24324
rect 52144 24284 52150 24296
rect 48498 24216 48504 24268
rect 48556 24256 48562 24268
rect 48869 24259 48927 24265
rect 48869 24256 48881 24259
rect 48556 24228 48881 24256
rect 48556 24216 48562 24228
rect 48869 24225 48881 24228
rect 48915 24225 48927 24259
rect 49510 24256 49516 24268
rect 48869 24219 48927 24225
rect 48976 24228 49516 24256
rect 42702 24148 42708 24200
rect 42760 24148 42766 24200
rect 43809 24191 43867 24197
rect 43809 24157 43821 24191
rect 43855 24157 43867 24191
rect 43809 24151 43867 24157
rect 43993 24191 44051 24197
rect 43993 24157 44005 24191
rect 44039 24188 44051 24191
rect 44269 24191 44327 24197
rect 44269 24188 44281 24191
rect 44039 24160 44281 24188
rect 44039 24157 44051 24160
rect 43993 24151 44051 24157
rect 44269 24157 44281 24160
rect 44315 24188 44327 24191
rect 44358 24188 44364 24200
rect 44315 24160 44364 24188
rect 44315 24157 44327 24160
rect 44269 24151 44327 24157
rect 42521 24123 42579 24129
rect 42521 24089 42533 24123
rect 42567 24089 42579 24123
rect 43824 24120 43852 24151
rect 44358 24148 44364 24160
rect 44416 24148 44422 24200
rect 44453 24191 44511 24197
rect 44453 24157 44465 24191
rect 44499 24157 44511 24191
rect 44453 24151 44511 24157
rect 44174 24120 44180 24132
rect 43824 24092 44180 24120
rect 42521 24083 42579 24089
rect 44174 24080 44180 24092
rect 44232 24120 44238 24132
rect 44468 24120 44496 24151
rect 48406 24148 48412 24200
rect 48464 24188 48470 24200
rect 48976 24197 49004 24228
rect 49510 24216 49516 24228
rect 49568 24216 49574 24268
rect 50801 24259 50859 24265
rect 50801 24225 50813 24259
rect 50847 24256 50859 24259
rect 52362 24256 52368 24268
rect 50847 24228 52368 24256
rect 50847 24225 50859 24228
rect 50801 24219 50859 24225
rect 52362 24216 52368 24228
rect 52420 24216 52426 24268
rect 48593 24191 48651 24197
rect 48593 24188 48605 24191
rect 48464 24160 48605 24188
rect 48464 24148 48470 24160
rect 48593 24157 48605 24160
rect 48639 24157 48651 24191
rect 48593 24151 48651 24157
rect 48685 24191 48743 24197
rect 48685 24157 48697 24191
rect 48731 24157 48743 24191
rect 48685 24151 48743 24157
rect 48961 24191 49019 24197
rect 48961 24157 48973 24191
rect 49007 24157 49019 24191
rect 48961 24151 49019 24157
rect 44232 24092 44496 24120
rect 44232 24080 44238 24092
rect 45738 24080 45744 24132
rect 45796 24080 45802 24132
rect 46966 24092 48636 24120
rect 48608 24064 48636 24092
rect 42886 24052 42892 24064
rect 42444 24024 42892 24052
rect 42886 24012 42892 24024
rect 42944 24012 42950 24064
rect 44085 24055 44143 24061
rect 44085 24021 44097 24055
rect 44131 24052 44143 24055
rect 44358 24052 44364 24064
rect 44131 24024 44364 24052
rect 44131 24021 44143 24024
rect 44085 24015 44143 24021
rect 44358 24012 44364 24024
rect 44416 24012 44422 24064
rect 48590 24012 48596 24064
rect 48648 24012 48654 24064
rect 48700 24052 48728 24151
rect 49234 24148 49240 24200
rect 49292 24148 49298 24200
rect 49418 24148 49424 24200
rect 49476 24148 49482 24200
rect 49602 24148 49608 24200
rect 49660 24148 49666 24200
rect 49973 24191 50031 24197
rect 49973 24157 49985 24191
rect 50019 24188 50031 24191
rect 50062 24188 50068 24200
rect 50019 24160 50068 24188
rect 50019 24157 50031 24160
rect 49973 24151 50031 24157
rect 50062 24148 50068 24160
rect 50120 24148 50126 24200
rect 52825 24191 52883 24197
rect 52825 24188 52837 24191
rect 52564 24160 52837 24188
rect 48774 24080 48780 24132
rect 48832 24120 48838 24132
rect 49329 24123 49387 24129
rect 48832 24092 49188 24120
rect 48832 24080 48838 24092
rect 49053 24055 49111 24061
rect 49053 24052 49065 24055
rect 48700 24024 49065 24052
rect 49053 24021 49065 24024
rect 49099 24021 49111 24055
rect 49160 24052 49188 24092
rect 49329 24089 49341 24123
rect 49375 24120 49387 24123
rect 49878 24120 49884 24132
rect 49375 24092 49884 24120
rect 49375 24089 49387 24092
rect 49329 24083 49387 24089
rect 49878 24080 49884 24092
rect 49936 24080 49942 24132
rect 51074 24080 51080 24132
rect 51132 24080 51138 24132
rect 51184 24092 51566 24120
rect 51184 24052 51212 24092
rect 52564 24064 52592 24160
rect 52825 24157 52837 24160
rect 52871 24157 52883 24191
rect 52825 24151 52883 24157
rect 52914 24148 52920 24200
rect 52972 24188 52978 24200
rect 53208 24197 53236 24296
rect 54938 24216 54944 24268
rect 54996 24256 55002 24268
rect 54996 24228 55720 24256
rect 54996 24216 55002 24228
rect 53101 24191 53159 24197
rect 53101 24188 53113 24191
rect 52972 24160 53113 24188
rect 52972 24148 52978 24160
rect 53101 24157 53113 24160
rect 53147 24157 53159 24191
rect 53101 24151 53159 24157
rect 53193 24191 53251 24197
rect 53193 24157 53205 24191
rect 53239 24157 53251 24191
rect 53193 24151 53251 24157
rect 53006 24080 53012 24132
rect 53064 24080 53070 24132
rect 53208 24120 53236 24151
rect 54754 24148 54760 24200
rect 54812 24188 54818 24200
rect 55692 24197 55720 24228
rect 55309 24191 55367 24197
rect 55309 24188 55321 24191
rect 54812 24160 55321 24188
rect 54812 24148 54818 24160
rect 55309 24157 55321 24160
rect 55355 24157 55367 24191
rect 55309 24151 55367 24157
rect 55677 24191 55735 24197
rect 55677 24157 55689 24191
rect 55723 24157 55735 24191
rect 55677 24151 55735 24157
rect 54938 24120 54944 24132
rect 53208 24092 54944 24120
rect 54938 24080 54944 24092
rect 54996 24080 55002 24132
rect 55493 24123 55551 24129
rect 55493 24120 55505 24123
rect 55186 24092 55505 24120
rect 49160 24024 51212 24052
rect 49053 24015 49111 24021
rect 52546 24012 52552 24064
rect 52604 24012 52610 24064
rect 53024 24052 53052 24080
rect 53742 24052 53748 24064
rect 53024 24024 53748 24052
rect 53742 24012 53748 24024
rect 53800 24052 53806 24064
rect 55186 24052 55214 24092
rect 55493 24089 55505 24092
rect 55539 24089 55551 24123
rect 55493 24083 55551 24089
rect 55582 24080 55588 24132
rect 55640 24080 55646 24132
rect 53800 24024 55214 24052
rect 53800 24012 53806 24024
rect 1104 23962 78844 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 66314 23962
rect 66366 23910 66378 23962
rect 66430 23910 66442 23962
rect 66494 23910 66506 23962
rect 66558 23910 66570 23962
rect 66622 23910 78844 23962
rect 1104 23888 78844 23910
rect 1302 23808 1308 23860
rect 1360 23848 1366 23860
rect 1857 23851 1915 23857
rect 1857 23848 1869 23851
rect 1360 23820 1869 23848
rect 1360 23808 1366 23820
rect 1857 23817 1869 23820
rect 1903 23817 1915 23851
rect 9674 23848 9680 23860
rect 1857 23811 1915 23817
rect 8772 23820 9680 23848
rect 2038 23672 2044 23724
rect 2096 23672 2102 23724
rect 7742 23672 7748 23724
rect 7800 23712 7806 23724
rect 8772 23721 8800 23820
rect 9674 23808 9680 23820
rect 9732 23848 9738 23860
rect 10962 23848 10968 23860
rect 9732 23820 10968 23848
rect 9732 23808 9738 23820
rect 10962 23808 10968 23820
rect 11020 23808 11026 23860
rect 14093 23851 14151 23857
rect 14093 23817 14105 23851
rect 14139 23848 14151 23851
rect 14274 23848 14280 23860
rect 14139 23820 14280 23848
rect 14139 23817 14151 23820
rect 14093 23811 14151 23817
rect 14274 23808 14280 23820
rect 14332 23808 14338 23860
rect 17678 23848 17684 23860
rect 17236 23820 17684 23848
rect 9030 23740 9036 23792
rect 9088 23740 9094 23792
rect 10318 23780 10324 23792
rect 10258 23752 10324 23780
rect 10318 23740 10324 23752
rect 10376 23740 10382 23792
rect 10594 23740 10600 23792
rect 10652 23740 10658 23792
rect 17236 23789 17264 23820
rect 17678 23808 17684 23820
rect 17736 23848 17742 23860
rect 19061 23851 19119 23857
rect 19061 23848 19073 23851
rect 17736 23820 19073 23848
rect 17736 23808 17742 23820
rect 19061 23817 19073 23820
rect 19107 23817 19119 23851
rect 19061 23811 19119 23817
rect 21082 23808 21088 23860
rect 21140 23848 21146 23860
rect 21545 23851 21603 23857
rect 21545 23848 21557 23851
rect 21140 23820 21557 23848
rect 21140 23808 21146 23820
rect 21545 23817 21557 23820
rect 21591 23817 21603 23851
rect 22830 23848 22836 23860
rect 21545 23811 21603 23817
rect 22066 23820 22836 23848
rect 17221 23783 17279 23789
rect 17221 23749 17233 23783
rect 17267 23749 17279 23783
rect 17221 23743 17279 23749
rect 17586 23740 17592 23792
rect 17644 23740 17650 23792
rect 18046 23740 18052 23792
rect 18104 23740 18110 23792
rect 20073 23783 20131 23789
rect 20073 23780 20085 23783
rect 19720 23752 20085 23780
rect 8757 23715 8815 23721
rect 8757 23712 8769 23715
rect 7800 23684 8769 23712
rect 7800 23672 7806 23684
rect 8757 23681 8769 23684
rect 8803 23681 8815 23715
rect 10781 23715 10839 23721
rect 10781 23712 10793 23715
rect 8757 23675 8815 23681
rect 10520 23684 10793 23712
rect 2130 23604 2136 23656
rect 2188 23604 2194 23656
rect 10520 23653 10548 23684
rect 10781 23681 10793 23684
rect 10827 23712 10839 23715
rect 10870 23712 10876 23724
rect 10827 23684 10876 23712
rect 10827 23681 10839 23684
rect 10781 23675 10839 23681
rect 10870 23672 10876 23684
rect 10928 23672 10934 23724
rect 10965 23715 11023 23721
rect 10965 23681 10977 23715
rect 11011 23681 11023 23715
rect 10965 23675 11023 23681
rect 11057 23715 11115 23721
rect 11057 23681 11069 23715
rect 11103 23712 11115 23715
rect 11146 23712 11152 23724
rect 11103 23684 11152 23712
rect 11103 23681 11115 23684
rect 11057 23675 11115 23681
rect 10505 23647 10563 23653
rect 10505 23613 10517 23647
rect 10551 23613 10563 23647
rect 10980 23644 11008 23675
rect 11146 23672 11152 23684
rect 11204 23672 11210 23724
rect 16942 23672 16948 23724
rect 17000 23672 17006 23724
rect 17034 23672 17040 23724
rect 17092 23672 17098 23724
rect 19337 23715 19395 23721
rect 19337 23681 19349 23715
rect 19383 23712 19395 23715
rect 19518 23712 19524 23724
rect 19383 23684 19524 23712
rect 19383 23681 19395 23684
rect 19337 23675 19395 23681
rect 19518 23672 19524 23684
rect 19576 23672 19582 23724
rect 10980 23616 11100 23644
rect 10505 23607 10563 23613
rect 11072 23588 11100 23616
rect 11054 23536 11060 23588
rect 11112 23536 11118 23588
rect 10870 23468 10876 23520
rect 10928 23508 10934 23520
rect 11164 23508 11192 23672
rect 14458 23604 14464 23656
rect 14516 23644 14522 23656
rect 14645 23647 14703 23653
rect 14645 23644 14657 23647
rect 14516 23616 14657 23644
rect 14516 23604 14522 23616
rect 14645 23613 14657 23616
rect 14691 23613 14703 23647
rect 14645 23607 14703 23613
rect 16666 23604 16672 23656
rect 16724 23644 16730 23656
rect 17313 23647 17371 23653
rect 17313 23644 17325 23647
rect 16724 23616 17325 23644
rect 16724 23604 16730 23616
rect 17313 23613 17325 23616
rect 17359 23613 17371 23647
rect 17313 23607 17371 23613
rect 17218 23536 17224 23588
rect 17276 23536 17282 23588
rect 10928 23480 11192 23508
rect 17328 23508 17356 23607
rect 17586 23604 17592 23656
rect 17644 23644 17650 23656
rect 19242 23644 19248 23656
rect 17644 23616 19248 23644
rect 17644 23604 17650 23616
rect 19242 23604 19248 23616
rect 19300 23644 19306 23656
rect 19720 23653 19748 23752
rect 20073 23749 20085 23752
rect 20119 23749 20131 23783
rect 21821 23783 21879 23789
rect 21821 23780 21833 23783
rect 21298 23752 21833 23780
rect 20073 23743 20131 23749
rect 21821 23749 21833 23752
rect 21867 23780 21879 23783
rect 22066 23780 22094 23820
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 30098 23808 30104 23860
rect 30156 23848 30162 23860
rect 30926 23848 30932 23860
rect 30156 23820 30932 23848
rect 30156 23808 30162 23820
rect 30926 23808 30932 23820
rect 30984 23848 30990 23860
rect 35897 23851 35955 23857
rect 30984 23820 35664 23848
rect 30984 23808 30990 23820
rect 21867 23752 22094 23780
rect 21867 23749 21879 23752
rect 21821 23743 21879 23749
rect 30834 23740 30840 23792
rect 30892 23740 30898 23792
rect 34146 23740 34152 23792
rect 34204 23740 34210 23792
rect 34698 23740 34704 23792
rect 34756 23780 34762 23792
rect 35069 23783 35127 23789
rect 35069 23780 35081 23783
rect 34756 23752 35081 23780
rect 34756 23740 34762 23752
rect 35069 23749 35081 23752
rect 35115 23749 35127 23783
rect 35069 23743 35127 23749
rect 35434 23740 35440 23792
rect 35492 23780 35498 23792
rect 35636 23789 35664 23820
rect 35897 23817 35909 23851
rect 35943 23848 35955 23851
rect 37090 23848 37096 23860
rect 35943 23820 36124 23848
rect 35943 23817 35955 23820
rect 35897 23811 35955 23817
rect 35529 23783 35587 23789
rect 35529 23780 35541 23783
rect 35492 23752 35541 23780
rect 35492 23740 35498 23752
rect 35529 23749 35541 23752
rect 35575 23749 35587 23783
rect 35529 23743 35587 23749
rect 35621 23783 35679 23789
rect 35621 23749 35633 23783
rect 35667 23749 35679 23783
rect 35986 23780 35992 23792
rect 35621 23743 35679 23749
rect 35728 23752 35992 23780
rect 28442 23672 28448 23724
rect 28500 23712 28506 23724
rect 30101 23715 30159 23721
rect 30101 23712 30113 23715
rect 28500 23684 30113 23712
rect 28500 23672 28506 23684
rect 30101 23681 30113 23684
rect 30147 23681 30159 23715
rect 30101 23675 30159 23681
rect 31294 23672 31300 23724
rect 31352 23712 31358 23724
rect 31895 23715 31953 23721
rect 31895 23712 31907 23715
rect 31352 23684 31907 23712
rect 31352 23672 31358 23684
rect 31895 23681 31907 23684
rect 31941 23712 31953 23715
rect 34563 23715 34621 23721
rect 31941 23684 33272 23712
rect 31941 23681 31953 23684
rect 31895 23675 31953 23681
rect 19429 23647 19487 23653
rect 19429 23644 19441 23647
rect 19300 23616 19441 23644
rect 19300 23604 19306 23616
rect 19429 23613 19441 23616
rect 19475 23613 19487 23647
rect 19429 23607 19487 23613
rect 19705 23647 19763 23653
rect 19705 23613 19717 23647
rect 19751 23613 19763 23647
rect 19705 23607 19763 23613
rect 19797 23647 19855 23653
rect 19797 23613 19809 23647
rect 19843 23613 19855 23647
rect 19797 23607 19855 23613
rect 19812 23508 19840 23607
rect 30466 23604 30472 23656
rect 30524 23604 30530 23656
rect 30834 23604 30840 23656
rect 30892 23644 30898 23656
rect 30892 23616 31248 23644
rect 30892 23604 30898 23616
rect 31220 23576 31248 23616
rect 32122 23604 32128 23656
rect 32180 23644 32186 23656
rect 32766 23644 32772 23656
rect 32180 23616 32772 23644
rect 32180 23604 32186 23616
rect 32766 23604 32772 23616
rect 32824 23604 32830 23656
rect 33134 23604 33140 23656
rect 33192 23604 33198 23656
rect 33244 23644 33272 23684
rect 34563 23681 34575 23715
rect 34609 23712 34621 23715
rect 34790 23712 34796 23724
rect 34609 23684 34796 23712
rect 34609 23681 34621 23684
rect 34563 23675 34621 23681
rect 34790 23672 34796 23684
rect 34848 23672 34854 23724
rect 34885 23715 34943 23721
rect 34885 23681 34897 23715
rect 34931 23681 34943 23715
rect 34885 23675 34943 23681
rect 34977 23715 35035 23721
rect 34977 23681 34989 23715
rect 35023 23681 35035 23715
rect 34977 23675 35035 23681
rect 33318 23644 33324 23656
rect 33244 23616 33324 23644
rect 33318 23604 33324 23616
rect 33376 23604 33382 23656
rect 34900 23644 34928 23675
rect 33888 23616 34928 23644
rect 32217 23579 32275 23585
rect 32217 23576 32229 23579
rect 31220 23548 32229 23576
rect 32217 23545 32229 23548
rect 32263 23545 32275 23579
rect 32217 23539 32275 23545
rect 17328 23480 19840 23508
rect 10928 23468 10934 23480
rect 30374 23468 30380 23520
rect 30432 23508 30438 23520
rect 31018 23508 31024 23520
rect 30432 23480 31024 23508
rect 30432 23468 30438 23480
rect 31018 23468 31024 23480
rect 31076 23468 31082 23520
rect 32950 23468 32956 23520
rect 33008 23508 33014 23520
rect 33888 23508 33916 23616
rect 33962 23536 33968 23588
rect 34020 23576 34026 23588
rect 34992 23576 35020 23675
rect 35250 23672 35256 23724
rect 35308 23672 35314 23724
rect 35342 23672 35348 23724
rect 35400 23672 35406 23724
rect 35728 23721 35756 23752
rect 35986 23740 35992 23752
rect 36044 23740 36050 23792
rect 36096 23721 36124 23820
rect 36372 23820 37096 23848
rect 36372 23789 36400 23820
rect 37090 23808 37096 23820
rect 37148 23808 37154 23860
rect 38194 23848 38200 23860
rect 37660 23820 38200 23848
rect 36357 23783 36415 23789
rect 36357 23749 36369 23783
rect 36403 23749 36415 23783
rect 36357 23743 36415 23749
rect 36449 23783 36507 23789
rect 36449 23749 36461 23783
rect 36495 23780 36507 23783
rect 37182 23780 37188 23792
rect 36495 23752 37188 23780
rect 36495 23749 36507 23752
rect 36449 23743 36507 23749
rect 37182 23740 37188 23752
rect 37240 23740 37246 23792
rect 37550 23740 37556 23792
rect 37608 23740 37614 23792
rect 37660 23789 37688 23820
rect 38194 23808 38200 23820
rect 38252 23808 38258 23860
rect 39206 23808 39212 23860
rect 39264 23808 39270 23860
rect 40034 23808 40040 23860
rect 40092 23848 40098 23860
rect 41049 23851 41107 23857
rect 41049 23848 41061 23851
rect 40092 23820 41061 23848
rect 40092 23808 40098 23820
rect 41049 23817 41061 23820
rect 41095 23848 41107 23851
rect 43806 23848 43812 23860
rect 41095 23820 43812 23848
rect 41095 23817 41107 23820
rect 41049 23811 41107 23817
rect 43806 23808 43812 23820
rect 43864 23808 43870 23860
rect 45738 23808 45744 23860
rect 45796 23848 45802 23860
rect 45925 23851 45983 23857
rect 45925 23848 45937 23851
rect 45796 23820 45937 23848
rect 45796 23808 45802 23820
rect 45925 23817 45937 23820
rect 45971 23817 45983 23851
rect 45925 23811 45983 23817
rect 49326 23808 49332 23860
rect 49384 23848 49390 23860
rect 49789 23851 49847 23857
rect 49789 23848 49801 23851
rect 49384 23820 49801 23848
rect 49384 23808 49390 23820
rect 49789 23817 49801 23820
rect 49835 23848 49847 23851
rect 52086 23848 52092 23860
rect 49835 23820 52092 23848
rect 49835 23817 49847 23820
rect 49789 23811 49847 23817
rect 52086 23808 52092 23820
rect 52144 23808 52150 23860
rect 37645 23783 37703 23789
rect 37645 23749 37657 23783
rect 37691 23749 37703 23783
rect 39224 23780 39252 23808
rect 39482 23780 39488 23792
rect 37645 23743 37703 23749
rect 38948 23752 39488 23780
rect 35713 23715 35771 23721
rect 35713 23681 35725 23715
rect 35759 23681 35771 23715
rect 35713 23675 35771 23681
rect 36081 23715 36139 23721
rect 36081 23681 36093 23715
rect 36127 23681 36139 23715
rect 36081 23675 36139 23681
rect 36174 23715 36232 23721
rect 36174 23681 36186 23715
rect 36220 23681 36232 23715
rect 36174 23675 36232 23681
rect 36546 23715 36604 23721
rect 36546 23681 36558 23715
rect 36592 23681 36604 23715
rect 37461 23715 37519 23721
rect 37461 23712 37473 23715
rect 36546 23675 36604 23681
rect 37292 23684 37473 23712
rect 36189 23644 36217 23675
rect 35544 23616 36217 23644
rect 35544 23576 35572 23616
rect 34020 23548 35572 23576
rect 34020 23536 34026 23548
rect 36078 23536 36084 23588
rect 36136 23576 36142 23588
rect 36556 23576 36584 23675
rect 36817 23579 36875 23585
rect 36817 23576 36829 23579
rect 36136 23548 36829 23576
rect 36136 23536 36142 23548
rect 36817 23545 36829 23548
rect 36863 23545 36875 23579
rect 37292 23576 37320 23684
rect 37461 23681 37473 23684
rect 37507 23681 37519 23715
rect 37461 23675 37519 23681
rect 37826 23672 37832 23724
rect 37884 23672 37890 23724
rect 38948 23721 38976 23752
rect 39482 23740 39488 23752
rect 39540 23740 39546 23792
rect 39577 23783 39635 23789
rect 39577 23749 39589 23783
rect 39623 23780 39635 23783
rect 39914 23783 39972 23789
rect 39914 23780 39926 23783
rect 39623 23752 39926 23780
rect 39623 23749 39635 23752
rect 39577 23743 39635 23749
rect 39914 23749 39926 23752
rect 39960 23749 39972 23783
rect 39914 23743 39972 23749
rect 42058 23740 42064 23792
rect 42116 23780 42122 23792
rect 42429 23783 42487 23789
rect 42429 23780 42441 23783
rect 42116 23752 42441 23780
rect 42116 23740 42122 23752
rect 42429 23749 42441 23752
rect 42475 23749 42487 23783
rect 42429 23743 42487 23749
rect 42702 23740 42708 23792
rect 42760 23780 42766 23792
rect 42981 23783 43039 23789
rect 42981 23780 42993 23783
rect 42760 23752 42993 23780
rect 42760 23740 42766 23752
rect 42981 23749 42993 23752
rect 43027 23749 43039 23783
rect 44634 23780 44640 23792
rect 42981 23743 43039 23749
rect 44284 23752 44640 23780
rect 38933 23715 38991 23721
rect 38933 23681 38945 23715
rect 38979 23681 38991 23715
rect 38933 23675 38991 23681
rect 39114 23672 39120 23724
rect 39172 23672 39178 23724
rect 39209 23715 39267 23721
rect 39209 23681 39221 23715
rect 39255 23681 39267 23715
rect 39209 23675 39267 23681
rect 39301 23715 39359 23721
rect 39301 23681 39313 23715
rect 39347 23712 39359 23715
rect 40310 23712 40316 23724
rect 39347 23684 40316 23712
rect 39347 23681 39359 23684
rect 39301 23675 39359 23681
rect 37366 23604 37372 23656
rect 37424 23644 37430 23656
rect 39224 23644 39252 23675
rect 40310 23672 40316 23684
rect 40368 23672 40374 23724
rect 42889 23715 42947 23721
rect 43165 23715 43223 23721
rect 42889 23681 42901 23715
rect 42935 23687 43024 23715
rect 42935 23681 42947 23687
rect 42889 23675 42947 23681
rect 37424 23616 39252 23644
rect 37424 23604 37430 23616
rect 39666 23604 39672 23656
rect 39724 23604 39730 23656
rect 42996 23644 43024 23687
rect 43165 23681 43177 23715
rect 43211 23712 43223 23715
rect 43714 23712 43720 23724
rect 43211 23684 43720 23712
rect 43211 23681 43223 23684
rect 43165 23675 43223 23681
rect 43714 23672 43720 23684
rect 43772 23672 43778 23724
rect 44174 23672 44180 23724
rect 44232 23712 44238 23724
rect 44284 23721 44312 23752
rect 44634 23740 44640 23752
rect 44692 23740 44698 23792
rect 45278 23740 45284 23792
rect 45336 23780 45342 23792
rect 46293 23783 46351 23789
rect 46293 23780 46305 23783
rect 45336 23752 46305 23780
rect 45336 23740 45342 23752
rect 46293 23749 46305 23752
rect 46339 23749 46351 23783
rect 48406 23780 48412 23792
rect 46293 23743 46351 23749
rect 48240 23752 48412 23780
rect 44269 23715 44327 23721
rect 44269 23712 44281 23715
rect 44232 23684 44281 23712
rect 44232 23672 44238 23684
rect 44269 23681 44281 23684
rect 44315 23681 44327 23715
rect 44269 23675 44327 23681
rect 44358 23672 44364 23724
rect 44416 23672 44422 23724
rect 44450 23672 44456 23724
rect 44508 23672 44514 23724
rect 46382 23672 46388 23724
rect 46440 23672 46446 23724
rect 48240 23721 48268 23752
rect 48406 23740 48412 23752
rect 48464 23740 48470 23792
rect 50893 23783 50951 23789
rect 50893 23749 50905 23783
rect 50939 23780 50951 23783
rect 52546 23780 52552 23792
rect 50939 23752 52552 23780
rect 50939 23749 50951 23752
rect 50893 23743 50951 23749
rect 52546 23740 52552 23752
rect 52604 23740 52610 23792
rect 55306 23780 55312 23792
rect 54312 23752 55312 23780
rect 47949 23715 48007 23721
rect 47949 23681 47961 23715
rect 47995 23712 48007 23715
rect 48225 23715 48283 23721
rect 48225 23712 48237 23715
rect 47995 23684 48237 23712
rect 47995 23681 48007 23684
rect 47949 23675 48007 23681
rect 48225 23681 48237 23684
rect 48271 23681 48283 23715
rect 48225 23675 48283 23681
rect 48314 23672 48320 23724
rect 48372 23672 48378 23724
rect 48593 23715 48651 23721
rect 48593 23681 48605 23715
rect 48639 23712 48651 23715
rect 48869 23715 48927 23721
rect 48869 23712 48881 23715
rect 48639 23684 48881 23712
rect 48639 23681 48651 23684
rect 48593 23675 48651 23681
rect 48869 23681 48881 23684
rect 48915 23681 48927 23715
rect 48869 23675 48927 23681
rect 48958 23672 48964 23724
rect 49016 23712 49022 23724
rect 49605 23715 49663 23721
rect 49605 23712 49617 23715
rect 49016 23684 49617 23712
rect 49016 23672 49022 23684
rect 49605 23681 49617 23684
rect 49651 23712 49663 23715
rect 49973 23715 50031 23721
rect 49973 23712 49985 23715
rect 49651 23684 49985 23712
rect 49651 23681 49663 23684
rect 49605 23675 49663 23681
rect 49973 23681 49985 23684
rect 50019 23712 50031 23715
rect 50522 23712 50528 23724
rect 50019 23684 50528 23712
rect 50019 23681 50031 23684
rect 49973 23675 50031 23681
rect 50522 23672 50528 23684
rect 50580 23672 50586 23724
rect 50617 23715 50675 23721
rect 50617 23681 50629 23715
rect 50663 23712 50675 23715
rect 50706 23712 50712 23724
rect 50663 23684 50712 23712
rect 50663 23681 50675 23684
rect 50617 23675 50675 23681
rect 50706 23672 50712 23684
rect 50764 23672 50770 23724
rect 50801 23715 50859 23721
rect 50801 23681 50813 23715
rect 50847 23681 50859 23715
rect 51009 23715 51067 23721
rect 51009 23712 51021 23715
rect 50801 23675 50859 23681
rect 51005 23681 51021 23712
rect 51055 23681 51067 23715
rect 51005 23675 51067 23681
rect 43622 23644 43628 23656
rect 42996 23616 43628 23644
rect 43622 23604 43628 23616
rect 43680 23644 43686 23656
rect 44545 23647 44603 23653
rect 44545 23644 44557 23647
rect 43680 23616 44557 23644
rect 43680 23604 43686 23616
rect 44545 23613 44557 23616
rect 44591 23613 44603 23647
rect 44545 23607 44603 23613
rect 45830 23604 45836 23656
rect 45888 23644 45894 23656
rect 46569 23647 46627 23653
rect 46569 23644 46581 23647
rect 45888 23616 46581 23644
rect 45888 23604 45894 23616
rect 46569 23613 46581 23616
rect 46615 23644 46627 23647
rect 46615 23616 48314 23644
rect 46615 23613 46627 23616
rect 46569 23607 46627 23613
rect 38013 23579 38071 23585
rect 38013 23576 38025 23579
rect 37292 23548 38025 23576
rect 36817 23539 36875 23545
rect 38013 23545 38025 23548
rect 38059 23576 38071 23579
rect 38470 23576 38476 23588
rect 38059 23548 38476 23576
rect 38059 23545 38071 23548
rect 38013 23539 38071 23545
rect 38470 23536 38476 23548
rect 38528 23536 38534 23588
rect 42242 23536 42248 23588
rect 42300 23576 42306 23588
rect 43257 23579 43315 23585
rect 43257 23576 43269 23579
rect 42300 23548 43269 23576
rect 42300 23536 42306 23548
rect 43257 23545 43269 23548
rect 43303 23545 43315 23579
rect 43257 23539 43315 23545
rect 33008 23480 33916 23508
rect 33008 23468 33014 23480
rect 34698 23468 34704 23520
rect 34756 23468 34762 23520
rect 36722 23468 36728 23520
rect 36780 23468 36786 23520
rect 37274 23468 37280 23520
rect 37332 23468 37338 23520
rect 41690 23468 41696 23520
rect 41748 23508 41754 23520
rect 44174 23508 44180 23520
rect 41748 23480 44180 23508
rect 41748 23468 41754 23480
rect 44174 23468 44180 23480
rect 44232 23468 44238 23520
rect 44450 23468 44456 23520
rect 44508 23508 44514 23520
rect 44729 23511 44787 23517
rect 44729 23508 44741 23511
rect 44508 23480 44741 23508
rect 44508 23468 44514 23480
rect 44729 23477 44741 23480
rect 44775 23477 44787 23511
rect 44729 23471 44787 23477
rect 48038 23468 48044 23520
rect 48096 23468 48102 23520
rect 48286 23508 48314 23616
rect 48498 23604 48504 23656
rect 48556 23604 48562 23656
rect 49234 23604 49240 23656
rect 49292 23644 49298 23656
rect 49418 23644 49424 23656
rect 49292 23616 49424 23644
rect 49292 23604 49298 23616
rect 49418 23604 49424 23616
rect 49476 23604 49482 23656
rect 50246 23604 50252 23656
rect 50304 23644 50310 23656
rect 50816 23644 50844 23675
rect 51005 23644 51033 23675
rect 52914 23672 52920 23724
rect 52972 23712 52978 23724
rect 54312 23721 54340 23752
rect 55306 23740 55312 23752
rect 55364 23740 55370 23792
rect 54297 23715 54355 23721
rect 54297 23712 54309 23715
rect 52972 23684 54309 23712
rect 52972 23672 52978 23684
rect 54297 23681 54309 23684
rect 54343 23681 54355 23715
rect 54297 23675 54355 23681
rect 54481 23715 54539 23721
rect 54481 23681 54493 23715
rect 54527 23681 54539 23715
rect 54481 23675 54539 23681
rect 50304 23616 50844 23644
rect 50908 23616 51033 23644
rect 50304 23604 50310 23616
rect 48516 23576 48544 23604
rect 49050 23576 49056 23588
rect 48516 23548 49056 23576
rect 49050 23536 49056 23548
rect 49108 23536 49114 23588
rect 50522 23536 50528 23588
rect 50580 23576 50586 23588
rect 50908 23576 50936 23616
rect 53742 23604 53748 23656
rect 53800 23644 53806 23656
rect 54496 23644 54524 23675
rect 54570 23672 54576 23724
rect 54628 23672 54634 23724
rect 54665 23715 54723 23721
rect 54665 23681 54677 23715
rect 54711 23712 54723 23715
rect 54938 23712 54944 23724
rect 54711 23684 54944 23712
rect 54711 23681 54723 23684
rect 54665 23675 54723 23681
rect 54938 23672 54944 23684
rect 54996 23672 55002 23724
rect 58526 23672 58532 23724
rect 58584 23712 58590 23724
rect 77849 23715 77907 23721
rect 77849 23712 77861 23715
rect 58584 23684 77861 23712
rect 58584 23672 58590 23684
rect 77849 23681 77861 23684
rect 77895 23712 77907 23715
rect 78033 23715 78091 23721
rect 78033 23712 78045 23715
rect 77895 23684 78045 23712
rect 77895 23681 77907 23684
rect 77849 23675 77907 23681
rect 78033 23681 78045 23684
rect 78079 23681 78091 23715
rect 78033 23675 78091 23681
rect 53800 23616 54524 23644
rect 53800 23604 53806 23616
rect 56042 23576 56048 23588
rect 50580 23548 50936 23576
rect 51000 23548 56048 23576
rect 50580 23536 50586 23548
rect 51000 23508 51028 23548
rect 56042 23536 56048 23548
rect 56100 23536 56106 23588
rect 48286 23480 51028 23508
rect 51074 23468 51080 23520
rect 51132 23508 51138 23520
rect 51169 23511 51227 23517
rect 51169 23508 51181 23511
rect 51132 23480 51181 23508
rect 51132 23468 51138 23480
rect 51169 23477 51181 23480
rect 51215 23477 51227 23511
rect 51169 23471 51227 23477
rect 54849 23511 54907 23517
rect 54849 23477 54861 23511
rect 54895 23508 54907 23511
rect 55122 23508 55128 23520
rect 54895 23480 55128 23508
rect 54895 23477 54907 23480
rect 54849 23471 54907 23477
rect 55122 23468 55128 23480
rect 55180 23468 55186 23520
rect 78214 23468 78220 23520
rect 78272 23468 78278 23520
rect 1104 23418 78844 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 78844 23418
rect 1104 23344 78844 23366
rect 17405 23307 17463 23313
rect 17405 23273 17417 23307
rect 17451 23304 17463 23307
rect 17494 23304 17500 23316
rect 17451 23276 17500 23304
rect 17451 23273 17463 23276
rect 17405 23267 17463 23273
rect 17494 23264 17500 23276
rect 17552 23264 17558 23316
rect 17589 23307 17647 23313
rect 17589 23273 17601 23307
rect 17635 23304 17647 23307
rect 17770 23304 17776 23316
rect 17635 23276 17776 23304
rect 17635 23273 17647 23276
rect 17589 23267 17647 23273
rect 1210 23196 1216 23248
rect 1268 23236 1274 23248
rect 2317 23239 2375 23245
rect 2317 23236 2329 23239
rect 1268 23208 2329 23236
rect 1268 23196 1274 23208
rect 2317 23205 2329 23208
rect 2363 23205 2375 23239
rect 2317 23199 2375 23205
rect 17034 23196 17040 23248
rect 17092 23236 17098 23248
rect 17604 23236 17632 23267
rect 17770 23264 17776 23276
rect 17828 23264 17834 23316
rect 18693 23307 18751 23313
rect 18693 23273 18705 23307
rect 18739 23304 18751 23307
rect 19334 23304 19340 23316
rect 18739 23276 19340 23304
rect 18739 23273 18751 23276
rect 18693 23267 18751 23273
rect 17092 23208 17632 23236
rect 17092 23196 17098 23208
rect 2501 23171 2559 23177
rect 2501 23168 2513 23171
rect 2056 23140 2513 23168
rect 2056 23109 2084 23140
rect 2501 23137 2513 23140
rect 2547 23137 2559 23171
rect 2501 23131 2559 23137
rect 10870 23128 10876 23180
rect 10928 23128 10934 23180
rect 11146 23128 11152 23180
rect 11204 23128 11210 23180
rect 15470 23128 15476 23180
rect 15528 23168 15534 23180
rect 17957 23171 18015 23177
rect 17957 23168 17969 23171
rect 15528 23140 17969 23168
rect 15528 23128 15534 23140
rect 17957 23137 17969 23140
rect 18003 23168 18015 23171
rect 18230 23168 18236 23180
rect 18003 23140 18236 23168
rect 18003 23137 18015 23140
rect 17957 23131 18015 23137
rect 18230 23128 18236 23140
rect 18288 23128 18294 23180
rect 2041 23103 2099 23109
rect 2041 23069 2053 23103
rect 2087 23069 2099 23103
rect 2041 23063 2099 23069
rect 2130 23060 2136 23112
rect 2188 23060 2194 23112
rect 10686 23060 10692 23112
rect 10744 23100 10750 23112
rect 10781 23103 10839 23109
rect 10781 23100 10793 23103
rect 10744 23072 10793 23100
rect 10744 23060 10750 23072
rect 10781 23069 10793 23072
rect 10827 23069 10839 23103
rect 10781 23063 10839 23069
rect 14458 23060 14464 23112
rect 14516 23100 14522 23112
rect 14645 23103 14703 23109
rect 14645 23100 14657 23103
rect 14516 23072 14657 23100
rect 14516 23060 14522 23072
rect 14645 23069 14657 23072
rect 14691 23069 14703 23103
rect 14645 23063 14703 23069
rect 16393 23103 16451 23109
rect 16393 23069 16405 23103
rect 16439 23100 16451 23103
rect 18708 23100 18736 23267
rect 19334 23264 19340 23276
rect 19392 23264 19398 23316
rect 29917 23307 29975 23313
rect 29917 23273 29929 23307
rect 29963 23304 29975 23307
rect 30006 23304 30012 23316
rect 29963 23276 30012 23304
rect 29963 23273 29975 23276
rect 29917 23267 29975 23273
rect 30006 23264 30012 23276
rect 30064 23304 30070 23316
rect 30374 23304 30380 23316
rect 30064 23276 30380 23304
rect 30064 23264 30070 23276
rect 30374 23264 30380 23276
rect 30432 23264 30438 23316
rect 30466 23264 30472 23316
rect 30524 23304 30530 23316
rect 30745 23307 30803 23313
rect 30745 23304 30757 23307
rect 30524 23276 30757 23304
rect 30524 23264 30530 23276
rect 30745 23273 30757 23276
rect 30791 23273 30803 23307
rect 30745 23267 30803 23273
rect 31110 23264 31116 23316
rect 31168 23304 31174 23316
rect 31205 23307 31263 23313
rect 31205 23304 31217 23307
rect 31168 23276 31217 23304
rect 31168 23264 31174 23276
rect 31205 23273 31217 23276
rect 31251 23304 31263 23307
rect 32582 23304 32588 23316
rect 31251 23276 32588 23304
rect 31251 23273 31263 23276
rect 31205 23267 31263 23273
rect 32582 23264 32588 23276
rect 32640 23264 32646 23316
rect 33134 23264 33140 23316
rect 33192 23304 33198 23316
rect 33321 23307 33379 23313
rect 33321 23304 33333 23307
rect 33192 23276 33333 23304
rect 33192 23264 33198 23276
rect 33321 23273 33333 23276
rect 33367 23273 33379 23307
rect 33321 23267 33379 23273
rect 35986 23264 35992 23316
rect 36044 23304 36050 23316
rect 36170 23304 36176 23316
rect 36044 23276 36176 23304
rect 36044 23264 36050 23276
rect 36170 23264 36176 23276
rect 36228 23264 36234 23316
rect 40310 23264 40316 23316
rect 40368 23304 40374 23316
rect 40497 23307 40555 23313
rect 40497 23304 40509 23307
rect 40368 23276 40509 23304
rect 40368 23264 40374 23276
rect 40497 23273 40509 23276
rect 40543 23273 40555 23307
rect 40497 23267 40555 23273
rect 42153 23307 42211 23313
rect 42153 23273 42165 23307
rect 42199 23304 42211 23307
rect 42334 23304 42340 23316
rect 42199 23276 42340 23304
rect 42199 23273 42211 23276
rect 42153 23267 42211 23273
rect 42334 23264 42340 23276
rect 42392 23264 42398 23316
rect 48222 23304 48228 23316
rect 42628 23276 48228 23304
rect 31386 23236 31392 23248
rect 30392 23208 31392 23236
rect 30282 23168 30288 23180
rect 16439 23072 18736 23100
rect 22066 23140 30288 23168
rect 16439 23069 16451 23072
rect 16393 23063 16451 23069
rect 13722 22992 13728 23044
rect 13780 23032 13786 23044
rect 16408 23032 16436 23063
rect 13780 23004 16436 23032
rect 13780 22992 13786 23004
rect 16666 22992 16672 23044
rect 16724 23032 16730 23044
rect 17129 23035 17187 23041
rect 17129 23032 17141 23035
rect 16724 23004 17141 23032
rect 16724 22992 16730 23004
rect 17129 23001 17141 23004
rect 17175 23001 17187 23035
rect 17129 22995 17187 23001
rect 17678 22992 17684 23044
rect 17736 23032 17742 23044
rect 17773 23035 17831 23041
rect 17773 23032 17785 23035
rect 17736 23004 17785 23032
rect 17736 22992 17742 23004
rect 17773 23001 17785 23004
rect 17819 23001 17831 23035
rect 17773 22995 17831 23001
rect 18233 23035 18291 23041
rect 18233 23001 18245 23035
rect 18279 23032 18291 23035
rect 18509 23035 18567 23041
rect 18509 23032 18521 23035
rect 18279 23004 18521 23032
rect 18279 23001 18291 23004
rect 18233 22995 18291 23001
rect 18509 23001 18521 23004
rect 18555 23032 18567 23035
rect 19150 23032 19156 23044
rect 18555 23004 19156 23032
rect 18555 23001 18567 23004
rect 18509 22995 18567 23001
rect 19150 22992 19156 23004
rect 19208 23032 19214 23044
rect 22066 23032 22094 23140
rect 30282 23128 30288 23140
rect 30340 23128 30346 23180
rect 29641 23103 29699 23109
rect 29641 23069 29653 23103
rect 29687 23100 29699 23103
rect 29733 23103 29791 23109
rect 29733 23100 29745 23103
rect 29687 23072 29745 23100
rect 29687 23069 29699 23072
rect 29641 23063 29699 23069
rect 29733 23069 29745 23072
rect 29779 23100 29791 23103
rect 29822 23100 29828 23112
rect 29779 23072 29828 23100
rect 29779 23069 29791 23072
rect 29733 23063 29791 23069
rect 29822 23060 29828 23072
rect 29880 23060 29886 23112
rect 29914 23060 29920 23112
rect 29972 23060 29978 23112
rect 30098 23060 30104 23112
rect 30156 23060 30162 23112
rect 30392 23100 30420 23208
rect 31386 23196 31392 23208
rect 31444 23236 31450 23248
rect 32858 23236 32864 23248
rect 31444 23208 32864 23236
rect 31444 23196 31450 23208
rect 32858 23196 32864 23208
rect 32916 23196 32922 23248
rect 35805 23239 35863 23245
rect 35805 23205 35817 23239
rect 35851 23236 35863 23239
rect 35851 23208 36308 23236
rect 35851 23205 35863 23208
rect 35805 23199 35863 23205
rect 31202 23168 31208 23180
rect 30484 23140 31208 23168
rect 30484 23109 30512 23140
rect 31202 23128 31208 23140
rect 31260 23128 31266 23180
rect 32582 23128 32588 23180
rect 32640 23168 32646 23180
rect 33781 23171 33839 23177
rect 33781 23168 33793 23171
rect 32640 23140 33793 23168
rect 32640 23128 32646 23140
rect 33781 23137 33793 23140
rect 33827 23137 33839 23171
rect 36170 23168 36176 23180
rect 33781 23131 33839 23137
rect 35452 23140 36176 23168
rect 30300 23072 30420 23100
rect 30469 23103 30527 23109
rect 19208 23004 22094 23032
rect 29932 23032 29960 23060
rect 30300 23041 30328 23072
rect 30469 23069 30481 23103
rect 30515 23069 30527 23103
rect 30469 23063 30527 23069
rect 30285 23035 30343 23041
rect 30285 23032 30297 23035
rect 29932 23004 30297 23032
rect 19208 22992 19214 23004
rect 30285 23001 30297 23004
rect 30331 23001 30343 23035
rect 30285 22995 30343 23001
rect 30374 22992 30380 23044
rect 30432 22992 30438 23044
rect 934 22924 940 22976
rect 992 22964 998 22976
rect 1857 22967 1915 22973
rect 1857 22964 1869 22967
rect 992 22936 1869 22964
rect 992 22924 998 22936
rect 1857 22933 1869 22936
rect 1903 22933 1915 22967
rect 1857 22927 1915 22933
rect 13078 22924 13084 22976
rect 13136 22964 13142 22976
rect 14093 22967 14151 22973
rect 14093 22964 14105 22967
rect 13136 22936 14105 22964
rect 13136 22924 13142 22936
rect 14093 22933 14105 22936
rect 14139 22933 14151 22967
rect 14093 22927 14151 22933
rect 16942 22924 16948 22976
rect 17000 22964 17006 22976
rect 17586 22973 17592 22976
rect 17563 22967 17592 22973
rect 17563 22964 17575 22967
rect 17000 22936 17575 22964
rect 17000 22924 17006 22936
rect 17563 22933 17575 22936
rect 17563 22927 17592 22933
rect 17586 22924 17592 22927
rect 17644 22924 17650 22976
rect 18598 22924 18604 22976
rect 18656 22964 18662 22976
rect 19242 22964 19248 22976
rect 18656 22936 19248 22964
rect 18656 22924 18662 22936
rect 19242 22924 19248 22936
rect 19300 22964 19306 22976
rect 19337 22967 19395 22973
rect 19337 22964 19349 22967
rect 19300 22936 19349 22964
rect 19300 22924 19306 22936
rect 19337 22933 19349 22936
rect 19383 22933 19395 22967
rect 19337 22927 19395 22933
rect 30098 22924 30104 22976
rect 30156 22964 30162 22976
rect 30484 22964 30512 23063
rect 30650 23060 30656 23112
rect 30708 23100 30714 23112
rect 30929 23103 30987 23109
rect 30929 23100 30941 23103
rect 30708 23072 30941 23100
rect 30708 23060 30714 23072
rect 30929 23069 30941 23072
rect 30975 23069 30987 23103
rect 30929 23063 30987 23069
rect 31021 23103 31079 23109
rect 31021 23069 31033 23103
rect 31067 23069 31079 23103
rect 31021 23063 31079 23069
rect 31036 23032 31064 23063
rect 31294 23060 31300 23112
rect 31352 23060 31358 23112
rect 31846 23060 31852 23112
rect 31904 23100 31910 23112
rect 32306 23100 32312 23112
rect 31904 23072 32312 23100
rect 31904 23060 31910 23072
rect 32306 23060 32312 23072
rect 32364 23100 32370 23112
rect 33505 23103 33563 23109
rect 33505 23100 33517 23103
rect 32364 23072 33517 23100
rect 32364 23060 32370 23072
rect 33505 23069 33517 23072
rect 33551 23069 33563 23103
rect 33505 23063 33563 23069
rect 33597 23103 33655 23109
rect 33597 23069 33609 23103
rect 33643 23069 33655 23103
rect 33597 23063 33655 23069
rect 33873 23103 33931 23109
rect 33873 23069 33885 23103
rect 33919 23100 33931 23103
rect 34790 23100 34796 23112
rect 33919 23072 34796 23100
rect 33919 23069 33931 23072
rect 33873 23063 33931 23069
rect 30668 23004 31064 23032
rect 30668 22973 30696 23004
rect 31754 22992 31760 23044
rect 31812 23032 31818 23044
rect 33226 23032 33232 23044
rect 31812 23004 33232 23032
rect 31812 22992 31818 23004
rect 33226 22992 33232 23004
rect 33284 22992 33290 23044
rect 33612 23032 33640 23063
rect 34790 23060 34796 23072
rect 34848 23060 34854 23112
rect 35253 23103 35311 23109
rect 35253 23069 35265 23103
rect 35299 23100 35311 23103
rect 35342 23100 35348 23112
rect 35299 23072 35348 23100
rect 35299 23069 35311 23072
rect 35253 23063 35311 23069
rect 35342 23060 35348 23072
rect 35400 23060 35406 23112
rect 35452 23109 35480 23140
rect 36170 23128 36176 23140
rect 36228 23128 36234 23180
rect 36280 23109 36308 23208
rect 39942 23196 39948 23248
rect 40000 23236 40006 23248
rect 42628 23236 42656 23276
rect 48222 23264 48228 23276
rect 48280 23264 48286 23316
rect 48314 23264 48320 23316
rect 48372 23304 48378 23316
rect 49145 23307 49203 23313
rect 49145 23304 49157 23307
rect 48372 23276 49157 23304
rect 48372 23264 48378 23276
rect 49145 23273 49157 23276
rect 49191 23273 49203 23307
rect 49145 23267 49203 23273
rect 50890 23264 50896 23316
rect 50948 23304 50954 23316
rect 51534 23304 51540 23316
rect 50948 23276 51540 23304
rect 50948 23264 50954 23276
rect 51534 23264 51540 23276
rect 51592 23264 51598 23316
rect 51902 23264 51908 23316
rect 51960 23304 51966 23316
rect 53377 23307 53435 23313
rect 53377 23304 53389 23307
rect 51960 23276 53389 23304
rect 51960 23264 51966 23276
rect 53377 23273 53389 23276
rect 53423 23304 53435 23307
rect 53745 23307 53803 23313
rect 53745 23304 53757 23307
rect 53423 23276 53757 23304
rect 53423 23273 53435 23276
rect 53377 23267 53435 23273
rect 53745 23273 53757 23276
rect 53791 23304 53803 23307
rect 55214 23304 55220 23316
rect 53791 23276 55220 23304
rect 53791 23273 53803 23276
rect 53745 23267 53803 23273
rect 55214 23264 55220 23276
rect 55272 23264 55278 23316
rect 55306 23264 55312 23316
rect 55364 23304 55370 23316
rect 55582 23304 55588 23316
rect 55364 23276 55588 23304
rect 55364 23264 55370 23276
rect 55582 23264 55588 23276
rect 55640 23264 55646 23316
rect 58526 23264 58532 23316
rect 58584 23264 58590 23316
rect 40000 23208 42656 23236
rect 40000 23196 40006 23208
rect 37274 23168 37280 23180
rect 36372 23140 37280 23168
rect 36372 23109 36400 23140
rect 37274 23128 37280 23140
rect 37332 23128 37338 23180
rect 39758 23128 39764 23180
rect 39816 23168 39822 23180
rect 41432 23177 41460 23208
rect 42702 23196 42708 23248
rect 42760 23236 42766 23248
rect 42760 23208 44588 23236
rect 42760 23196 42766 23208
rect 41417 23171 41475 23177
rect 39816 23140 39988 23168
rect 39816 23128 39822 23140
rect 35437 23103 35495 23109
rect 35437 23069 35449 23103
rect 35483 23069 35495 23103
rect 35437 23063 35495 23069
rect 35621 23103 35679 23109
rect 35621 23069 35633 23103
rect 35667 23069 35679 23103
rect 35621 23063 35679 23069
rect 36265 23103 36323 23109
rect 36265 23069 36277 23103
rect 36311 23069 36323 23103
rect 36265 23063 36323 23069
rect 36357 23103 36415 23109
rect 36357 23069 36369 23103
rect 36403 23069 36415 23103
rect 36357 23063 36415 23069
rect 34698 23032 34704 23044
rect 33612 23004 34704 23032
rect 34698 22992 34704 23004
rect 34756 22992 34762 23044
rect 35529 23035 35587 23041
rect 35529 23001 35541 23035
rect 35575 23001 35587 23035
rect 35636 23032 35664 23063
rect 36538 23060 36544 23112
rect 36596 23060 36602 23112
rect 36633 23103 36691 23109
rect 36633 23069 36645 23103
rect 36679 23100 36691 23103
rect 36814 23100 36820 23112
rect 36679 23072 36820 23100
rect 36679 23069 36691 23072
rect 36633 23063 36691 23069
rect 36814 23060 36820 23072
rect 36872 23100 36878 23112
rect 36909 23103 36967 23109
rect 36909 23100 36921 23103
rect 36872 23072 36921 23100
rect 36872 23060 36878 23072
rect 36909 23069 36921 23072
rect 36955 23069 36967 23103
rect 36909 23063 36967 23069
rect 39114 23060 39120 23112
rect 39172 23100 39178 23112
rect 39960 23109 39988 23140
rect 41417 23137 41429 23171
rect 41463 23137 41475 23171
rect 41417 23131 41475 23137
rect 42518 23128 42524 23180
rect 42576 23128 42582 23180
rect 43070 23128 43076 23180
rect 43128 23128 43134 23180
rect 44082 23128 44088 23180
rect 44140 23168 44146 23180
rect 44177 23171 44235 23177
rect 44177 23168 44189 23171
rect 44140 23140 44189 23168
rect 44140 23128 44146 23140
rect 44177 23137 44189 23140
rect 44223 23137 44235 23171
rect 44177 23131 44235 23137
rect 44266 23128 44272 23180
rect 44324 23128 44330 23180
rect 44461 23171 44519 23177
rect 44461 23137 44473 23171
rect 44507 23168 44519 23171
rect 44560 23168 44588 23208
rect 44836 23208 45324 23236
rect 44726 23168 44732 23180
rect 44507 23140 44732 23168
rect 44507 23137 44519 23140
rect 44461 23131 44519 23137
rect 44726 23128 44732 23140
rect 44784 23128 44790 23180
rect 39853 23103 39911 23109
rect 39853 23100 39865 23103
rect 39172 23072 39865 23100
rect 39172 23060 39178 23072
rect 39853 23069 39865 23072
rect 39899 23069 39911 23103
rect 39853 23063 39911 23069
rect 39946 23103 40004 23109
rect 39946 23069 39958 23103
rect 39992 23069 40004 23103
rect 40318 23103 40376 23109
rect 40318 23100 40330 23103
rect 39946 23063 40004 23069
rect 40052 23072 40330 23100
rect 35989 23035 36047 23041
rect 35989 23032 36001 23035
rect 35636 23004 36001 23032
rect 35529 22995 35587 23001
rect 35989 23001 36001 23004
rect 36035 23032 36047 23035
rect 37182 23032 37188 23044
rect 36035 23004 37188 23032
rect 36035 23001 36047 23004
rect 35989 22995 36047 23001
rect 30156 22936 30512 22964
rect 30653 22967 30711 22973
rect 30156 22924 30162 22936
rect 30653 22933 30665 22967
rect 30699 22933 30711 22967
rect 30653 22927 30711 22933
rect 31570 22924 31576 22976
rect 31628 22964 31634 22976
rect 35544 22964 35572 22995
rect 37182 22992 37188 23004
rect 37240 22992 37246 23044
rect 39574 22992 39580 23044
rect 39632 23032 39638 23044
rect 40052 23032 40080 23072
rect 40318 23069 40330 23072
rect 40364 23100 40376 23103
rect 41877 23103 41935 23109
rect 41877 23100 41889 23103
rect 40364 23072 41889 23100
rect 40364 23069 40376 23072
rect 40318 23063 40376 23069
rect 41877 23069 41889 23072
rect 41923 23069 41935 23103
rect 41877 23063 41935 23069
rect 39632 23004 40080 23032
rect 40129 23035 40187 23041
rect 39632 22992 39638 23004
rect 40129 23001 40141 23035
rect 40175 23001 40187 23035
rect 40129 22995 40187 23001
rect 31628 22936 35572 22964
rect 31628 22924 31634 22936
rect 36170 22924 36176 22976
rect 36228 22924 36234 22976
rect 36538 22924 36544 22976
rect 36596 22964 36602 22976
rect 36817 22967 36875 22973
rect 36817 22964 36829 22967
rect 36596 22936 36829 22964
rect 36596 22924 36602 22936
rect 36817 22933 36829 22936
rect 36863 22933 36875 22967
rect 40144 22964 40172 22995
rect 40218 22992 40224 23044
rect 40276 22992 40282 23044
rect 40494 22964 40500 22976
rect 40144 22936 40500 22964
rect 36817 22927 36875 22933
rect 40494 22924 40500 22936
rect 40552 22964 40558 22976
rect 40589 22967 40647 22973
rect 40589 22964 40601 22967
rect 40552 22936 40601 22964
rect 40552 22924 40558 22936
rect 40589 22933 40601 22936
rect 40635 22933 40647 22967
rect 41892 22964 41920 23063
rect 42242 23060 42248 23112
rect 42300 23060 42306 23112
rect 42536 23100 42564 23128
rect 42978 23100 42984 23112
rect 42536 23072 42984 23100
rect 42978 23060 42984 23072
rect 43036 23100 43042 23112
rect 43622 23100 43628 23112
rect 43036 23072 43628 23100
rect 43036 23060 43042 23072
rect 43622 23060 43628 23072
rect 43680 23100 43686 23112
rect 43717 23103 43775 23109
rect 43717 23100 43729 23103
rect 43680 23072 43729 23100
rect 43680 23060 43686 23072
rect 43717 23069 43729 23072
rect 43763 23069 43775 23103
rect 43717 23063 43775 23069
rect 43806 23060 43812 23112
rect 43864 23060 43870 23112
rect 43898 23060 43904 23112
rect 43956 23060 43962 23112
rect 44361 23103 44419 23109
rect 44361 23069 44373 23103
rect 44407 23100 44419 23103
rect 44836 23100 44864 23208
rect 45186 23128 45192 23180
rect 45244 23128 45250 23180
rect 45296 23177 45324 23208
rect 45370 23196 45376 23248
rect 45428 23196 45434 23248
rect 49050 23196 49056 23248
rect 49108 23236 49114 23248
rect 49108 23208 53328 23236
rect 49108 23196 49114 23208
rect 45281 23171 45339 23177
rect 45281 23137 45293 23171
rect 45327 23137 45339 23171
rect 45388 23168 45416 23196
rect 45465 23171 45523 23177
rect 45465 23168 45477 23171
rect 45388 23140 45477 23168
rect 45281 23131 45339 23137
rect 45465 23137 45477 23140
rect 45511 23137 45523 23171
rect 45465 23131 45523 23137
rect 47581 23171 47639 23177
rect 47581 23137 47593 23171
rect 47627 23168 47639 23171
rect 48038 23168 48044 23180
rect 47627 23140 48044 23168
rect 47627 23137 47639 23140
rect 47581 23131 47639 23137
rect 48038 23128 48044 23140
rect 48096 23128 48102 23180
rect 48590 23128 48596 23180
rect 48648 23168 48654 23180
rect 49142 23168 49148 23180
rect 48648 23140 49148 23168
rect 48648 23128 48654 23140
rect 49142 23128 49148 23140
rect 49200 23168 49206 23180
rect 49513 23171 49571 23177
rect 49513 23168 49525 23171
rect 49200 23140 49525 23168
rect 49200 23128 49206 23140
rect 49513 23137 49525 23140
rect 49559 23137 49571 23171
rect 52914 23168 52920 23180
rect 49513 23131 49571 23137
rect 51460 23140 52920 23168
rect 44407 23072 44864 23100
rect 44407 23069 44419 23072
rect 44361 23063 44419 23069
rect 41969 23035 42027 23041
rect 41969 23001 41981 23035
rect 42015 23032 42027 23035
rect 42518 23032 42524 23044
rect 42015 23004 42524 23032
rect 42015 23001 42027 23004
rect 41969 22995 42027 23001
rect 42518 22992 42524 23004
rect 42576 22992 42582 23044
rect 42886 22992 42892 23044
rect 42944 23032 42950 23044
rect 43257 23035 43315 23041
rect 43257 23032 43269 23035
rect 42944 23004 43269 23032
rect 42944 22992 42950 23004
rect 43257 23001 43269 23004
rect 43303 23001 43315 23035
rect 43257 22995 43315 23001
rect 42610 22964 42616 22976
rect 41892 22936 42616 22964
rect 40589 22927 40647 22933
rect 42610 22924 42616 22936
rect 42668 22964 42674 22976
rect 43438 22964 43444 22976
rect 42668 22936 43444 22964
rect 42668 22924 42674 22936
rect 43438 22924 43444 22936
rect 43496 22964 43502 22976
rect 44376 22964 44404 23063
rect 45370 23060 45376 23112
rect 45428 23060 45434 23112
rect 46014 23060 46020 23112
rect 46072 23100 46078 23112
rect 46109 23103 46167 23109
rect 46109 23100 46121 23103
rect 46072 23072 46121 23100
rect 46072 23060 46078 23072
rect 46109 23069 46121 23072
rect 46155 23069 46167 23103
rect 46109 23063 46167 23069
rect 46382 23060 46388 23112
rect 46440 23060 46446 23112
rect 47302 23060 47308 23112
rect 47360 23060 47366 23112
rect 48682 23060 48688 23112
rect 48740 23060 48746 23112
rect 49326 23060 49332 23112
rect 49384 23060 49390 23112
rect 50614 23100 50620 23112
rect 49436 23072 50620 23100
rect 44726 22992 44732 23044
rect 44784 23032 44790 23044
rect 45186 23032 45192 23044
rect 44784 23004 45192 23032
rect 44784 22992 44790 23004
rect 45186 22992 45192 23004
rect 45244 23032 45250 23044
rect 46477 23035 46535 23041
rect 46477 23032 46489 23035
rect 45244 23004 46489 23032
rect 45244 22992 45250 23004
rect 46477 23001 46489 23004
rect 46523 23032 46535 23035
rect 46658 23032 46664 23044
rect 46523 23004 46664 23032
rect 46523 23001 46535 23004
rect 46477 22995 46535 23001
rect 46658 22992 46664 23004
rect 46716 22992 46722 23044
rect 49436 23032 49464 23072
rect 50614 23060 50620 23072
rect 50672 23060 50678 23112
rect 51074 23060 51080 23112
rect 51132 23060 51138 23112
rect 51225 23103 51283 23109
rect 51225 23069 51237 23103
rect 51271 23100 51283 23103
rect 51460 23100 51488 23140
rect 52914 23128 52920 23140
rect 52972 23128 52978 23180
rect 51271 23072 51488 23100
rect 51271 23069 51283 23072
rect 51225 23063 51283 23069
rect 51534 23060 51540 23112
rect 51592 23109 51598 23112
rect 51592 23063 51600 23109
rect 51592 23060 51598 23063
rect 52270 23060 52276 23112
rect 52328 23100 52334 23112
rect 53101 23103 53159 23109
rect 53101 23100 53113 23103
rect 52328 23072 53113 23100
rect 52328 23060 52334 23072
rect 53101 23069 53113 23072
rect 53147 23069 53159 23103
rect 53101 23063 53159 23069
rect 53190 23060 53196 23112
rect 53248 23060 53254 23112
rect 48884 23004 49464 23032
rect 43496 22936 44404 22964
rect 43496 22924 43502 22936
rect 44634 22924 44640 22976
rect 44692 22924 44698 22976
rect 45002 22924 45008 22976
rect 45060 22924 45066 22976
rect 45094 22924 45100 22976
rect 45152 22964 45158 22976
rect 48884 22964 48912 23004
rect 49878 22992 49884 23044
rect 49936 23032 49942 23044
rect 50890 23032 50896 23044
rect 49936 23004 50896 23032
rect 49936 22992 49942 23004
rect 50890 22992 50896 23004
rect 50948 22992 50954 23044
rect 51353 23035 51411 23041
rect 51353 23032 51365 23035
rect 51046 23004 51365 23032
rect 45152 22936 48912 22964
rect 49053 22967 49111 22973
rect 45152 22924 45158 22936
rect 49053 22933 49065 22967
rect 49099 22964 49111 22967
rect 49234 22964 49240 22976
rect 49099 22936 49240 22964
rect 49099 22933 49111 22936
rect 49053 22927 49111 22933
rect 49234 22924 49240 22936
rect 49292 22924 49298 22976
rect 49694 22924 49700 22976
rect 49752 22964 49758 22976
rect 50154 22964 50160 22976
rect 49752 22936 50160 22964
rect 49752 22924 49758 22936
rect 50154 22924 50160 22936
rect 50212 22924 50218 22976
rect 50706 22924 50712 22976
rect 50764 22964 50770 22976
rect 51046 22964 51074 23004
rect 51353 23001 51365 23004
rect 51399 23001 51411 23035
rect 51353 22995 51411 23001
rect 51445 23035 51503 23041
rect 51445 23001 51457 23035
rect 51491 23032 51503 23035
rect 52546 23032 52552 23044
rect 51491 23004 52552 23032
rect 51491 23001 51503 23004
rect 51445 22995 51503 23001
rect 52546 22992 52552 23004
rect 52604 22992 52610 23044
rect 53300 23032 53328 23208
rect 54478 23128 54484 23180
rect 54536 23168 54542 23180
rect 56226 23168 56232 23180
rect 54536 23140 56232 23168
rect 54536 23128 54542 23140
rect 56226 23128 56232 23140
rect 56284 23128 56290 23180
rect 53469 23103 53527 23109
rect 53469 23069 53481 23103
rect 53515 23100 53527 23103
rect 54021 23103 54079 23109
rect 54021 23100 54033 23103
rect 53515 23072 54033 23100
rect 53515 23069 53527 23072
rect 53469 23063 53527 23069
rect 54021 23069 54033 23072
rect 54067 23069 54079 23103
rect 54021 23063 54079 23069
rect 54570 23060 54576 23112
rect 54628 23060 54634 23112
rect 57054 23060 57060 23112
rect 57112 23100 57118 23112
rect 57149 23103 57207 23109
rect 57149 23100 57161 23103
rect 57112 23072 57161 23100
rect 57112 23060 57118 23072
rect 57149 23069 57161 23072
rect 57195 23069 57207 23103
rect 57149 23063 57207 23069
rect 53653 23035 53711 23041
rect 53653 23032 53665 23035
rect 53300 23004 53665 23032
rect 53653 23001 53665 23004
rect 53699 23001 53711 23035
rect 53653 22995 53711 23001
rect 56226 22992 56232 23044
rect 56284 22992 56290 23044
rect 56781 23035 56839 23041
rect 56781 23001 56793 23035
rect 56827 23001 56839 23035
rect 56781 22995 56839 23001
rect 50764 22936 51074 22964
rect 50764 22924 50770 22936
rect 51534 22924 51540 22976
rect 51592 22964 51598 22976
rect 51721 22967 51779 22973
rect 51721 22964 51733 22967
rect 51592 22936 51733 22964
rect 51592 22924 51598 22936
rect 51721 22933 51733 22936
rect 51767 22933 51779 22967
rect 51721 22927 51779 22933
rect 52917 22967 52975 22973
rect 52917 22933 52929 22967
rect 52963 22964 52975 22967
rect 53006 22964 53012 22976
rect 52963 22936 53012 22964
rect 52963 22933 52975 22936
rect 52917 22927 52975 22933
rect 53006 22924 53012 22936
rect 53064 22924 53070 22976
rect 54846 22924 54852 22976
rect 54904 22964 54910 22976
rect 55306 22964 55312 22976
rect 54904 22936 55312 22964
rect 54904 22924 54910 22936
rect 55306 22924 55312 22936
rect 55364 22924 55370 22976
rect 55398 22924 55404 22976
rect 55456 22964 55462 22976
rect 56796 22964 56824 22995
rect 56870 22992 56876 23044
rect 56928 23032 56934 23044
rect 57394 23035 57452 23041
rect 57394 23032 57406 23035
rect 56928 23004 57406 23032
rect 56928 22992 56934 23004
rect 57394 23001 57406 23004
rect 57440 23001 57452 23035
rect 57394 22995 57452 23001
rect 55456 22936 56824 22964
rect 55456 22924 55462 22936
rect 1104 22874 78844 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 66314 22874
rect 66366 22822 66378 22874
rect 66430 22822 66442 22874
rect 66494 22822 66506 22874
rect 66558 22822 66570 22874
rect 66622 22822 78844 22874
rect 1104 22800 78844 22822
rect 10686 22720 10692 22772
rect 10744 22720 10750 22772
rect 13633 22763 13691 22769
rect 13633 22729 13645 22763
rect 13679 22760 13691 22763
rect 14458 22760 14464 22772
rect 13679 22732 14464 22760
rect 13679 22729 13691 22732
rect 13633 22723 13691 22729
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 17126 22720 17132 22772
rect 17184 22760 17190 22772
rect 17862 22760 17868 22772
rect 17184 22732 17868 22760
rect 17184 22720 17190 22732
rect 17862 22720 17868 22732
rect 17920 22760 17926 22772
rect 18509 22763 18567 22769
rect 18509 22760 18521 22763
rect 17920 22732 18521 22760
rect 17920 22720 17926 22732
rect 18509 22729 18521 22732
rect 18555 22729 18567 22763
rect 18509 22723 18567 22729
rect 19242 22720 19248 22772
rect 19300 22760 19306 22772
rect 19429 22763 19487 22769
rect 19429 22760 19441 22763
rect 19300 22732 19441 22760
rect 19300 22720 19306 22732
rect 19429 22729 19441 22732
rect 19475 22729 19487 22763
rect 30466 22760 30472 22772
rect 19429 22723 19487 22729
rect 30024 22732 30472 22760
rect 9674 22652 9680 22704
rect 9732 22652 9738 22704
rect 10505 22695 10563 22701
rect 10505 22661 10517 22695
rect 10551 22692 10563 22695
rect 11609 22695 11667 22701
rect 11609 22692 11621 22695
rect 10551 22664 11621 22692
rect 10551 22661 10563 22664
rect 10505 22655 10563 22661
rect 11609 22661 11621 22664
rect 11655 22692 11667 22695
rect 13722 22692 13728 22704
rect 11655 22664 13728 22692
rect 11655 22661 11667 22664
rect 11609 22655 11667 22661
rect 13722 22652 13728 22664
rect 13780 22652 13786 22704
rect 15470 22692 15476 22704
rect 14674 22664 15476 22692
rect 15470 22652 15476 22664
rect 15528 22652 15534 22704
rect 18230 22652 18236 22704
rect 18288 22692 18294 22704
rect 19337 22695 19395 22701
rect 19337 22692 19349 22695
rect 18288 22664 19349 22692
rect 18288 22652 18294 22664
rect 19337 22661 19349 22664
rect 19383 22692 19395 22695
rect 19797 22695 19855 22701
rect 19797 22692 19809 22695
rect 19383 22664 19809 22692
rect 19383 22661 19395 22664
rect 19337 22655 19395 22661
rect 19797 22661 19809 22664
rect 19843 22661 19855 22695
rect 30024 22692 30052 22732
rect 30466 22720 30472 22732
rect 30524 22760 30530 22772
rect 30653 22763 30711 22769
rect 30653 22760 30665 22763
rect 30524 22732 30665 22760
rect 30524 22720 30530 22732
rect 30653 22729 30665 22732
rect 30699 22760 30711 22763
rect 30834 22760 30840 22772
rect 30699 22732 30840 22760
rect 30699 22729 30711 22732
rect 30653 22723 30711 22729
rect 30834 22720 30840 22732
rect 30892 22720 30898 22772
rect 32030 22720 32036 22772
rect 32088 22760 32094 22772
rect 32674 22760 32680 22772
rect 32088 22732 32680 22760
rect 32088 22720 32094 22732
rect 32674 22720 32680 22732
rect 32732 22720 32738 22772
rect 32769 22763 32827 22769
rect 32769 22729 32781 22763
rect 32815 22729 32827 22763
rect 38289 22763 38347 22769
rect 38289 22760 38301 22763
rect 32769 22723 32827 22729
rect 33244 22732 37596 22760
rect 32784 22692 32812 22723
rect 29394 22664 30052 22692
rect 32416 22664 32812 22692
rect 19797 22655 19855 22661
rect 13078 22584 13084 22636
rect 13136 22584 13142 22636
rect 18046 22584 18052 22636
rect 18104 22624 18110 22636
rect 18598 22624 18604 22636
rect 18104 22596 18604 22624
rect 18104 22584 18110 22596
rect 18598 22584 18604 22596
rect 18656 22584 18662 22636
rect 27985 22627 28043 22633
rect 27985 22593 27997 22627
rect 28031 22624 28043 22627
rect 28442 22624 28448 22636
rect 28031 22596 28448 22624
rect 28031 22593 28043 22596
rect 27985 22587 28043 22593
rect 28442 22584 28448 22596
rect 28500 22584 28506 22636
rect 30098 22584 30104 22636
rect 30156 22584 30162 22636
rect 30190 22584 30196 22636
rect 30248 22584 30254 22636
rect 30285 22627 30343 22633
rect 30285 22593 30297 22627
rect 30331 22593 30343 22627
rect 30285 22587 30343 22593
rect 11054 22516 11060 22568
rect 11112 22556 11118 22568
rect 11241 22559 11299 22565
rect 11241 22556 11253 22559
rect 11112 22528 11253 22556
rect 11112 22516 11118 22528
rect 11241 22525 11253 22528
rect 11287 22525 11299 22559
rect 11241 22519 11299 22525
rect 12434 22516 12440 22568
rect 12492 22556 12498 22568
rect 12894 22556 12900 22568
rect 12492 22528 12900 22556
rect 12492 22516 12498 22528
rect 12894 22516 12900 22528
rect 12952 22556 12958 22568
rect 12989 22559 13047 22565
rect 12989 22556 13001 22559
rect 12952 22528 13001 22556
rect 12952 22516 12958 22528
rect 12989 22525 13001 22528
rect 13035 22525 13047 22559
rect 12989 22519 13047 22525
rect 15102 22516 15108 22568
rect 15160 22516 15166 22568
rect 15381 22559 15439 22565
rect 15381 22525 15393 22559
rect 15427 22556 15439 22559
rect 16666 22556 16672 22568
rect 15427 22528 16672 22556
rect 15427 22525 15439 22528
rect 15381 22519 15439 22525
rect 13449 22491 13507 22497
rect 13449 22457 13461 22491
rect 13495 22488 13507 22491
rect 14090 22488 14096 22500
rect 13495 22460 14096 22488
rect 13495 22457 13507 22460
rect 13449 22451 13507 22457
rect 14090 22448 14096 22460
rect 14148 22448 14154 22500
rect 14366 22380 14372 22432
rect 14424 22420 14430 22432
rect 15396 22420 15424 22519
rect 16666 22516 16672 22528
rect 16724 22516 16730 22568
rect 16942 22516 16948 22568
rect 17000 22516 17006 22568
rect 17954 22516 17960 22568
rect 18012 22556 18018 22568
rect 18417 22559 18475 22565
rect 18417 22556 18429 22559
rect 18012 22528 18429 22556
rect 18012 22516 18018 22528
rect 18417 22525 18429 22528
rect 18463 22556 18475 22559
rect 19061 22559 19119 22565
rect 19061 22556 19073 22559
rect 18463 22528 19073 22556
rect 18463 22525 18475 22528
rect 18417 22519 18475 22525
rect 19061 22525 19073 22528
rect 19107 22525 19119 22559
rect 19061 22519 19119 22525
rect 28353 22559 28411 22565
rect 28353 22525 28365 22559
rect 28399 22556 28411 22559
rect 29546 22556 29552 22568
rect 28399 22528 29552 22556
rect 28399 22525 28411 22528
rect 28353 22519 28411 22525
rect 29546 22516 29552 22528
rect 29604 22516 29610 22568
rect 29914 22516 29920 22568
rect 29972 22556 29978 22568
rect 30300 22556 30328 22587
rect 30374 22584 30380 22636
rect 30432 22624 30438 22636
rect 30469 22627 30527 22633
rect 30469 22624 30481 22627
rect 30432 22596 30481 22624
rect 30432 22584 30438 22596
rect 30469 22593 30481 22596
rect 30515 22593 30527 22627
rect 30469 22587 30527 22593
rect 29972 22528 30328 22556
rect 30484 22556 30512 22587
rect 30650 22584 30656 22636
rect 30708 22624 30714 22636
rect 31846 22624 31852 22636
rect 30708 22596 31852 22624
rect 30708 22584 30714 22596
rect 31846 22584 31852 22596
rect 31904 22584 31910 22636
rect 32306 22584 32312 22636
rect 32364 22584 32370 22636
rect 32416 22633 32444 22664
rect 32858 22652 32864 22704
rect 32916 22692 32922 22704
rect 33137 22695 33195 22701
rect 33137 22692 33149 22695
rect 32916 22664 33149 22692
rect 32916 22652 32922 22664
rect 33137 22661 33149 22664
rect 33183 22661 33195 22695
rect 33137 22655 33195 22661
rect 32401 22627 32459 22633
rect 32401 22593 32413 22627
rect 32447 22593 32459 22627
rect 32401 22587 32459 22593
rect 32674 22584 32680 22636
rect 32732 22584 32738 22636
rect 32950 22584 32956 22636
rect 33008 22584 33014 22636
rect 33042 22584 33048 22636
rect 33100 22624 33106 22636
rect 33244 22624 33272 22732
rect 35161 22695 35219 22701
rect 35161 22692 35173 22695
rect 33428 22664 35173 22692
rect 33318 22633 33324 22636
rect 33100 22596 33272 22624
rect 33301 22627 33324 22633
rect 33100 22584 33106 22596
rect 33301 22593 33313 22627
rect 33376 22624 33382 22636
rect 33428 22624 33456 22664
rect 35161 22661 35173 22664
rect 35207 22661 35219 22695
rect 35161 22655 35219 22661
rect 35805 22695 35863 22701
rect 35805 22661 35817 22695
rect 35851 22692 35863 22695
rect 35851 22664 36768 22692
rect 35851 22661 35863 22664
rect 35805 22655 35863 22661
rect 33376 22596 33456 22624
rect 33301 22587 33324 22593
rect 33318 22584 33324 22587
rect 33376 22584 33382 22596
rect 33778 22584 33784 22636
rect 33836 22624 33842 22636
rect 34885 22627 34943 22633
rect 34885 22624 34897 22627
rect 33836 22596 34897 22624
rect 33836 22584 33842 22596
rect 34885 22593 34897 22596
rect 34931 22593 34943 22627
rect 34885 22587 34943 22593
rect 35069 22627 35127 22633
rect 35069 22593 35081 22627
rect 35115 22593 35127 22627
rect 35069 22587 35127 22593
rect 35253 22627 35311 22633
rect 35253 22593 35265 22627
rect 35299 22624 35311 22627
rect 35618 22624 35624 22636
rect 35299 22596 35624 22624
rect 35299 22593 35311 22596
rect 35253 22587 35311 22593
rect 32030 22556 32036 22568
rect 30484 22528 32036 22556
rect 29972 22516 29978 22528
rect 32030 22516 32036 22528
rect 32088 22516 32094 22568
rect 35084 22556 35112 22587
rect 35618 22584 35624 22596
rect 35676 22584 35682 22636
rect 35820 22556 35848 22655
rect 36538 22584 36544 22636
rect 36596 22584 36602 22636
rect 35084 22528 35848 22556
rect 36633 22559 36691 22565
rect 36633 22525 36645 22559
rect 36679 22525 36691 22559
rect 36740 22556 36768 22664
rect 37568 22633 37596 22732
rect 37752 22732 38301 22760
rect 37752 22704 37780 22732
rect 38289 22729 38301 22732
rect 38335 22760 38347 22763
rect 38378 22760 38384 22772
rect 38335 22732 38384 22760
rect 38335 22729 38347 22732
rect 38289 22723 38347 22729
rect 38378 22720 38384 22732
rect 38436 22720 38442 22772
rect 38473 22763 38531 22769
rect 38473 22729 38485 22763
rect 38519 22729 38531 22763
rect 38473 22723 38531 22729
rect 37734 22652 37740 22704
rect 37792 22652 37798 22704
rect 37829 22695 37887 22701
rect 37829 22661 37841 22695
rect 37875 22692 37887 22695
rect 38102 22692 38108 22704
rect 37875 22664 38108 22692
rect 37875 22661 37887 22664
rect 37829 22655 37887 22661
rect 38102 22652 38108 22664
rect 38160 22652 38166 22704
rect 38194 22652 38200 22704
rect 38252 22692 38258 22704
rect 38488 22692 38516 22723
rect 39114 22720 39120 22772
rect 39172 22720 39178 22772
rect 39942 22760 39948 22772
rect 39224 22732 39948 22760
rect 39224 22704 39252 22732
rect 39942 22720 39948 22732
rect 40000 22720 40006 22772
rect 40218 22720 40224 22772
rect 40276 22760 40282 22772
rect 41230 22760 41236 22772
rect 40276 22732 41236 22760
rect 40276 22720 40282 22732
rect 41230 22720 41236 22732
rect 41288 22760 41294 22772
rect 41288 22732 41414 22760
rect 41288 22720 41294 22732
rect 38252 22664 38516 22692
rect 38252 22652 38258 22664
rect 39206 22652 39212 22704
rect 39264 22652 39270 22704
rect 41386 22692 41414 22732
rect 41506 22720 41512 22772
rect 41564 22760 41570 22772
rect 42058 22760 42064 22772
rect 41564 22732 42064 22760
rect 41564 22720 41570 22732
rect 42058 22720 42064 22732
rect 42116 22760 42122 22772
rect 43349 22763 43407 22769
rect 43349 22760 43361 22763
rect 42116 22732 43361 22760
rect 42116 22720 42122 22732
rect 43349 22729 43361 22732
rect 43395 22729 43407 22763
rect 43349 22723 43407 22729
rect 44174 22720 44180 22772
rect 44232 22760 44238 22772
rect 45186 22760 45192 22772
rect 44232 22732 45192 22760
rect 44232 22720 44238 22732
rect 45186 22720 45192 22732
rect 45244 22720 45250 22772
rect 48222 22720 48228 22772
rect 48280 22760 48286 22772
rect 49053 22763 49111 22769
rect 48280 22732 49004 22760
rect 48280 22720 48286 22732
rect 44358 22692 44364 22704
rect 41386 22664 44364 22692
rect 37553 22627 37611 22633
rect 37553 22593 37565 22627
rect 37599 22593 37611 22627
rect 37553 22587 37611 22593
rect 37921 22627 37979 22633
rect 37921 22593 37933 22627
rect 37967 22624 37979 22627
rect 38286 22624 38292 22636
rect 37967 22596 38292 22624
rect 37967 22593 37979 22596
rect 37921 22587 37979 22593
rect 38286 22584 38292 22596
rect 38344 22584 38350 22636
rect 38381 22627 38439 22633
rect 38381 22593 38393 22627
rect 38427 22593 38439 22627
rect 38381 22587 38439 22593
rect 38396 22556 38424 22587
rect 38746 22584 38752 22636
rect 38804 22624 38810 22636
rect 39301 22627 39359 22633
rect 39301 22624 39313 22627
rect 38804 22596 39313 22624
rect 38804 22584 38810 22596
rect 39301 22593 39313 22596
rect 39347 22593 39359 22627
rect 39301 22587 39359 22593
rect 39574 22584 39580 22636
rect 39632 22584 39638 22636
rect 39669 22627 39727 22633
rect 39669 22593 39681 22627
rect 39715 22624 39727 22627
rect 42334 22624 42340 22636
rect 39715 22596 42340 22624
rect 39715 22593 39727 22596
rect 39669 22587 39727 22593
rect 42334 22584 42340 22596
rect 42392 22624 42398 22636
rect 42429 22627 42487 22633
rect 42429 22624 42441 22627
rect 42392 22596 42441 22624
rect 42392 22584 42398 22596
rect 42429 22593 42441 22596
rect 42475 22593 42487 22627
rect 42429 22587 42487 22593
rect 42610 22584 42616 22636
rect 42668 22584 42674 22636
rect 42702 22584 42708 22636
rect 42760 22584 42766 22636
rect 43640 22633 43668 22664
rect 44358 22652 44364 22664
rect 44416 22652 44422 22704
rect 44634 22652 44640 22704
rect 44692 22692 44698 22704
rect 48130 22692 48136 22704
rect 44692 22664 48136 22692
rect 44692 22652 44698 22664
rect 48130 22652 48136 22664
rect 48188 22652 48194 22704
rect 48240 22664 48912 22692
rect 43625 22627 43683 22633
rect 43625 22593 43637 22627
rect 43671 22593 43683 22627
rect 43625 22587 43683 22593
rect 43809 22627 43867 22633
rect 43809 22593 43821 22627
rect 43855 22624 43867 22627
rect 45002 22624 45008 22636
rect 43855 22596 45008 22624
rect 43855 22593 43867 22596
rect 43809 22587 43867 22593
rect 45002 22584 45008 22596
rect 45060 22584 45066 22636
rect 45738 22584 45744 22636
rect 45796 22624 45802 22636
rect 48240 22633 48268 22664
rect 48225 22627 48283 22633
rect 48225 22624 48237 22627
rect 45796 22596 48237 22624
rect 45796 22584 45802 22596
rect 48225 22593 48237 22596
rect 48271 22593 48283 22627
rect 48225 22587 48283 22593
rect 48314 22584 48320 22636
rect 48372 22624 48378 22636
rect 48590 22633 48596 22636
rect 48409 22627 48467 22633
rect 48409 22624 48421 22627
rect 48372 22596 48421 22624
rect 48372 22584 48378 22596
rect 48409 22593 48421 22596
rect 48455 22593 48467 22627
rect 48409 22587 48467 22593
rect 48557 22627 48596 22633
rect 48557 22593 48569 22627
rect 48557 22587 48596 22593
rect 48590 22584 48596 22587
rect 48648 22584 48654 22636
rect 48884 22633 48912 22664
rect 48685 22627 48743 22633
rect 48685 22593 48697 22627
rect 48731 22593 48743 22627
rect 48685 22587 48743 22593
rect 48777 22627 48835 22633
rect 48777 22593 48789 22627
rect 48823 22593 48835 22627
rect 48777 22587 48835 22593
rect 48874 22627 48932 22633
rect 48874 22593 48886 22627
rect 48920 22593 48932 22627
rect 48976 22624 49004 22732
rect 49053 22729 49065 22763
rect 49099 22729 49111 22763
rect 49053 22723 49111 22729
rect 49068 22692 49096 22723
rect 50614 22720 50620 22772
rect 50672 22760 50678 22772
rect 51169 22763 51227 22769
rect 50672 22732 50844 22760
rect 50672 22720 50678 22732
rect 50816 22701 50844 22732
rect 51169 22729 51181 22763
rect 51215 22760 51227 22763
rect 51721 22763 51779 22769
rect 51215 22732 51304 22760
rect 51215 22729 51227 22732
rect 51169 22723 51227 22729
rect 51276 22701 51304 22732
rect 51721 22729 51733 22763
rect 51767 22760 51779 22763
rect 51767 22732 56272 22760
rect 51767 22729 51779 22732
rect 51721 22723 51779 22729
rect 50801 22695 50859 22701
rect 49068 22664 50568 22692
rect 49605 22627 49663 22633
rect 49605 22624 49617 22627
rect 48976 22596 49617 22624
rect 48874 22587 48932 22593
rect 49605 22593 49617 22596
rect 49651 22593 49663 22627
rect 49605 22587 49663 22593
rect 38654 22556 38660 22568
rect 36740 22528 37872 22556
rect 38396 22528 38660 22556
rect 36633 22519 36691 22525
rect 29779 22491 29837 22497
rect 29779 22457 29791 22491
rect 29825 22488 29837 22491
rect 30098 22488 30104 22500
rect 29825 22460 30104 22488
rect 29825 22457 29837 22460
rect 29779 22451 29837 22457
rect 30098 22448 30104 22460
rect 30156 22488 30162 22500
rect 33042 22488 33048 22500
rect 30156 22460 33048 22488
rect 30156 22448 30162 22460
rect 33042 22448 33048 22460
rect 33100 22448 33106 22500
rect 35437 22491 35495 22497
rect 35437 22457 35449 22491
rect 35483 22488 35495 22491
rect 36648 22488 36676 22519
rect 37844 22500 37872 22528
rect 38654 22516 38660 22528
rect 38712 22516 38718 22568
rect 43162 22516 43168 22568
rect 43220 22516 43226 22568
rect 43530 22516 43536 22568
rect 43588 22516 43594 22568
rect 43717 22559 43775 22565
rect 43717 22525 43729 22559
rect 43763 22556 43775 22559
rect 44266 22556 44272 22568
rect 43763 22528 44272 22556
rect 43763 22525 43775 22528
rect 43717 22519 43775 22525
rect 44266 22516 44272 22528
rect 44324 22516 44330 22568
rect 47210 22516 47216 22568
rect 47268 22556 47274 22568
rect 47946 22556 47952 22568
rect 47268 22528 47952 22556
rect 47268 22516 47274 22528
rect 47946 22516 47952 22528
rect 48004 22516 48010 22568
rect 48700 22556 48728 22587
rect 48056 22528 48728 22556
rect 48792 22556 48820 22587
rect 49510 22556 49516 22568
rect 48792 22528 49516 22556
rect 35483 22460 36676 22488
rect 36909 22491 36967 22497
rect 35483 22457 35495 22460
rect 35437 22451 35495 22457
rect 36909 22457 36921 22491
rect 36955 22488 36967 22491
rect 37366 22488 37372 22500
rect 36955 22460 37372 22488
rect 36955 22457 36967 22460
rect 36909 22451 36967 22457
rect 37366 22448 37372 22460
rect 37424 22448 37430 22500
rect 37826 22448 37832 22500
rect 37884 22448 37890 22500
rect 38105 22491 38163 22497
rect 38105 22457 38117 22491
rect 38151 22488 38163 22491
rect 38749 22491 38807 22497
rect 38749 22488 38761 22491
rect 38151 22460 38761 22488
rect 38151 22457 38163 22460
rect 38105 22451 38163 22457
rect 38749 22457 38761 22460
rect 38795 22457 38807 22491
rect 38749 22451 38807 22457
rect 38841 22491 38899 22497
rect 38841 22457 38853 22491
rect 38887 22488 38899 22491
rect 39853 22491 39911 22497
rect 39853 22488 39865 22491
rect 38887 22460 39865 22488
rect 38887 22457 38899 22460
rect 38841 22451 38899 22457
rect 39853 22457 39865 22460
rect 39899 22457 39911 22491
rect 39853 22451 39911 22457
rect 14424 22392 15424 22420
rect 14424 22380 14430 22392
rect 29914 22380 29920 22432
rect 29972 22380 29978 22432
rect 30190 22380 30196 22432
rect 30248 22420 30254 22432
rect 31110 22420 31116 22432
rect 30248 22392 31116 22420
rect 30248 22380 30254 22392
rect 31110 22380 31116 22392
rect 31168 22380 31174 22432
rect 32125 22423 32183 22429
rect 32125 22389 32137 22423
rect 32171 22420 32183 22423
rect 32398 22420 32404 22432
rect 32171 22392 32404 22420
rect 32171 22389 32183 22392
rect 32125 22383 32183 22389
rect 32398 22380 32404 22392
rect 32456 22380 32462 22432
rect 32582 22380 32588 22432
rect 32640 22380 32646 22432
rect 32674 22380 32680 22432
rect 32732 22420 32738 22432
rect 33778 22420 33784 22432
rect 32732 22392 33784 22420
rect 32732 22380 32738 22392
rect 33778 22380 33784 22392
rect 33836 22380 33842 22432
rect 35618 22380 35624 22432
rect 35676 22380 35682 22432
rect 36722 22380 36728 22432
rect 36780 22380 36786 22432
rect 38657 22423 38715 22429
rect 38657 22389 38669 22423
rect 38703 22420 38715 22423
rect 40218 22420 40224 22432
rect 38703 22392 40224 22420
rect 38703 22389 38715 22392
rect 38657 22383 38715 22389
rect 40218 22380 40224 22392
rect 40276 22380 40282 22432
rect 40494 22380 40500 22432
rect 40552 22420 40558 22432
rect 44910 22420 44916 22432
rect 40552 22392 44916 22420
rect 40552 22380 40558 22392
rect 44910 22380 44916 22392
rect 44968 22420 44974 22432
rect 48056 22429 48084 22528
rect 49510 22516 49516 22528
rect 49568 22516 49574 22568
rect 49620 22556 49648 22587
rect 49694 22584 49700 22636
rect 49752 22584 49758 22636
rect 49786 22584 49792 22636
rect 49844 22624 49850 22636
rect 49973 22627 50031 22633
rect 49844 22596 49889 22624
rect 49844 22584 49850 22596
rect 49973 22593 49985 22627
rect 50019 22593 50031 22627
rect 49973 22587 50031 22593
rect 50065 22627 50123 22633
rect 50065 22593 50077 22627
rect 50111 22593 50123 22627
rect 50065 22587 50123 22593
rect 49988 22556 50016 22587
rect 49620 22528 50016 22556
rect 49786 22488 49792 22500
rect 49160 22460 49792 22488
rect 48041 22423 48099 22429
rect 48041 22420 48053 22423
rect 44968 22392 48053 22420
rect 44968 22380 44974 22392
rect 48041 22389 48053 22392
rect 48087 22389 48099 22423
rect 48041 22383 48099 22389
rect 48590 22380 48596 22432
rect 48648 22420 48654 22432
rect 49160 22429 49188 22460
rect 49786 22448 49792 22460
rect 49844 22448 49850 22500
rect 49145 22423 49203 22429
rect 49145 22420 49157 22423
rect 48648 22392 49157 22420
rect 48648 22380 48654 22392
rect 49145 22389 49157 22392
rect 49191 22389 49203 22423
rect 49145 22383 49203 22389
rect 49421 22423 49479 22429
rect 49421 22389 49433 22423
rect 49467 22420 49479 22423
rect 49510 22420 49516 22432
rect 49467 22392 49516 22420
rect 49467 22389 49479 22392
rect 49421 22383 49479 22389
rect 49510 22380 49516 22392
rect 49568 22380 49574 22432
rect 49896 22420 49924 22528
rect 49970 22448 49976 22500
rect 50028 22488 50034 22500
rect 50080 22488 50108 22587
rect 50154 22584 50160 22636
rect 50212 22633 50218 22636
rect 50540 22633 50568 22664
rect 50801 22661 50813 22695
rect 50847 22661 50859 22695
rect 50801 22655 50859 22661
rect 50893 22695 50951 22701
rect 50893 22661 50905 22695
rect 50939 22692 50951 22695
rect 51261 22695 51319 22701
rect 50939 22664 51212 22692
rect 50939 22661 50951 22664
rect 50893 22655 50951 22661
rect 51184 22636 51212 22664
rect 51261 22661 51273 22695
rect 51307 22661 51319 22695
rect 51261 22655 51319 22661
rect 53006 22652 53012 22704
rect 53064 22652 53070 22704
rect 54478 22692 54484 22704
rect 54234 22664 54484 22692
rect 54478 22652 54484 22664
rect 54536 22652 54542 22704
rect 55398 22652 55404 22704
rect 55456 22652 55462 22704
rect 56042 22652 56048 22704
rect 56100 22652 56106 22704
rect 50212 22624 50220 22633
rect 50525 22627 50583 22633
rect 50212 22596 50257 22624
rect 50212 22587 50220 22596
rect 50525 22593 50537 22627
rect 50571 22593 50583 22627
rect 50525 22587 50583 22593
rect 50673 22627 50731 22633
rect 50673 22593 50685 22627
rect 50719 22624 50731 22627
rect 50982 22624 50988 22636
rect 51040 22633 51046 22636
rect 50719 22593 50752 22624
rect 50948 22596 50988 22624
rect 50673 22587 50752 22593
rect 50212 22584 50218 22587
rect 50724 22556 50752 22587
rect 50982 22584 50988 22596
rect 51040 22587 51048 22633
rect 51040 22584 51046 22587
rect 51166 22584 51172 22636
rect 51224 22584 51230 22636
rect 51276 22596 51488 22624
rect 51276 22556 51304 22596
rect 50724 22528 51304 22556
rect 51350 22516 51356 22568
rect 51408 22516 51414 22568
rect 51460 22556 51488 22596
rect 51534 22584 51540 22636
rect 51592 22584 51598 22636
rect 54846 22584 54852 22636
rect 54904 22584 54910 22636
rect 55122 22584 55128 22636
rect 55180 22584 55186 22636
rect 55217 22627 55275 22633
rect 55217 22593 55229 22627
rect 55263 22593 55275 22627
rect 55217 22587 55275 22593
rect 52638 22556 52644 22568
rect 51460 22528 52644 22556
rect 52638 22516 52644 22528
rect 52696 22516 52702 22568
rect 52730 22516 52736 22568
rect 52788 22516 52794 22568
rect 54864 22556 54892 22584
rect 55232 22556 55260 22587
rect 52840 22528 54892 22556
rect 54956 22528 55260 22556
rect 56060 22556 56088 22652
rect 56244 22633 56272 22732
rect 56870 22720 56876 22772
rect 56928 22720 56934 22772
rect 58526 22720 58532 22772
rect 58584 22760 58590 22772
rect 58621 22763 58679 22769
rect 58621 22760 58633 22763
rect 58584 22732 58633 22760
rect 58584 22720 58590 22732
rect 58621 22729 58633 22732
rect 58667 22729 58679 22763
rect 58621 22723 58679 22729
rect 56229 22627 56287 22633
rect 56229 22593 56241 22627
rect 56275 22593 56287 22627
rect 56229 22587 56287 22593
rect 56318 22584 56324 22636
rect 56376 22624 56382 22636
rect 58544 22633 58572 22720
rect 56413 22627 56471 22633
rect 56413 22624 56425 22627
rect 56376 22596 56425 22624
rect 56376 22584 56382 22596
rect 56413 22593 56425 22596
rect 56459 22593 56471 22627
rect 56413 22587 56471 22593
rect 56505 22627 56563 22633
rect 56505 22593 56517 22627
rect 56551 22593 56563 22627
rect 56505 22587 56563 22593
rect 56597 22627 56655 22633
rect 56597 22593 56609 22627
rect 56643 22624 56655 22627
rect 57885 22627 57943 22633
rect 57885 22624 57897 22627
rect 56643 22596 57897 22624
rect 56643 22593 56655 22596
rect 56597 22587 56655 22593
rect 57885 22593 57897 22596
rect 57931 22593 57943 22627
rect 57885 22587 57943 22593
rect 58529 22627 58587 22633
rect 58529 22593 58541 22627
rect 58575 22593 58587 22627
rect 58529 22587 58587 22593
rect 56520 22556 56548 22587
rect 56060 22528 56548 22556
rect 50028 22460 50108 22488
rect 50341 22491 50399 22497
rect 50028 22448 50034 22460
rect 50341 22457 50353 22491
rect 50387 22488 50399 22491
rect 52656 22488 52684 22516
rect 52840 22488 52868 22528
rect 50387 22460 51304 22488
rect 52656 22460 52868 22488
rect 50387 22457 50399 22460
rect 50341 22451 50399 22457
rect 50154 22420 50160 22432
rect 49896 22392 50160 22420
rect 50154 22380 50160 22392
rect 50212 22380 50218 22432
rect 51276 22429 51304 22460
rect 54110 22448 54116 22500
rect 54168 22488 54174 22500
rect 54665 22491 54723 22497
rect 54665 22488 54677 22491
rect 54168 22460 54677 22488
rect 54168 22448 54174 22460
rect 54665 22457 54677 22460
rect 54711 22488 54723 22491
rect 54956 22488 54984 22528
rect 55214 22488 55220 22500
rect 54711 22460 54984 22488
rect 54711 22457 54723 22460
rect 54665 22451 54723 22457
rect 55186 22448 55220 22488
rect 55272 22448 55278 22500
rect 51261 22423 51319 22429
rect 51261 22389 51273 22423
rect 51307 22389 51319 22423
rect 51261 22383 51319 22389
rect 54478 22380 54484 22432
rect 54536 22380 54542 22432
rect 54941 22423 54999 22429
rect 54941 22389 54953 22423
rect 54987 22420 54999 22423
rect 55186 22420 55214 22448
rect 54987 22392 55214 22420
rect 54987 22389 54999 22392
rect 54941 22383 54999 22389
rect 1104 22330 78844 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 78844 22330
rect 1104 22256 78844 22278
rect 11146 22176 11152 22228
rect 11204 22216 11210 22228
rect 11713 22219 11771 22225
rect 11713 22216 11725 22219
rect 11204 22188 11725 22216
rect 11204 22176 11210 22188
rect 11713 22185 11725 22188
rect 11759 22185 11771 22219
rect 11713 22179 11771 22185
rect 14921 22219 14979 22225
rect 14921 22185 14933 22219
rect 14967 22216 14979 22219
rect 15102 22216 15108 22228
rect 14967 22188 15108 22216
rect 14967 22185 14979 22188
rect 14921 22179 14979 22185
rect 15102 22176 15108 22188
rect 15160 22176 15166 22228
rect 16577 22219 16635 22225
rect 16577 22185 16589 22219
rect 16623 22216 16635 22219
rect 16942 22216 16948 22228
rect 16623 22188 16948 22216
rect 16623 22185 16635 22188
rect 16577 22179 16635 22185
rect 16942 22176 16948 22188
rect 17000 22176 17006 22228
rect 29181 22219 29239 22225
rect 29181 22185 29193 22219
rect 29227 22216 29239 22219
rect 29822 22216 29828 22228
rect 29227 22188 29828 22216
rect 29227 22185 29239 22188
rect 29181 22179 29239 22185
rect 29822 22176 29828 22188
rect 29880 22176 29886 22228
rect 30006 22176 30012 22228
rect 30064 22176 30070 22228
rect 31110 22176 31116 22228
rect 31168 22216 31174 22228
rect 38194 22216 38200 22228
rect 31168 22188 38200 22216
rect 31168 22176 31174 22188
rect 38194 22176 38200 22188
rect 38252 22176 38258 22228
rect 40586 22216 40592 22228
rect 38580 22188 40592 22216
rect 12986 22108 12992 22160
rect 13044 22108 13050 22160
rect 30190 22108 30196 22160
rect 30248 22148 30254 22160
rect 30466 22148 30472 22160
rect 30248 22120 30472 22148
rect 30248 22108 30254 22120
rect 30466 22108 30472 22120
rect 30524 22108 30530 22160
rect 30558 22108 30564 22160
rect 30616 22148 30622 22160
rect 31021 22151 31079 22157
rect 31021 22148 31033 22151
rect 30616 22120 31033 22148
rect 30616 22108 30622 22120
rect 31021 22117 31033 22120
rect 31067 22148 31079 22151
rect 31202 22148 31208 22160
rect 31067 22120 31208 22148
rect 31067 22117 31079 22120
rect 31021 22111 31079 22117
rect 31202 22108 31208 22120
rect 31260 22108 31266 22160
rect 35618 22108 35624 22160
rect 35676 22148 35682 22160
rect 38580 22148 38608 22188
rect 40586 22176 40592 22188
rect 40644 22176 40650 22228
rect 44266 22176 44272 22228
rect 44324 22216 44330 22228
rect 45005 22219 45063 22225
rect 45005 22216 45017 22219
rect 44324 22188 45017 22216
rect 44324 22176 44330 22188
rect 45005 22185 45017 22188
rect 45051 22216 45063 22219
rect 45278 22216 45284 22228
rect 45051 22188 45284 22216
rect 45051 22185 45063 22188
rect 45005 22179 45063 22185
rect 45278 22176 45284 22188
rect 45336 22216 45342 22228
rect 45833 22219 45891 22225
rect 45833 22216 45845 22219
rect 45336 22188 45845 22216
rect 45336 22176 45342 22188
rect 45833 22185 45845 22188
rect 45879 22185 45891 22219
rect 47210 22216 47216 22228
rect 45833 22179 45891 22185
rect 46676 22188 47216 22216
rect 43990 22148 43996 22160
rect 35676 22120 38608 22148
rect 38672 22120 43996 22148
rect 35676 22108 35682 22120
rect 9674 22040 9680 22092
rect 9732 22080 9738 22092
rect 11977 22083 12035 22089
rect 11977 22080 11989 22083
rect 9732 22052 11989 22080
rect 9732 22040 9738 22052
rect 11977 22049 11989 22052
rect 12023 22049 12035 22083
rect 11977 22043 12035 22049
rect 12434 22040 12440 22092
rect 12492 22080 12498 22092
rect 12713 22083 12771 22089
rect 12713 22080 12725 22083
rect 12492 22052 12725 22080
rect 12492 22040 12498 22052
rect 12713 22049 12725 22052
rect 12759 22049 12771 22083
rect 12713 22043 12771 22049
rect 14090 22040 14096 22092
rect 14148 22080 14154 22092
rect 14277 22083 14335 22089
rect 14277 22080 14289 22083
rect 14148 22052 14289 22080
rect 14148 22040 14154 22052
rect 14277 22049 14289 22052
rect 14323 22049 14335 22083
rect 14277 22043 14335 22049
rect 17037 22083 17095 22089
rect 17037 22049 17049 22083
rect 17083 22080 17095 22083
rect 17494 22080 17500 22092
rect 17083 22052 17500 22080
rect 17083 22049 17095 22052
rect 17037 22043 17095 22049
rect 17494 22040 17500 22052
rect 17552 22040 17558 22092
rect 18598 22040 18604 22092
rect 18656 22040 18662 22092
rect 29546 22040 29552 22092
rect 29604 22040 29610 22092
rect 29656 22052 32352 22080
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 22012 1731 22015
rect 7006 22012 7012 22024
rect 1719 21984 7012 22012
rect 1719 21981 1731 21984
rect 1673 21975 1731 21981
rect 7006 21972 7012 21984
rect 7064 21972 7070 22024
rect 16945 22015 17003 22021
rect 16945 21981 16957 22015
rect 16991 22012 17003 22015
rect 17126 22012 17132 22024
rect 16991 21984 17132 22012
rect 16991 21981 17003 21984
rect 16945 21975 17003 21981
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 29365 22015 29423 22021
rect 29365 21981 29377 22015
rect 29411 22012 29423 22015
rect 29656 22012 29684 22052
rect 29411 21984 29684 22012
rect 29733 22015 29791 22021
rect 29411 21981 29423 21984
rect 29365 21975 29423 21981
rect 29733 21981 29745 22015
rect 29779 21981 29791 22015
rect 29733 21975 29791 21981
rect 29825 22015 29883 22021
rect 29825 21981 29837 22015
rect 29871 22012 29883 22015
rect 29914 22012 29920 22024
rect 29871 21984 29920 22012
rect 29871 21981 29883 21984
rect 29825 21975 29883 21981
rect 10042 21904 10048 21956
rect 10100 21944 10106 21956
rect 29748 21944 29776 21975
rect 29914 21972 29920 21984
rect 29972 21972 29978 22024
rect 30098 21972 30104 22024
rect 30156 21972 30162 22024
rect 30282 21972 30288 22024
rect 30340 22012 30346 22024
rect 31110 22012 31116 22024
rect 30340 21984 31116 22012
rect 30340 21972 30346 21984
rect 31110 21972 31116 21984
rect 31168 21972 31174 22024
rect 31389 22015 31447 22021
rect 31389 22012 31401 22015
rect 31220 21984 31401 22012
rect 30650 21944 30656 21956
rect 10100 21916 10534 21944
rect 29748 21916 30656 21944
rect 10100 21904 10106 21916
rect 30650 21904 30656 21916
rect 30708 21904 30714 21956
rect 30742 21904 30748 21956
rect 30800 21944 30806 21956
rect 30837 21947 30895 21953
rect 30837 21944 30849 21947
rect 30800 21916 30849 21944
rect 30800 21904 30806 21916
rect 30837 21913 30849 21916
rect 30883 21944 30895 21947
rect 31220 21944 31248 21984
rect 31389 21981 31401 21984
rect 31435 22012 31447 22015
rect 32033 22015 32091 22021
rect 31435 21984 31754 22012
rect 31435 21981 31447 21984
rect 31389 21975 31447 21981
rect 30883 21916 31248 21944
rect 31726 21944 31754 21984
rect 32033 21981 32045 22015
rect 32079 22012 32091 22015
rect 32122 22012 32128 22024
rect 32079 21984 32128 22012
rect 32079 21981 32091 21984
rect 32033 21975 32091 21981
rect 32122 21972 32128 21984
rect 32180 21972 32186 22024
rect 32324 22012 32352 22052
rect 32398 22040 32404 22092
rect 32456 22040 32462 22092
rect 32508 22052 33732 22080
rect 32508 22012 32536 22052
rect 32324 21984 32536 22012
rect 33704 22012 33732 22052
rect 33778 22040 33784 22092
rect 33836 22089 33842 22092
rect 33836 22083 33885 22089
rect 33836 22049 33839 22083
rect 33873 22049 33885 22083
rect 33836 22043 33885 22049
rect 33836 22040 33842 22043
rect 37182 22040 37188 22092
rect 37240 22080 37246 22092
rect 38672 22080 38700 22120
rect 43990 22108 43996 22120
rect 44048 22108 44054 22160
rect 45186 22108 45192 22160
rect 45244 22148 45250 22160
rect 46676 22157 46704 22188
rect 47210 22176 47216 22188
rect 47268 22176 47274 22228
rect 47394 22176 47400 22228
rect 47452 22216 47458 22228
rect 47452 22188 49648 22216
rect 47452 22176 47458 22188
rect 46661 22151 46719 22157
rect 46661 22148 46673 22151
rect 45244 22120 46673 22148
rect 45244 22108 45250 22120
rect 46661 22117 46673 22120
rect 46707 22117 46719 22151
rect 46661 22111 46719 22117
rect 46750 22108 46756 22160
rect 46808 22148 46814 22160
rect 49620 22148 49648 22188
rect 49694 22176 49700 22228
rect 49752 22216 49758 22228
rect 49789 22219 49847 22225
rect 49789 22216 49801 22219
rect 49752 22188 49801 22216
rect 49752 22176 49758 22188
rect 49789 22185 49801 22188
rect 49835 22185 49847 22219
rect 49789 22179 49847 22185
rect 49970 22176 49976 22228
rect 50028 22216 50034 22228
rect 50154 22216 50160 22228
rect 50028 22188 50160 22216
rect 50028 22176 50034 22188
rect 50154 22176 50160 22188
rect 50212 22176 50218 22228
rect 53190 22176 53196 22228
rect 53248 22216 53254 22228
rect 53285 22219 53343 22225
rect 53285 22216 53297 22219
rect 53248 22188 53297 22216
rect 53248 22176 53254 22188
rect 53285 22185 53297 22188
rect 53331 22185 53343 22219
rect 53285 22179 53343 22185
rect 46808 22120 49188 22148
rect 49620 22120 49740 22148
rect 46808 22108 46814 22120
rect 42518 22080 42524 22092
rect 37240 22052 38700 22080
rect 42260 22052 42524 22080
rect 37240 22040 37246 22052
rect 34606 22012 34612 22024
rect 33704 21984 34612 22012
rect 34606 21972 34612 21984
rect 34664 21972 34670 22024
rect 31938 21944 31944 21956
rect 31726 21916 31944 21944
rect 30883 21913 30895 21916
rect 30837 21907 30895 21913
rect 31938 21904 31944 21916
rect 31996 21904 32002 21956
rect 33410 21904 33416 21956
rect 33468 21944 33474 21956
rect 35986 21944 35992 21956
rect 33468 21916 35992 21944
rect 33468 21904 33474 21916
rect 35986 21904 35992 21916
rect 36044 21944 36050 21956
rect 37185 21947 37243 21953
rect 37185 21944 37197 21947
rect 36044 21916 37197 21944
rect 36044 21904 36050 21916
rect 37185 21913 37197 21916
rect 37231 21913 37243 21947
rect 37185 21907 37243 21913
rect 37553 21947 37611 21953
rect 37553 21913 37565 21947
rect 37599 21944 37611 21947
rect 37829 21947 37887 21953
rect 37829 21944 37841 21947
rect 37599 21916 37841 21944
rect 37599 21913 37611 21916
rect 37553 21907 37611 21913
rect 37829 21913 37841 21916
rect 37875 21944 37887 21947
rect 41598 21944 41604 21956
rect 37875 21916 41604 21944
rect 37875 21913 37887 21916
rect 37829 21907 37887 21913
rect 41598 21904 41604 21916
rect 41656 21904 41662 21956
rect 41782 21904 41788 21956
rect 41840 21904 41846 21956
rect 41966 21904 41972 21956
rect 42024 21944 42030 21956
rect 42150 21944 42156 21956
rect 42024 21916 42156 21944
rect 42024 21904 42030 21916
rect 42150 21904 42156 21916
rect 42208 21904 42214 21956
rect 42260 21953 42288 22052
rect 42518 22040 42524 22052
rect 42576 22080 42582 22092
rect 43070 22080 43076 22092
rect 42576 22052 43076 22080
rect 42576 22040 42582 22052
rect 43070 22040 43076 22052
rect 43128 22080 43134 22092
rect 43898 22080 43904 22092
rect 43128 22052 43904 22080
rect 43128 22040 43134 22052
rect 43898 22040 43904 22052
rect 43956 22080 43962 22092
rect 46569 22083 46627 22089
rect 43956 22052 46244 22080
rect 43956 22040 43962 22052
rect 42610 21972 42616 22024
rect 42668 21972 42674 22024
rect 45204 22021 45232 22052
rect 46032 22021 46060 22052
rect 45189 22015 45247 22021
rect 42904 21984 43208 22012
rect 42245 21947 42303 21953
rect 42245 21913 42257 21947
rect 42291 21913 42303 21947
rect 42245 21907 42303 21913
rect 42521 21947 42579 21953
rect 42521 21913 42533 21947
rect 42567 21944 42579 21947
rect 42794 21944 42800 21956
rect 42567 21916 42800 21944
rect 42567 21913 42579 21916
rect 42521 21907 42579 21913
rect 42794 21904 42800 21916
rect 42852 21904 42858 21956
rect 842 21836 848 21888
rect 900 21876 906 21888
rect 1489 21879 1547 21885
rect 1489 21876 1501 21879
rect 900 21848 1501 21876
rect 900 21836 906 21848
rect 1489 21845 1501 21848
rect 1535 21845 1547 21879
rect 1489 21839 1547 21845
rect 10229 21879 10287 21885
rect 10229 21845 10241 21879
rect 10275 21876 10287 21879
rect 11054 21876 11060 21888
rect 10275 21848 11060 21876
rect 10275 21845 10287 21848
rect 10229 21839 10287 21845
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 13173 21879 13231 21885
rect 13173 21845 13185 21879
rect 13219 21876 13231 21879
rect 13906 21876 13912 21888
rect 13219 21848 13912 21876
rect 13219 21845 13231 21848
rect 13173 21839 13231 21845
rect 13906 21836 13912 21848
rect 13964 21836 13970 21888
rect 29730 21836 29736 21888
rect 29788 21876 29794 21888
rect 34238 21876 34244 21888
rect 29788 21848 34244 21876
rect 29788 21836 29794 21848
rect 34238 21836 34244 21848
rect 34296 21836 34302 21888
rect 37458 21836 37464 21888
rect 37516 21876 37522 21888
rect 37918 21876 37924 21888
rect 37516 21848 37924 21876
rect 37516 21836 37522 21848
rect 37918 21836 37924 21848
rect 37976 21836 37982 21888
rect 38286 21836 38292 21888
rect 38344 21836 38350 21888
rect 38654 21836 38660 21888
rect 38712 21876 38718 21888
rect 39301 21879 39359 21885
rect 39301 21876 39313 21879
rect 38712 21848 39313 21876
rect 38712 21836 38718 21848
rect 39301 21845 39313 21848
rect 39347 21876 39359 21879
rect 39850 21876 39856 21888
rect 39347 21848 39856 21876
rect 39347 21845 39359 21848
rect 39301 21839 39359 21845
rect 39850 21836 39856 21848
rect 39908 21836 39914 21888
rect 42337 21879 42395 21885
rect 42337 21845 42349 21879
rect 42383 21876 42395 21879
rect 42904 21876 42932 21984
rect 42978 21904 42984 21956
rect 43036 21904 43042 21956
rect 43070 21904 43076 21956
rect 43128 21904 43134 21956
rect 43180 21885 43208 21984
rect 45189 21981 45201 22015
rect 45235 21981 45247 22015
rect 45189 21975 45247 21981
rect 45281 22015 45339 22021
rect 45281 21981 45293 22015
rect 45327 21981 45339 22015
rect 45281 21975 45339 21981
rect 46017 22015 46075 22021
rect 46017 21981 46029 22015
rect 46063 21981 46075 22015
rect 46017 21975 46075 21981
rect 46109 22015 46167 22021
rect 46109 21981 46121 22015
rect 46155 21981 46167 22015
rect 46216 22012 46244 22052
rect 46569 22049 46581 22083
rect 46615 22080 46627 22083
rect 46768 22080 46796 22108
rect 46615 22052 46796 22080
rect 46615 22049 46627 22052
rect 46569 22043 46627 22049
rect 47394 22040 47400 22092
rect 47452 22040 47458 22092
rect 49160 22089 49188 22120
rect 49712 22092 49740 22120
rect 49145 22083 49203 22089
rect 49145 22049 49157 22083
rect 49191 22080 49203 22083
rect 49191 22052 49648 22080
rect 49191 22049 49203 22052
rect 49145 22043 49203 22049
rect 49620 22024 49648 22052
rect 49694 22040 49700 22092
rect 49752 22040 49758 22092
rect 49786 22040 49792 22092
rect 49844 22080 49850 22092
rect 50341 22083 50399 22089
rect 50341 22080 50353 22083
rect 49844 22052 50353 22080
rect 49844 22040 49850 22052
rect 50341 22049 50353 22052
rect 50387 22080 50399 22083
rect 50982 22080 50988 22092
rect 50387 22052 50988 22080
rect 50387 22049 50399 22052
rect 50341 22043 50399 22049
rect 50982 22040 50988 22052
rect 51040 22040 51046 22092
rect 52546 22040 52552 22092
rect 52604 22080 52610 22092
rect 52604 22052 52868 22080
rect 52604 22040 52610 22052
rect 46382 22012 46388 22024
rect 46216 21984 46388 22012
rect 46109 21975 46167 21981
rect 43346 21904 43352 21956
rect 43404 21904 43410 21956
rect 43530 21904 43536 21956
rect 43588 21944 43594 21956
rect 43898 21944 43904 21956
rect 43588 21916 43904 21944
rect 43588 21904 43594 21916
rect 43898 21904 43904 21916
rect 43956 21944 43962 21956
rect 45094 21944 45100 21956
rect 43956 21916 45100 21944
rect 43956 21904 43962 21916
rect 45094 21904 45100 21916
rect 45152 21944 45158 21956
rect 45296 21944 45324 21975
rect 45152 21916 45324 21944
rect 45152 21904 45158 21916
rect 45554 21904 45560 21956
rect 45612 21944 45618 21956
rect 45738 21944 45744 21956
rect 45612 21916 45744 21944
rect 45612 21904 45618 21916
rect 45738 21904 45744 21916
rect 45796 21904 45802 21956
rect 42383 21848 42932 21876
rect 43165 21879 43223 21885
rect 42383 21845 42395 21848
rect 42337 21839 42395 21845
rect 43165 21845 43177 21879
rect 43211 21876 43223 21879
rect 44266 21876 44272 21888
rect 43211 21848 44272 21876
rect 43211 21845 43223 21848
rect 43165 21839 43223 21845
rect 44266 21836 44272 21848
rect 44324 21836 44330 21888
rect 46124 21876 46152 21975
rect 46382 21972 46388 21984
rect 46440 22012 46446 22024
rect 46937 22015 46995 22021
rect 46440 21984 46888 22012
rect 46440 21972 46446 21984
rect 46860 21953 46888 21984
rect 46937 21981 46949 22015
rect 46983 22012 46995 22015
rect 47026 22012 47032 22024
rect 46983 21984 47032 22012
rect 46983 21981 46995 21984
rect 46937 21975 46995 21981
rect 47026 21972 47032 21984
rect 47084 21972 47090 22024
rect 49234 21972 49240 22024
rect 49292 21972 49298 22024
rect 49602 21972 49608 22024
rect 49660 21972 49666 22024
rect 52638 21972 52644 22024
rect 52696 22012 52702 22024
rect 52733 22015 52791 22021
rect 52733 22012 52745 22015
rect 52696 21984 52745 22012
rect 52696 21972 52702 21984
rect 52733 21981 52745 21984
rect 52779 21981 52791 22015
rect 52840 22012 52868 22052
rect 52914 22040 52920 22092
rect 52972 22080 52978 22092
rect 54113 22083 54171 22089
rect 54113 22080 54125 22083
rect 52972 22052 54125 22080
rect 52972 22040 52978 22052
rect 54113 22049 54125 22052
rect 54159 22080 54171 22083
rect 56962 22080 56968 22092
rect 54159 22052 56968 22080
rect 54159 22049 54171 22052
rect 54113 22043 54171 22049
rect 56962 22040 56968 22052
rect 57020 22040 57026 22092
rect 53006 22012 53012 22024
rect 52840 21984 53012 22012
rect 52733 21975 52791 21981
rect 53006 21972 53012 21984
rect 53064 21972 53070 22024
rect 53101 22015 53159 22021
rect 53101 21981 53113 22015
rect 53147 22012 53159 22015
rect 54938 22012 54944 22024
rect 53147 21984 54944 22012
rect 53147 21981 53159 21984
rect 53101 21975 53159 21981
rect 54938 21972 54944 21984
rect 54996 21972 55002 22024
rect 46845 21947 46903 21953
rect 46845 21913 46857 21947
rect 46891 21944 46903 21947
rect 47762 21944 47768 21956
rect 46891 21916 47768 21944
rect 46891 21913 46903 21916
rect 46845 21907 46903 21913
rect 47762 21904 47768 21916
rect 47820 21904 47826 21956
rect 48866 21904 48872 21956
rect 48924 21944 48930 21956
rect 48961 21947 49019 21953
rect 48961 21944 48973 21947
rect 48924 21916 48973 21944
rect 48924 21904 48930 21916
rect 48961 21913 48973 21916
rect 49007 21944 49019 21947
rect 49326 21944 49332 21956
rect 49007 21916 49332 21944
rect 49007 21913 49019 21916
rect 48961 21907 49019 21913
rect 49326 21904 49332 21916
rect 49384 21944 49390 21956
rect 49421 21947 49479 21953
rect 49421 21944 49433 21947
rect 49384 21916 49433 21944
rect 49384 21904 49390 21916
rect 49421 21913 49433 21916
rect 49467 21913 49479 21947
rect 49421 21907 49479 21913
rect 49513 21947 49571 21953
rect 49513 21913 49525 21947
rect 49559 21944 49571 21947
rect 52822 21944 52828 21956
rect 49559 21916 52828 21944
rect 49559 21913 49571 21916
rect 49513 21907 49571 21913
rect 52822 21904 52828 21916
rect 52880 21904 52886 21956
rect 52917 21947 52975 21953
rect 52917 21913 52929 21947
rect 52963 21913 52975 21947
rect 52917 21907 52975 21913
rect 46934 21876 46940 21888
rect 46124 21848 46940 21876
rect 46934 21836 46940 21848
rect 46992 21836 46998 21888
rect 48130 21836 48136 21888
rect 48188 21876 48194 21888
rect 49878 21876 49884 21888
rect 48188 21848 49884 21876
rect 48188 21836 48194 21848
rect 49878 21836 49884 21848
rect 49936 21836 49942 21888
rect 50154 21836 50160 21888
rect 50212 21876 50218 21888
rect 50614 21876 50620 21888
rect 50212 21848 50620 21876
rect 50212 21836 50218 21848
rect 50614 21836 50620 21848
rect 50672 21836 50678 21888
rect 52932 21876 52960 21907
rect 53374 21904 53380 21956
rect 53432 21904 53438 21956
rect 53742 21876 53748 21888
rect 52932 21848 53748 21876
rect 53742 21836 53748 21848
rect 53800 21836 53806 21888
rect 1104 21786 78844 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 66314 21786
rect 66366 21734 66378 21786
rect 66430 21734 66442 21786
rect 66494 21734 66506 21786
rect 66558 21734 66570 21786
rect 66622 21734 78844 21786
rect 1104 21712 78844 21734
rect 12434 21632 12440 21684
rect 12492 21632 12498 21684
rect 12636 21644 13584 21672
rect 7742 21604 7748 21616
rect 7576 21576 7748 21604
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 7374 21536 7380 21548
rect 1719 21508 7380 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 7374 21496 7380 21508
rect 7432 21496 7438 21548
rect 7576 21545 7604 21576
rect 7742 21564 7748 21576
rect 7800 21564 7806 21616
rect 9674 21604 9680 21616
rect 9062 21576 9680 21604
rect 9674 21564 9680 21576
rect 9732 21604 9738 21616
rect 10042 21604 10048 21616
rect 9732 21576 10048 21604
rect 9732 21564 9738 21576
rect 10042 21564 10048 21576
rect 10100 21604 10106 21616
rect 12636 21604 12664 21644
rect 10100 21576 12664 21604
rect 10100 21564 10106 21576
rect 13446 21564 13452 21616
rect 13504 21604 13510 21616
rect 13556 21604 13584 21644
rect 29822 21632 29828 21684
rect 29880 21632 29886 21684
rect 30116 21644 30880 21672
rect 13504 21576 13584 21604
rect 13504 21564 13510 21576
rect 13906 21564 13912 21616
rect 13964 21564 13970 21616
rect 29840 21604 29868 21632
rect 30116 21616 30144 21644
rect 30009 21607 30067 21613
rect 30009 21604 30021 21607
rect 29840 21576 30021 21604
rect 30009 21573 30021 21576
rect 30055 21573 30067 21607
rect 30009 21567 30067 21573
rect 30098 21564 30104 21616
rect 30156 21564 30162 21616
rect 30852 21604 30880 21644
rect 31110 21632 31116 21684
rect 31168 21672 31174 21684
rect 31205 21675 31263 21681
rect 31205 21672 31217 21675
rect 31168 21644 31217 21672
rect 31168 21632 31174 21644
rect 31205 21641 31217 21644
rect 31251 21641 31263 21675
rect 38746 21672 38752 21684
rect 31205 21635 31263 21641
rect 31726 21644 38752 21672
rect 31726 21604 31754 21644
rect 38746 21632 38752 21644
rect 38804 21632 38810 21684
rect 49786 21672 49792 21684
rect 45112 21644 49792 21672
rect 30852 21576 31754 21604
rect 33410 21564 33416 21616
rect 33468 21604 33474 21616
rect 37553 21607 37611 21613
rect 33468 21576 34638 21604
rect 33468 21564 33474 21576
rect 37553 21573 37565 21607
rect 37599 21604 37611 21607
rect 39482 21604 39488 21616
rect 37599 21576 38332 21604
rect 39330 21576 39488 21604
rect 37599 21573 37611 21576
rect 37553 21567 37611 21573
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21505 7619 21539
rect 7561 21499 7619 21505
rect 29730 21496 29736 21548
rect 29788 21496 29794 21548
rect 29825 21539 29883 21545
rect 29825 21505 29837 21539
rect 29871 21536 29883 21539
rect 29914 21536 29920 21548
rect 29871 21508 29920 21536
rect 29871 21505 29883 21508
rect 29825 21499 29883 21505
rect 29914 21496 29920 21508
rect 29972 21496 29978 21548
rect 30193 21539 30251 21545
rect 30193 21505 30205 21539
rect 30239 21536 30251 21539
rect 30558 21536 30564 21548
rect 30239 21508 30564 21536
rect 30239 21505 30251 21508
rect 30193 21499 30251 21505
rect 30558 21496 30564 21508
rect 30616 21496 30622 21548
rect 30650 21496 30656 21548
rect 30708 21496 30714 21548
rect 30745 21539 30803 21545
rect 30745 21505 30757 21539
rect 30791 21505 30803 21539
rect 30745 21499 30803 21505
rect 7837 21471 7895 21477
rect 7837 21468 7849 21471
rect 7576 21440 7849 21468
rect 7576 21412 7604 21440
rect 7837 21437 7849 21440
rect 7883 21437 7895 21471
rect 7837 21431 7895 21437
rect 14185 21471 14243 21477
rect 14185 21437 14197 21471
rect 14231 21468 14243 21471
rect 14274 21468 14280 21480
rect 14231 21440 14280 21468
rect 14231 21437 14243 21440
rect 14185 21431 14243 21437
rect 14274 21428 14280 21440
rect 14332 21428 14338 21480
rect 30466 21428 30472 21480
rect 30524 21428 30530 21480
rect 7558 21360 7564 21412
rect 7616 21360 7622 21412
rect 29549 21403 29607 21409
rect 29549 21369 29561 21403
rect 29595 21400 29607 21403
rect 30668 21400 30696 21496
rect 29595 21372 30696 21400
rect 29595 21369 29607 21372
rect 29549 21363 29607 21369
rect 842 21292 848 21344
rect 900 21332 906 21344
rect 1489 21335 1547 21341
rect 1489 21332 1501 21335
rect 900 21304 1501 21332
rect 900 21292 906 21304
rect 1489 21301 1501 21304
rect 1535 21301 1547 21335
rect 1489 21295 1547 21301
rect 8202 21292 8208 21344
rect 8260 21332 8266 21344
rect 9309 21335 9367 21341
rect 9309 21332 9321 21335
rect 8260 21304 9321 21332
rect 8260 21292 8266 21304
rect 9309 21301 9321 21304
rect 9355 21301 9367 21335
rect 9309 21295 9367 21301
rect 30377 21335 30435 21341
rect 30377 21301 30389 21335
rect 30423 21332 30435 21335
rect 30760 21332 30788 21499
rect 31018 21496 31024 21548
rect 31076 21496 31082 21548
rect 31386 21496 31392 21548
rect 31444 21496 31450 21548
rect 32122 21496 32128 21548
rect 32180 21536 32186 21548
rect 33873 21539 33931 21545
rect 33873 21536 33885 21539
rect 32180 21508 33885 21536
rect 32180 21496 32186 21508
rect 33873 21505 33885 21508
rect 33919 21505 33931 21539
rect 33873 21499 33931 21505
rect 37458 21496 37464 21548
rect 37516 21496 37522 21548
rect 37642 21496 37648 21548
rect 37700 21496 37706 21548
rect 37829 21539 37887 21545
rect 37829 21505 37841 21539
rect 37875 21505 37887 21539
rect 37829 21499 37887 21505
rect 34149 21471 34207 21477
rect 34149 21437 34161 21471
rect 34195 21468 34207 21471
rect 34698 21468 34704 21480
rect 34195 21440 34704 21468
rect 34195 21437 34207 21440
rect 34149 21431 34207 21437
rect 34698 21428 34704 21440
rect 34756 21428 34762 21480
rect 35434 21428 35440 21480
rect 35492 21468 35498 21480
rect 35621 21471 35679 21477
rect 35621 21468 35633 21471
rect 35492 21440 35633 21468
rect 35492 21428 35498 21440
rect 35621 21437 35633 21440
rect 35667 21468 35679 21471
rect 36357 21471 36415 21477
rect 36357 21468 36369 21471
rect 35667 21440 36369 21468
rect 35667 21437 35679 21440
rect 35621 21431 35679 21437
rect 36357 21437 36369 21440
rect 36403 21468 36415 21471
rect 37844 21468 37872 21499
rect 36403 21440 37872 21468
rect 36403 21437 36415 21440
rect 36357 21431 36415 21437
rect 30929 21403 30987 21409
rect 30929 21369 30941 21403
rect 30975 21400 30987 21403
rect 30975 21372 31754 21400
rect 30975 21369 30987 21372
rect 30929 21363 30987 21369
rect 30423 21304 30788 21332
rect 30423 21301 30435 21304
rect 30377 21295 30435 21301
rect 30834 21292 30840 21344
rect 30892 21332 30898 21344
rect 31386 21332 31392 21344
rect 30892 21304 31392 21332
rect 30892 21292 30898 21304
rect 31386 21292 31392 21304
rect 31444 21332 31450 21344
rect 31481 21335 31539 21341
rect 31481 21332 31493 21335
rect 31444 21304 31493 21332
rect 31444 21292 31450 21304
rect 31481 21301 31493 21304
rect 31527 21301 31539 21335
rect 31726 21332 31754 21372
rect 35342 21360 35348 21412
rect 35400 21400 35406 21412
rect 35713 21403 35771 21409
rect 35713 21400 35725 21403
rect 35400 21372 35725 21400
rect 35400 21360 35406 21372
rect 35713 21369 35725 21372
rect 35759 21369 35771 21403
rect 35713 21363 35771 21369
rect 34330 21332 34336 21344
rect 31726 21304 34336 21332
rect 31481 21295 31539 21301
rect 34330 21292 34336 21304
rect 34388 21292 34394 21344
rect 37274 21292 37280 21344
rect 37332 21292 37338 21344
rect 37550 21292 37556 21344
rect 37608 21332 37614 21344
rect 37826 21332 37832 21344
rect 37608 21304 37832 21332
rect 37608 21292 37614 21304
rect 37826 21292 37832 21304
rect 37884 21292 37890 21344
rect 38304 21341 38332 21576
rect 39482 21564 39488 21576
rect 39540 21564 39546 21616
rect 39666 21564 39672 21616
rect 39724 21604 39730 21616
rect 39724 21576 40080 21604
rect 39724 21564 39730 21576
rect 40052 21545 40080 21576
rect 42150 21564 42156 21616
rect 42208 21604 42214 21616
rect 45112 21604 45140 21644
rect 49786 21632 49792 21644
rect 49844 21632 49850 21684
rect 50062 21632 50068 21684
rect 50120 21672 50126 21684
rect 50338 21672 50344 21684
rect 50120 21644 50344 21672
rect 50120 21632 50126 21644
rect 50338 21632 50344 21644
rect 50396 21632 50402 21684
rect 51261 21675 51319 21681
rect 51261 21641 51273 21675
rect 51307 21672 51319 21675
rect 51350 21672 51356 21684
rect 51307 21644 51356 21672
rect 51307 21641 51319 21644
rect 51261 21635 51319 21641
rect 51350 21632 51356 21644
rect 51408 21632 51414 21684
rect 53285 21675 53343 21681
rect 53285 21641 53297 21675
rect 53331 21672 53343 21675
rect 53374 21672 53380 21684
rect 53331 21644 53380 21672
rect 53331 21641 53343 21644
rect 53285 21635 53343 21641
rect 53374 21632 53380 21644
rect 53432 21632 53438 21684
rect 54478 21672 54484 21684
rect 53668 21644 54484 21672
rect 42208 21576 45140 21604
rect 45189 21607 45247 21613
rect 42208 21564 42214 21576
rect 45189 21573 45201 21607
rect 45235 21604 45247 21607
rect 45370 21604 45376 21616
rect 45235 21576 45376 21604
rect 45235 21573 45247 21576
rect 45189 21567 45247 21573
rect 45370 21564 45376 21576
rect 45428 21604 45434 21616
rect 45925 21607 45983 21613
rect 45925 21604 45937 21607
rect 45428 21576 45937 21604
rect 45428 21564 45434 21576
rect 45925 21573 45937 21576
rect 45971 21604 45983 21607
rect 46658 21604 46664 21616
rect 45971 21576 46664 21604
rect 45971 21573 45983 21576
rect 45925 21567 45983 21573
rect 46658 21564 46664 21576
rect 46716 21564 46722 21616
rect 50249 21607 50307 21613
rect 46952 21576 47900 21604
rect 46952 21548 46980 21576
rect 40037 21539 40095 21545
rect 40037 21505 40049 21539
rect 40083 21505 40095 21539
rect 40037 21499 40095 21505
rect 45094 21496 45100 21548
rect 45152 21496 45158 21548
rect 45278 21496 45284 21548
rect 45336 21536 45342 21548
rect 45741 21539 45799 21545
rect 45741 21536 45753 21539
rect 45336 21508 45753 21536
rect 45336 21496 45342 21508
rect 45741 21505 45753 21508
rect 45787 21505 45799 21539
rect 45741 21499 45799 21505
rect 46017 21539 46075 21545
rect 46017 21505 46029 21539
rect 46063 21536 46075 21539
rect 46934 21536 46940 21548
rect 46063 21508 46940 21536
rect 46063 21505 46075 21508
rect 46017 21499 46075 21505
rect 46934 21496 46940 21508
rect 46992 21496 46998 21548
rect 47762 21496 47768 21548
rect 47820 21496 47826 21548
rect 47872 21545 47900 21576
rect 50249 21573 50261 21607
rect 50295 21604 50307 21607
rect 50798 21604 50804 21616
rect 50295 21576 50804 21604
rect 50295 21573 50307 21576
rect 50249 21567 50307 21573
rect 50798 21564 50804 21576
rect 50856 21564 50862 21616
rect 52822 21564 52828 21616
rect 52880 21604 52886 21616
rect 53668 21604 53696 21644
rect 54478 21632 54484 21644
rect 54536 21632 54542 21684
rect 52880 21576 53696 21604
rect 52880 21564 52886 21576
rect 53742 21564 53748 21616
rect 53800 21604 53806 21616
rect 54757 21607 54815 21613
rect 54757 21604 54769 21607
rect 53800 21576 54769 21604
rect 53800 21564 53806 21576
rect 54757 21573 54769 21576
rect 54803 21573 54815 21607
rect 54757 21567 54815 21573
rect 55306 21564 55312 21616
rect 55364 21604 55370 21616
rect 55364 21590 55522 21604
rect 55364 21576 55536 21590
rect 55364 21564 55370 21576
rect 47857 21539 47915 21545
rect 47857 21505 47869 21539
rect 47903 21505 47915 21539
rect 47857 21499 47915 21505
rect 49970 21496 49976 21548
rect 50028 21496 50034 21548
rect 50062 21496 50068 21548
rect 50120 21536 50126 21548
rect 50157 21539 50215 21545
rect 50157 21536 50169 21539
rect 50120 21508 50169 21536
rect 50120 21496 50126 21508
rect 50157 21505 50169 21508
rect 50203 21505 50215 21539
rect 50157 21499 50215 21505
rect 50341 21539 50399 21545
rect 50341 21505 50353 21539
rect 50387 21505 50399 21539
rect 50617 21539 50675 21545
rect 50617 21536 50629 21539
rect 50341 21499 50399 21505
rect 50540 21508 50629 21536
rect 39758 21428 39764 21480
rect 39816 21428 39822 21480
rect 44637 21471 44695 21477
rect 44637 21437 44649 21471
rect 44683 21468 44695 21471
rect 44910 21468 44916 21480
rect 44683 21440 44916 21468
rect 44683 21437 44695 21440
rect 44637 21431 44695 21437
rect 44910 21428 44916 21440
rect 44968 21428 44974 21480
rect 50356 21468 50384 21499
rect 49620 21440 50384 21468
rect 40586 21360 40592 21412
rect 40644 21400 40650 21412
rect 42610 21400 42616 21412
rect 40644 21372 42616 21400
rect 40644 21360 40650 21372
rect 42610 21360 42616 21372
rect 42668 21400 42674 21412
rect 46106 21400 46112 21412
rect 42668 21372 46112 21400
rect 42668 21360 42674 21372
rect 46106 21360 46112 21372
rect 46164 21360 46170 21412
rect 46216 21372 48176 21400
rect 46216 21344 46244 21372
rect 38289 21335 38347 21341
rect 38289 21301 38301 21335
rect 38335 21332 38347 21335
rect 38654 21332 38660 21344
rect 38335 21304 38660 21332
rect 38335 21301 38347 21304
rect 38289 21295 38347 21301
rect 38654 21292 38660 21304
rect 38712 21292 38718 21344
rect 46198 21292 46204 21344
rect 46256 21292 46262 21344
rect 47394 21292 47400 21344
rect 47452 21332 47458 21344
rect 47581 21335 47639 21341
rect 47581 21332 47593 21335
rect 47452 21304 47593 21332
rect 47452 21292 47458 21304
rect 47581 21301 47593 21304
rect 47627 21301 47639 21335
rect 47581 21295 47639 21301
rect 48038 21292 48044 21344
rect 48096 21292 48102 21344
rect 48148 21332 48176 21372
rect 49620 21332 49648 21440
rect 49694 21360 49700 21412
rect 49752 21400 49758 21412
rect 50062 21400 50068 21412
rect 49752 21372 50068 21400
rect 49752 21360 49758 21372
rect 50062 21360 50068 21372
rect 50120 21360 50126 21412
rect 50540 21409 50568 21508
rect 50617 21505 50629 21508
rect 50663 21505 50675 21539
rect 50617 21499 50675 21505
rect 50710 21539 50768 21545
rect 50710 21505 50722 21539
rect 50756 21505 50768 21539
rect 50710 21499 50768 21505
rect 50525 21403 50583 21409
rect 50525 21369 50537 21403
rect 50571 21369 50583 21403
rect 50525 21363 50583 21369
rect 49789 21335 49847 21341
rect 49789 21332 49801 21335
rect 48148 21304 49801 21332
rect 49789 21301 49801 21304
rect 49835 21301 49847 21335
rect 49789 21295 49847 21301
rect 50430 21292 50436 21344
rect 50488 21332 50494 21344
rect 50724 21332 50752 21499
rect 50890 21496 50896 21548
rect 50948 21496 50954 21548
rect 51166 21545 51172 21548
rect 50985 21539 51043 21545
rect 50985 21505 50997 21539
rect 51031 21505 51043 21539
rect 50985 21499 51043 21505
rect 51123 21539 51172 21545
rect 51123 21505 51135 21539
rect 51169 21505 51172 21539
rect 51123 21499 51172 21505
rect 51000 21468 51028 21499
rect 51166 21496 51172 21499
rect 51224 21496 51230 21548
rect 54478 21496 54484 21548
rect 54536 21536 54542 21548
rect 54573 21539 54631 21545
rect 54573 21536 54585 21539
rect 54536 21508 54585 21536
rect 54536 21496 54542 21508
rect 54573 21505 54585 21508
rect 54619 21505 54631 21539
rect 54573 21499 54631 21505
rect 54846 21496 54852 21548
rect 54904 21496 54910 21548
rect 54938 21496 54944 21548
rect 54996 21496 55002 21548
rect 52178 21468 52184 21480
rect 51000 21440 52184 21468
rect 52178 21428 52184 21440
rect 52236 21428 52242 21480
rect 55508 21468 55536 21576
rect 56962 21496 56968 21548
rect 57020 21496 57026 21548
rect 56226 21468 56232 21480
rect 55508 21440 56232 21468
rect 56226 21428 56232 21440
rect 56284 21428 56290 21480
rect 56594 21428 56600 21480
rect 56652 21468 56658 21480
rect 56689 21471 56747 21477
rect 56689 21468 56701 21471
rect 56652 21440 56701 21468
rect 56652 21428 56658 21440
rect 56689 21437 56701 21440
rect 56735 21437 56747 21471
rect 56689 21431 56747 21437
rect 51626 21360 51632 21412
rect 51684 21400 51690 21412
rect 52362 21400 52368 21412
rect 51684 21372 52368 21400
rect 51684 21360 51690 21372
rect 52362 21360 52368 21372
rect 52420 21400 52426 21412
rect 52914 21400 52920 21412
rect 52420 21372 52920 21400
rect 52420 21360 52426 21372
rect 52914 21360 52920 21372
rect 52972 21400 52978 21412
rect 55490 21400 55496 21412
rect 52972 21372 55496 21400
rect 52972 21360 52978 21372
rect 55490 21360 55496 21372
rect 55548 21360 55554 21412
rect 54202 21332 54208 21344
rect 50488 21304 54208 21332
rect 50488 21292 50494 21304
rect 54202 21292 54208 21304
rect 54260 21292 54266 21344
rect 55122 21292 55128 21344
rect 55180 21292 55186 21344
rect 55214 21292 55220 21344
rect 55272 21292 55278 21344
rect 1104 21242 78844 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 78844 21242
rect 1104 21168 78844 21190
rect 7558 21088 7564 21140
rect 7616 21088 7622 21140
rect 14737 21131 14795 21137
rect 14737 21097 14749 21131
rect 14783 21128 14795 21131
rect 14918 21128 14924 21140
rect 14783 21100 14924 21128
rect 14783 21097 14795 21100
rect 14737 21091 14795 21097
rect 7926 21060 7932 21072
rect 6886 21032 7932 21060
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 6886 20924 6914 21032
rect 7926 21020 7932 21032
rect 7984 21020 7990 21072
rect 7006 20952 7012 21004
rect 7064 20992 7070 21004
rect 8113 20995 8171 21001
rect 8113 20992 8125 20995
rect 7064 20964 8125 20992
rect 7064 20952 7070 20964
rect 8113 20961 8125 20964
rect 8159 20992 8171 20995
rect 8202 20992 8208 21004
rect 8159 20964 8208 20992
rect 8159 20961 8171 20964
rect 8113 20955 8171 20961
rect 8202 20952 8208 20964
rect 8260 20992 8266 21004
rect 9769 20995 9827 21001
rect 9769 20992 9781 20995
rect 8260 20964 9781 20992
rect 8260 20952 8266 20964
rect 9769 20961 9781 20964
rect 9815 20961 9827 20995
rect 12986 20992 12992 21004
rect 9769 20955 9827 20961
rect 11348 20964 12992 20992
rect 1719 20896 6914 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 7098 20884 7104 20936
rect 7156 20884 7162 20936
rect 11348 20933 11376 20964
rect 12986 20952 12992 20964
rect 13044 20952 13050 21004
rect 7285 20927 7343 20933
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 8389 20927 8447 20933
rect 8389 20924 8401 20927
rect 7331 20896 8401 20924
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 8389 20893 8401 20896
rect 8435 20893 8447 20927
rect 8389 20887 8447 20893
rect 11333 20927 11391 20933
rect 11333 20893 11345 20927
rect 11379 20893 11391 20927
rect 11333 20887 11391 20893
rect 11514 20884 11520 20936
rect 11572 20884 11578 20936
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20924 14519 20927
rect 14752 20924 14780 21091
rect 14918 21088 14924 21100
rect 14976 21088 14982 21140
rect 31938 21088 31944 21140
rect 31996 21128 32002 21140
rect 34514 21128 34520 21140
rect 31996 21100 34520 21128
rect 31996 21088 32002 21100
rect 34514 21088 34520 21100
rect 34572 21128 34578 21140
rect 34790 21128 34796 21140
rect 34572 21100 34796 21128
rect 34572 21088 34578 21100
rect 34790 21088 34796 21100
rect 34848 21088 34854 21140
rect 37366 21088 37372 21140
rect 37424 21128 37430 21140
rect 39669 21131 39727 21137
rect 37424 21100 38332 21128
rect 37424 21088 37430 21100
rect 38304 21072 38332 21100
rect 39669 21097 39681 21131
rect 39715 21128 39727 21131
rect 39758 21128 39764 21140
rect 39715 21100 39764 21128
rect 39715 21097 39727 21100
rect 39669 21091 39727 21097
rect 39758 21088 39764 21100
rect 39816 21088 39822 21140
rect 39850 21088 39856 21140
rect 39908 21128 39914 21140
rect 39908 21100 41414 21128
rect 39908 21088 39914 21100
rect 38286 21020 38292 21072
rect 38344 21060 38350 21072
rect 38344 21032 39344 21060
rect 38344 21020 38350 21032
rect 29917 20995 29975 21001
rect 29917 20961 29929 20995
rect 29963 20992 29975 20995
rect 30466 20992 30472 21004
rect 29963 20964 30472 20992
rect 29963 20961 29975 20964
rect 29917 20955 29975 20961
rect 30466 20952 30472 20964
rect 30524 20952 30530 21004
rect 37458 20992 37464 21004
rect 35268 20964 37464 20992
rect 14507 20896 14780 20924
rect 14507 20893 14519 20896
rect 14461 20887 14519 20893
rect 29546 20884 29552 20936
rect 29604 20884 29610 20936
rect 34514 20884 34520 20936
rect 34572 20924 34578 20936
rect 35268 20933 35296 20964
rect 37458 20952 37464 20964
rect 37516 20952 37522 21004
rect 37737 20995 37795 21001
rect 37737 20961 37749 20995
rect 37783 20992 37795 20995
rect 38562 20992 38568 21004
rect 37783 20964 38568 20992
rect 37783 20961 37795 20964
rect 37737 20955 37795 20961
rect 38562 20952 38568 20964
rect 38620 20952 38626 21004
rect 39206 20952 39212 21004
rect 39264 20952 39270 21004
rect 39316 20992 39344 21032
rect 39482 21020 39488 21072
rect 39540 21060 39546 21072
rect 41386 21060 41414 21100
rect 41782 21088 41788 21140
rect 41840 21128 41846 21140
rect 41840 21100 46060 21128
rect 41840 21088 41846 21100
rect 45554 21060 45560 21072
rect 39540 21032 39988 21060
rect 41386 21032 45560 21060
rect 39540 21020 39546 21032
rect 39316 20964 39620 20992
rect 34885 20927 34943 20933
rect 34885 20924 34897 20927
rect 34572 20896 34897 20924
rect 34572 20884 34578 20896
rect 34885 20893 34897 20896
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 35253 20927 35311 20933
rect 35253 20893 35265 20927
rect 35299 20893 35311 20927
rect 35253 20887 35311 20893
rect 35986 20884 35992 20936
rect 36044 20924 36050 20936
rect 38473 20927 38531 20933
rect 36044 20896 36386 20924
rect 36044 20884 36050 20896
rect 38473 20893 38485 20927
rect 38519 20924 38531 20927
rect 38654 20924 38660 20936
rect 38519 20896 38660 20924
rect 38519 20893 38531 20896
rect 38473 20887 38531 20893
rect 38654 20884 38660 20896
rect 38712 20924 38718 20936
rect 38930 20924 38936 20936
rect 38712 20896 38936 20924
rect 38712 20884 38718 20896
rect 38930 20884 38936 20896
rect 38988 20884 38994 20936
rect 39025 20927 39083 20933
rect 39025 20893 39037 20927
rect 39071 20924 39083 20927
rect 39117 20927 39175 20933
rect 39117 20924 39129 20927
rect 39071 20896 39129 20924
rect 39071 20893 39083 20896
rect 39025 20887 39083 20893
rect 39117 20893 39129 20896
rect 39163 20893 39175 20927
rect 39117 20887 39175 20893
rect 39390 20884 39396 20936
rect 39448 20884 39454 20936
rect 39485 20927 39543 20933
rect 39485 20893 39497 20927
rect 39531 20893 39543 20927
rect 39485 20887 39543 20893
rect 7116 20856 7144 20884
rect 8021 20859 8079 20865
rect 8021 20856 8033 20859
rect 7116 20828 8033 20856
rect 8021 20825 8033 20828
rect 8067 20825 8079 20859
rect 8021 20819 8079 20825
rect 8570 20816 8576 20868
rect 8628 20816 8634 20868
rect 8757 20859 8815 20865
rect 8757 20825 8769 20859
rect 8803 20856 8815 20859
rect 30282 20856 30288 20868
rect 8803 20828 10732 20856
rect 8803 20825 8815 20828
rect 8757 20819 8815 20825
rect 1486 20748 1492 20800
rect 1544 20748 1550 20800
rect 7466 20748 7472 20800
rect 7524 20748 7530 20800
rect 7742 20748 7748 20800
rect 7800 20788 7806 20800
rect 7929 20791 7987 20797
rect 7929 20788 7941 20791
rect 7800 20760 7941 20788
rect 7800 20748 7806 20760
rect 7929 20757 7941 20760
rect 7975 20788 7987 20791
rect 8772 20788 8800 20819
rect 10704 20800 10732 20828
rect 30208 20828 30288 20856
rect 7975 20760 8800 20788
rect 10413 20791 10471 20797
rect 7975 20757 7987 20760
rect 7929 20751 7987 20757
rect 10413 20757 10425 20791
rect 10459 20788 10471 20791
rect 10594 20788 10600 20800
rect 10459 20760 10600 20788
rect 10459 20757 10471 20760
rect 10413 20751 10471 20757
rect 10594 20748 10600 20760
rect 10652 20748 10658 20800
rect 10686 20748 10692 20800
rect 10744 20788 10750 20800
rect 11425 20791 11483 20797
rect 11425 20788 11437 20791
rect 10744 20760 11437 20788
rect 10744 20748 10750 20760
rect 11425 20757 11437 20760
rect 11471 20757 11483 20791
rect 11425 20751 11483 20757
rect 13538 20748 13544 20800
rect 13596 20788 13602 20800
rect 14185 20791 14243 20797
rect 14185 20788 14197 20791
rect 13596 20760 14197 20788
rect 13596 20748 13602 20760
rect 14185 20757 14197 20760
rect 14231 20757 14243 20791
rect 30208 20788 30236 20828
rect 30282 20816 30288 20828
rect 30340 20816 30346 20868
rect 31481 20859 31539 20865
rect 31481 20856 31493 20859
rect 31036 20828 31493 20856
rect 31036 20788 31064 20828
rect 31481 20825 31493 20828
rect 31527 20825 31539 20859
rect 31481 20819 31539 20825
rect 34606 20816 34612 20868
rect 34664 20856 34670 20868
rect 35069 20859 35127 20865
rect 35069 20856 35081 20859
rect 34664 20828 35081 20856
rect 34664 20816 34670 20828
rect 35069 20825 35081 20828
rect 35115 20825 35127 20859
rect 35069 20819 35127 20825
rect 35161 20859 35219 20865
rect 35161 20825 35173 20859
rect 35207 20856 35219 20859
rect 35207 20828 36032 20856
rect 35207 20825 35219 20828
rect 35161 20819 35219 20825
rect 30208 20760 31064 20788
rect 14185 20751 14243 20757
rect 31110 20748 31116 20800
rect 31168 20788 31174 20800
rect 31343 20791 31401 20797
rect 31343 20788 31355 20791
rect 31168 20760 31355 20788
rect 31168 20748 31174 20760
rect 31343 20757 31355 20760
rect 31389 20757 31401 20791
rect 31343 20751 31401 20757
rect 34974 20748 34980 20800
rect 35032 20788 35038 20800
rect 36004 20797 36032 20828
rect 37458 20816 37464 20868
rect 37516 20816 37522 20868
rect 35437 20791 35495 20797
rect 35437 20788 35449 20791
rect 35032 20760 35449 20788
rect 35032 20748 35038 20760
rect 35437 20757 35449 20760
rect 35483 20757 35495 20791
rect 35437 20751 35495 20757
rect 35989 20791 36047 20797
rect 35989 20757 36001 20791
rect 36035 20788 36047 20791
rect 36170 20788 36176 20800
rect 36035 20760 36176 20788
rect 36035 20757 36047 20760
rect 35989 20751 36047 20757
rect 36170 20748 36176 20760
rect 36228 20748 36234 20800
rect 36630 20748 36636 20800
rect 36688 20788 36694 20800
rect 39500 20788 39528 20887
rect 36688 20760 39528 20788
rect 39592 20788 39620 20964
rect 39666 20952 39672 21004
rect 39724 20992 39730 21004
rect 39853 20995 39911 21001
rect 39853 20992 39865 20995
rect 39724 20964 39865 20992
rect 39724 20952 39730 20964
rect 39853 20961 39865 20964
rect 39899 20961 39911 20995
rect 39960 20992 39988 21032
rect 45554 21020 45560 21032
rect 45612 21020 45618 21072
rect 45370 20992 45376 21004
rect 39960 20964 41184 20992
rect 39853 20955 39911 20961
rect 41156 20868 41184 20964
rect 42628 20964 45376 20992
rect 41966 20884 41972 20936
rect 42024 20924 42030 20936
rect 42628 20933 42656 20964
rect 42613 20927 42671 20933
rect 42024 20896 42564 20924
rect 42024 20884 42030 20896
rect 42536 20868 42564 20896
rect 42613 20893 42625 20927
rect 42659 20893 42671 20927
rect 42613 20887 42671 20893
rect 42978 20884 42984 20936
rect 43036 20924 43042 20936
rect 44376 20933 44404 20964
rect 45370 20952 45376 20964
rect 45428 20952 45434 21004
rect 46032 20992 46060 21100
rect 46106 21088 46112 21140
rect 46164 21128 46170 21140
rect 50525 21131 50583 21137
rect 50525 21128 50537 21131
rect 46164 21100 50537 21128
rect 46164 21088 46170 21100
rect 50525 21097 50537 21100
rect 50571 21128 50583 21131
rect 50798 21128 50804 21140
rect 50571 21100 50804 21128
rect 50571 21097 50583 21100
rect 50525 21091 50583 21097
rect 50798 21088 50804 21100
rect 50856 21088 50862 21140
rect 51077 21131 51135 21137
rect 51077 21097 51089 21131
rect 51123 21128 51135 21131
rect 53193 21131 53251 21137
rect 53193 21128 53205 21131
rect 51123 21100 53205 21128
rect 51123 21097 51135 21100
rect 51077 21091 51135 21097
rect 53193 21097 53205 21100
rect 53239 21128 53251 21131
rect 53650 21128 53656 21140
rect 53239 21100 53656 21128
rect 53239 21097 53251 21100
rect 53193 21091 53251 21097
rect 53650 21088 53656 21100
rect 53708 21088 53714 21140
rect 54938 21088 54944 21140
rect 54996 21128 55002 21140
rect 56137 21131 56195 21137
rect 56137 21128 56149 21131
rect 54996 21100 56149 21128
rect 54996 21088 55002 21100
rect 56137 21097 56149 21100
rect 56183 21097 56195 21131
rect 56137 21091 56195 21097
rect 56594 21088 56600 21140
rect 56652 21088 56658 21140
rect 47118 21020 47124 21072
rect 47176 21060 47182 21072
rect 50246 21060 50252 21072
rect 47176 21032 50252 21060
rect 47176 21020 47182 21032
rect 50246 21020 50252 21032
rect 50304 21020 50310 21072
rect 50341 21063 50399 21069
rect 50341 21029 50353 21063
rect 50387 21060 50399 21063
rect 50890 21060 50896 21072
rect 50387 21032 50896 21060
rect 50387 21029 50399 21032
rect 50341 21023 50399 21029
rect 50890 21020 50896 21032
rect 50948 21060 50954 21072
rect 51534 21060 51540 21072
rect 50948 21032 51540 21060
rect 50948 21020 50954 21032
rect 51534 21020 51540 21032
rect 51592 21020 51598 21072
rect 53006 21020 53012 21072
rect 53064 21060 53070 21072
rect 53064 21032 54984 21060
rect 53064 21020 53070 21032
rect 48406 20992 48412 21004
rect 46032 20964 48412 20992
rect 48406 20952 48412 20964
rect 48464 20952 48470 21004
rect 48590 20952 48596 21004
rect 48648 20992 48654 21004
rect 50522 20992 50528 21004
rect 48648 20964 49096 20992
rect 48648 20952 48654 20964
rect 44361 20927 44419 20933
rect 43036 20896 44220 20924
rect 43036 20884 43042 20896
rect 40126 20816 40132 20868
rect 40184 20816 40190 20868
rect 41138 20816 41144 20868
rect 41196 20816 41202 20868
rect 42150 20856 42156 20868
rect 41432 20828 42156 20856
rect 41432 20788 41460 20828
rect 42150 20816 42156 20828
rect 42208 20816 42214 20868
rect 42518 20816 42524 20868
rect 42576 20816 42582 20868
rect 42794 20816 42800 20868
rect 42852 20856 42858 20868
rect 42889 20859 42947 20865
rect 42889 20856 42901 20859
rect 42852 20828 42901 20856
rect 42852 20816 42858 20828
rect 42889 20825 42901 20828
rect 42935 20856 42947 20859
rect 43346 20856 43352 20868
rect 42935 20828 43352 20856
rect 42935 20825 42947 20828
rect 42889 20819 42947 20825
rect 43346 20816 43352 20828
rect 43404 20856 43410 20868
rect 44082 20856 44088 20868
rect 43404 20828 44088 20856
rect 43404 20816 43410 20828
rect 44082 20816 44088 20828
rect 44140 20816 44146 20868
rect 44192 20856 44220 20896
rect 44361 20893 44373 20927
rect 44407 20893 44419 20927
rect 44361 20887 44419 20893
rect 45005 20927 45063 20933
rect 45005 20893 45017 20927
rect 45051 20924 45063 20927
rect 45186 20924 45192 20936
rect 45051 20896 45192 20924
rect 45051 20893 45063 20896
rect 45005 20887 45063 20893
rect 45186 20884 45192 20896
rect 45244 20884 45250 20936
rect 45554 20884 45560 20936
rect 45612 20924 45618 20936
rect 46750 20924 46756 20936
rect 45612 20896 46756 20924
rect 45612 20884 45618 20896
rect 46750 20884 46756 20896
rect 46808 20884 46814 20936
rect 49068 20933 49096 20964
rect 49160 20964 50528 20992
rect 49160 20933 49188 20964
rect 50522 20952 50528 20964
rect 50580 20952 50586 21004
rect 51626 20992 51632 21004
rect 50816 20964 51632 20992
rect 48961 20927 49019 20933
rect 48961 20893 48973 20927
rect 49007 20893 49019 20927
rect 48961 20887 49019 20893
rect 49053 20927 49111 20933
rect 49053 20893 49065 20927
rect 49099 20893 49111 20927
rect 49053 20887 49111 20893
rect 49145 20927 49203 20933
rect 49145 20893 49157 20927
rect 49191 20893 49203 20927
rect 49145 20887 49203 20893
rect 49329 20927 49387 20933
rect 49329 20893 49341 20927
rect 49375 20924 49387 20927
rect 49970 20924 49976 20936
rect 49375 20896 49976 20924
rect 49375 20893 49387 20896
rect 49329 20887 49387 20893
rect 44453 20859 44511 20865
rect 44453 20856 44465 20859
rect 44192 20828 44465 20856
rect 44453 20825 44465 20828
rect 44499 20856 44511 20859
rect 44542 20856 44548 20868
rect 44499 20828 44548 20856
rect 44499 20825 44511 20828
rect 44453 20819 44511 20825
rect 44542 20816 44548 20828
rect 44600 20816 44606 20868
rect 44726 20816 44732 20868
rect 44784 20856 44790 20868
rect 44821 20859 44879 20865
rect 44821 20856 44833 20859
rect 44784 20828 44833 20856
rect 44784 20816 44790 20828
rect 44821 20825 44833 20828
rect 44867 20856 44879 20859
rect 47118 20856 47124 20868
rect 44867 20828 47124 20856
rect 44867 20825 44879 20828
rect 44821 20819 44879 20825
rect 47118 20816 47124 20828
rect 47176 20816 47182 20868
rect 39592 20760 41460 20788
rect 36688 20748 36694 20760
rect 41506 20748 41512 20800
rect 41564 20788 41570 20800
rect 41601 20791 41659 20797
rect 41601 20788 41613 20791
rect 41564 20760 41613 20788
rect 41564 20748 41570 20760
rect 41601 20757 41613 20760
rect 41647 20757 41659 20791
rect 41601 20751 41659 20757
rect 42702 20748 42708 20800
rect 42760 20788 42766 20800
rect 44266 20788 44272 20800
rect 42760 20760 44272 20788
rect 42760 20748 42766 20760
rect 44266 20748 44272 20760
rect 44324 20788 44330 20800
rect 45186 20788 45192 20800
rect 44324 20760 45192 20788
rect 44324 20748 44330 20760
rect 45186 20748 45192 20760
rect 45244 20748 45250 20800
rect 48590 20748 48596 20800
rect 48648 20748 48654 20800
rect 48777 20791 48835 20797
rect 48777 20757 48789 20791
rect 48823 20788 48835 20791
rect 48866 20788 48872 20800
rect 48823 20760 48872 20788
rect 48823 20757 48835 20760
rect 48777 20751 48835 20757
rect 48866 20748 48872 20760
rect 48924 20748 48930 20800
rect 48976 20788 49004 20887
rect 49970 20884 49976 20896
rect 50028 20884 50034 20936
rect 50816 20933 50844 20964
rect 51626 20952 51632 20964
rect 51684 20952 51690 21004
rect 52270 20992 52276 21004
rect 51828 20964 52276 20992
rect 50801 20927 50859 20933
rect 50801 20893 50813 20927
rect 50847 20893 50859 20927
rect 50801 20887 50859 20893
rect 50890 20884 50896 20936
rect 50948 20884 50954 20936
rect 51169 20927 51227 20933
rect 51169 20893 51181 20927
rect 51215 20924 51227 20927
rect 51721 20927 51779 20933
rect 51721 20924 51733 20927
rect 51215 20896 51733 20924
rect 51215 20893 51227 20896
rect 51169 20887 51227 20893
rect 51721 20893 51733 20896
rect 51767 20893 51779 20927
rect 51721 20887 51779 20893
rect 49988 20856 50016 20884
rect 51828 20856 51856 20964
rect 52270 20952 52276 20964
rect 52328 20952 52334 21004
rect 52914 20884 52920 20936
rect 52972 20884 52978 20936
rect 53009 20927 53067 20933
rect 53009 20893 53021 20927
rect 53055 20893 53067 20927
rect 53009 20887 53067 20893
rect 53285 20927 53343 20933
rect 53285 20893 53297 20927
rect 53331 20924 53343 20927
rect 53653 20927 53711 20933
rect 53653 20924 53665 20927
rect 53331 20896 53665 20924
rect 53331 20893 53343 20896
rect 53285 20887 53343 20893
rect 53653 20893 53665 20896
rect 53699 20893 53711 20927
rect 54128 20924 54156 21032
rect 54202 20952 54208 21004
rect 54260 20992 54266 21004
rect 54956 20992 54984 21032
rect 55122 21020 55128 21072
rect 55180 21060 55186 21072
rect 55180 21032 56364 21060
rect 55180 21020 55186 21032
rect 55214 20992 55220 21004
rect 54260 20964 54708 20992
rect 54956 20964 55220 20992
rect 54260 20952 54266 20964
rect 54680 20933 54708 20964
rect 55214 20952 55220 20964
rect 55272 20992 55278 21004
rect 55309 20995 55367 21001
rect 55309 20992 55321 20995
rect 55272 20964 55321 20992
rect 55272 20952 55278 20964
rect 55309 20961 55321 20964
rect 55355 20961 55367 20995
rect 55309 20955 55367 20961
rect 56336 20933 56364 21032
rect 54389 20927 54447 20933
rect 54389 20924 54401 20927
rect 54128 20896 54401 20924
rect 53653 20887 53711 20893
rect 54389 20893 54401 20896
rect 54435 20893 54447 20927
rect 54389 20887 54447 20893
rect 54665 20927 54723 20933
rect 54665 20893 54677 20927
rect 54711 20893 54723 20927
rect 54665 20887 54723 20893
rect 54757 20927 54815 20933
rect 54757 20893 54769 20927
rect 54803 20893 54815 20927
rect 54757 20887 54815 20893
rect 55953 20927 56011 20933
rect 55953 20893 55965 20927
rect 55999 20924 56011 20927
rect 56045 20927 56103 20933
rect 56045 20924 56057 20927
rect 55999 20896 56057 20924
rect 55999 20893 56011 20896
rect 55953 20887 56011 20893
rect 56045 20893 56057 20896
rect 56091 20893 56103 20927
rect 56045 20887 56103 20893
rect 56321 20927 56379 20933
rect 56321 20893 56333 20927
rect 56367 20893 56379 20927
rect 56321 20887 56379 20893
rect 56413 20927 56471 20933
rect 56413 20893 56425 20927
rect 56459 20893 56471 20927
rect 56413 20887 56471 20893
rect 49988 20828 51856 20856
rect 52822 20816 52828 20868
rect 52880 20856 52886 20868
rect 53024 20856 53052 20887
rect 52880 20828 53052 20856
rect 52880 20816 52886 20828
rect 54570 20816 54576 20868
rect 54628 20816 54634 20868
rect 50246 20788 50252 20800
rect 48976 20760 50252 20788
rect 50246 20748 50252 20760
rect 50304 20748 50310 20800
rect 50617 20791 50675 20797
rect 50617 20757 50629 20791
rect 50663 20788 50675 20791
rect 50798 20788 50804 20800
rect 50663 20760 50804 20788
rect 50663 20757 50675 20760
rect 50617 20751 50675 20757
rect 50798 20748 50804 20760
rect 50856 20748 50862 20800
rect 52733 20791 52791 20797
rect 52733 20757 52745 20791
rect 52779 20788 52791 20791
rect 53006 20788 53012 20800
rect 52779 20760 53012 20788
rect 52779 20757 52791 20760
rect 52733 20751 52791 20757
rect 53006 20748 53012 20760
rect 53064 20748 53070 20800
rect 53098 20748 53104 20800
rect 53156 20788 53162 20800
rect 54772 20788 54800 20887
rect 55490 20816 55496 20868
rect 55548 20856 55554 20868
rect 56428 20856 56456 20887
rect 55548 20828 56456 20856
rect 55548 20816 55554 20828
rect 53156 20760 54800 20788
rect 54941 20791 54999 20797
rect 53156 20748 53162 20760
rect 54941 20757 54953 20791
rect 54987 20788 54999 20791
rect 55122 20788 55128 20800
rect 54987 20760 55128 20788
rect 54987 20757 54999 20760
rect 54941 20751 54999 20757
rect 55122 20748 55128 20760
rect 55180 20748 55186 20800
rect 55950 20748 55956 20800
rect 56008 20788 56014 20800
rect 56689 20791 56747 20797
rect 56689 20788 56701 20791
rect 56008 20760 56701 20788
rect 56008 20748 56014 20760
rect 56689 20757 56701 20760
rect 56735 20757 56747 20791
rect 56689 20751 56747 20757
rect 1104 20698 78844 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 66314 20698
rect 66366 20646 66378 20698
rect 66430 20646 66442 20698
rect 66494 20646 66506 20698
rect 66558 20646 66570 20698
rect 66622 20646 78844 20698
rect 1104 20624 78844 20646
rect 7098 20544 7104 20596
rect 7156 20584 7162 20596
rect 7561 20587 7619 20593
rect 7561 20584 7573 20587
rect 7156 20556 7573 20584
rect 7156 20544 7162 20556
rect 7561 20553 7573 20556
rect 7607 20553 7619 20587
rect 7561 20547 7619 20553
rect 7926 20544 7932 20596
rect 7984 20584 7990 20596
rect 7984 20556 9812 20584
rect 7984 20544 7990 20556
rect 7466 20476 7472 20528
rect 7524 20516 7530 20528
rect 8113 20519 8171 20525
rect 8113 20516 8125 20519
rect 7524 20488 8125 20516
rect 7524 20476 7530 20488
rect 8113 20485 8125 20488
rect 8159 20485 8171 20519
rect 9674 20516 9680 20528
rect 9338 20488 9680 20516
rect 8113 20479 8171 20485
rect 9674 20476 9680 20488
rect 9732 20476 9738 20528
rect 9784 20516 9812 20556
rect 34698 20544 34704 20596
rect 34756 20544 34762 20596
rect 37274 20544 37280 20596
rect 37332 20544 37338 20596
rect 37550 20544 37556 20596
rect 37608 20584 37614 20596
rect 38565 20587 38623 20593
rect 37608 20556 38424 20584
rect 37608 20544 37614 20556
rect 9784 20488 10088 20516
rect 7374 20408 7380 20460
rect 7432 20448 7438 20460
rect 7561 20451 7619 20457
rect 7561 20448 7573 20451
rect 7432 20420 7573 20448
rect 7432 20408 7438 20420
rect 7561 20417 7573 20420
rect 7607 20417 7619 20451
rect 7561 20411 7619 20417
rect 7576 20380 7604 20411
rect 7650 20408 7656 20460
rect 7708 20448 7714 20460
rect 7745 20451 7803 20457
rect 7745 20448 7757 20451
rect 7708 20420 7757 20448
rect 7708 20408 7714 20420
rect 7745 20417 7757 20420
rect 7791 20417 7803 20451
rect 7745 20411 7803 20417
rect 7834 20408 7840 20460
rect 7892 20408 7898 20460
rect 9784 20457 9812 20488
rect 9769 20451 9827 20457
rect 9769 20417 9781 20451
rect 9815 20417 9827 20451
rect 9769 20411 9827 20417
rect 9953 20451 10011 20457
rect 9953 20417 9965 20451
rect 9999 20417 10011 20451
rect 9953 20411 10011 20417
rect 8570 20380 8576 20392
rect 7576 20352 8576 20380
rect 8570 20340 8576 20352
rect 8628 20380 8634 20392
rect 9490 20380 9496 20392
rect 8628 20352 9496 20380
rect 8628 20340 8634 20352
rect 9490 20340 9496 20352
rect 9548 20380 9554 20392
rect 9585 20383 9643 20389
rect 9585 20380 9597 20383
rect 9548 20352 9597 20380
rect 9548 20340 9554 20352
rect 9585 20349 9597 20352
rect 9631 20349 9643 20383
rect 9585 20343 9643 20349
rect 9968 20312 9996 20411
rect 10060 20380 10088 20488
rect 10134 20476 10140 20528
rect 10192 20516 10198 20528
rect 10192 20488 10456 20516
rect 10192 20476 10198 20488
rect 10428 20457 10456 20488
rect 11514 20476 11520 20528
rect 11572 20516 11578 20528
rect 12066 20516 12072 20528
rect 11572 20488 12072 20516
rect 11572 20476 11578 20488
rect 12066 20476 12072 20488
rect 12124 20516 12130 20528
rect 12529 20519 12587 20525
rect 12529 20516 12541 20519
rect 12124 20488 12541 20516
rect 12124 20476 12130 20488
rect 12529 20485 12541 20488
rect 12575 20485 12587 20519
rect 12529 20479 12587 20485
rect 13538 20476 13544 20528
rect 13596 20476 13602 20528
rect 19334 20476 19340 20528
rect 19392 20516 19398 20528
rect 19392 20488 22094 20516
rect 19392 20476 19398 20488
rect 10413 20451 10471 20457
rect 10413 20417 10425 20451
rect 10459 20417 10471 20451
rect 10413 20411 10471 20417
rect 10134 20380 10140 20392
rect 10060 20352 10140 20380
rect 10134 20340 10140 20352
rect 10192 20340 10198 20392
rect 10229 20383 10287 20389
rect 10229 20349 10241 20383
rect 10275 20380 10287 20383
rect 10686 20380 10692 20392
rect 10275 20352 10692 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 10244 20312 10272 20343
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 10962 20340 10968 20392
rect 11020 20380 11026 20392
rect 12253 20383 12311 20389
rect 12253 20380 12265 20383
rect 11020 20352 12265 20380
rect 11020 20340 11026 20352
rect 12253 20349 12265 20352
rect 12299 20349 12311 20383
rect 12253 20343 12311 20349
rect 14001 20383 14059 20389
rect 14001 20349 14013 20383
rect 14047 20380 14059 20383
rect 14277 20383 14335 20389
rect 14277 20380 14289 20383
rect 14047 20352 14289 20380
rect 14047 20349 14059 20352
rect 14001 20343 14059 20349
rect 14277 20349 14289 20352
rect 14323 20349 14335 20383
rect 14277 20343 14335 20349
rect 9968 20284 10272 20312
rect 9858 20204 9864 20256
rect 9916 20204 9922 20256
rect 10410 20204 10416 20256
rect 10468 20244 10474 20256
rect 10597 20247 10655 20253
rect 10597 20244 10609 20247
rect 10468 20216 10609 20244
rect 10468 20204 10474 20216
rect 10597 20213 10609 20216
rect 10643 20213 10655 20247
rect 10597 20207 10655 20213
rect 14550 20204 14556 20256
rect 14608 20244 14614 20256
rect 14921 20247 14979 20253
rect 14921 20244 14933 20247
rect 14608 20216 14933 20244
rect 14608 20204 14614 20216
rect 14921 20213 14933 20216
rect 14967 20213 14979 20247
rect 22066 20244 22094 20488
rect 33410 20476 33416 20528
rect 33468 20476 33474 20528
rect 37292 20516 37320 20544
rect 34900 20488 36676 20516
rect 23569 20451 23627 20457
rect 23569 20417 23581 20451
rect 23615 20448 23627 20451
rect 23615 20420 23796 20448
rect 23615 20417 23627 20420
rect 23569 20411 23627 20417
rect 23768 20321 23796 20420
rect 27890 20408 27896 20460
rect 27948 20408 27954 20460
rect 32122 20408 32128 20460
rect 32180 20408 32186 20460
rect 33686 20408 33692 20460
rect 33744 20448 33750 20460
rect 34900 20457 34928 20488
rect 36648 20460 36676 20488
rect 36740 20488 37320 20516
rect 34885 20451 34943 20457
rect 34885 20448 34897 20451
rect 33744 20420 34897 20448
rect 33744 20408 33750 20420
rect 34885 20417 34897 20420
rect 34931 20417 34943 20451
rect 34885 20411 34943 20417
rect 34974 20408 34980 20460
rect 35032 20408 35038 20460
rect 35253 20451 35311 20457
rect 35253 20417 35265 20451
rect 35299 20448 35311 20451
rect 35342 20448 35348 20460
rect 35299 20420 35348 20448
rect 35299 20417 35311 20420
rect 35253 20411 35311 20417
rect 35342 20408 35348 20420
rect 35400 20408 35406 20460
rect 36630 20408 36636 20460
rect 36688 20408 36694 20460
rect 36740 20457 36768 20488
rect 37642 20476 37648 20528
rect 37700 20516 37706 20528
rect 38194 20516 38200 20528
rect 37700 20488 38200 20516
rect 37700 20476 37706 20488
rect 38194 20476 38200 20488
rect 38252 20476 38258 20528
rect 38396 20457 38424 20556
rect 38565 20553 38577 20587
rect 38611 20584 38623 20587
rect 39390 20584 39396 20596
rect 38611 20556 39396 20584
rect 38611 20553 38623 20556
rect 38565 20547 38623 20553
rect 39390 20544 39396 20556
rect 39448 20544 39454 20596
rect 39669 20587 39727 20593
rect 39669 20553 39681 20587
rect 39715 20584 39727 20587
rect 40126 20584 40132 20596
rect 39715 20556 40132 20584
rect 39715 20553 39727 20556
rect 39669 20547 39727 20553
rect 40126 20544 40132 20556
rect 40184 20544 40190 20596
rect 41138 20544 41144 20596
rect 41196 20584 41202 20596
rect 41509 20587 41567 20593
rect 41509 20584 41521 20587
rect 41196 20556 41521 20584
rect 41196 20544 41202 20556
rect 41509 20553 41521 20556
rect 41555 20553 41567 20587
rect 41509 20547 41567 20553
rect 43898 20544 43904 20596
rect 43956 20584 43962 20596
rect 47026 20584 47032 20596
rect 43956 20556 47032 20584
rect 43956 20544 43962 20556
rect 43441 20519 43499 20525
rect 43441 20485 43453 20519
rect 43487 20516 43499 20519
rect 44082 20516 44088 20528
rect 43487 20488 44088 20516
rect 43487 20485 43499 20488
rect 43441 20479 43499 20485
rect 44082 20476 44088 20488
rect 44140 20476 44146 20528
rect 44358 20476 44364 20528
rect 44416 20516 44422 20528
rect 46014 20516 46020 20528
rect 44416 20488 46020 20516
rect 44416 20476 44422 20488
rect 46014 20476 46020 20488
rect 46072 20476 46078 20528
rect 36725 20451 36783 20457
rect 36725 20417 36737 20451
rect 36771 20417 36783 20451
rect 36725 20411 36783 20417
rect 37001 20451 37059 20457
rect 37001 20417 37013 20451
rect 37047 20448 37059 20451
rect 37277 20451 37335 20457
rect 37277 20448 37289 20451
rect 37047 20420 37289 20448
rect 37047 20417 37059 20420
rect 37001 20411 37059 20417
rect 37277 20417 37289 20420
rect 37323 20417 37335 20451
rect 37277 20411 37335 20417
rect 38013 20451 38071 20457
rect 38013 20417 38025 20451
rect 38059 20417 38071 20451
rect 38013 20411 38071 20417
rect 38289 20451 38347 20457
rect 38289 20417 38301 20451
rect 38335 20417 38347 20451
rect 38289 20411 38347 20417
rect 38381 20451 38439 20457
rect 38381 20417 38393 20451
rect 38427 20448 38439 20451
rect 39758 20448 39764 20460
rect 38427 20420 39764 20448
rect 38427 20417 38439 20420
rect 38381 20411 38439 20417
rect 26602 20340 26608 20392
rect 26660 20380 26666 20392
rect 28629 20383 28687 20389
rect 28629 20380 28641 20383
rect 26660 20352 28641 20380
rect 26660 20340 26666 20352
rect 28629 20349 28641 20352
rect 28675 20380 28687 20383
rect 29546 20380 29552 20392
rect 28675 20352 29552 20380
rect 28675 20349 28687 20352
rect 28629 20343 28687 20349
rect 29546 20340 29552 20352
rect 29604 20340 29610 20392
rect 32398 20340 32404 20392
rect 32456 20340 32462 20392
rect 33873 20383 33931 20389
rect 33873 20349 33885 20383
rect 33919 20380 33931 20383
rect 34514 20380 34520 20392
rect 33919 20352 34520 20380
rect 33919 20349 33931 20352
rect 33873 20343 33931 20349
rect 34514 20340 34520 20352
rect 34572 20380 34578 20392
rect 34609 20383 34667 20389
rect 34609 20380 34621 20383
rect 34572 20352 34621 20380
rect 34572 20340 34578 20352
rect 34609 20349 34621 20352
rect 34655 20349 34667 20383
rect 34609 20343 34667 20349
rect 36449 20383 36507 20389
rect 36449 20349 36461 20383
rect 36495 20380 36507 20383
rect 37458 20380 37464 20392
rect 36495 20352 37464 20380
rect 36495 20349 36507 20352
rect 36449 20343 36507 20349
rect 37458 20340 37464 20352
rect 37516 20340 37522 20392
rect 37829 20383 37887 20389
rect 37829 20349 37841 20383
rect 37875 20380 37887 20383
rect 38028 20380 38056 20411
rect 38304 20380 38332 20411
rect 39758 20408 39764 20420
rect 39816 20408 39822 20460
rect 39850 20408 39856 20460
rect 39908 20408 39914 20460
rect 39945 20451 40003 20457
rect 39945 20417 39957 20451
rect 39991 20448 40003 20451
rect 40034 20448 40040 20460
rect 39991 20420 40040 20448
rect 39991 20417 40003 20420
rect 39945 20411 40003 20417
rect 40034 20408 40040 20420
rect 40092 20408 40098 20460
rect 40221 20451 40279 20457
rect 40221 20417 40233 20451
rect 40267 20448 40279 20451
rect 40681 20451 40739 20457
rect 40681 20448 40693 20451
rect 40267 20420 40693 20448
rect 40267 20417 40279 20420
rect 40221 20411 40279 20417
rect 40681 20417 40693 20420
rect 40727 20417 40739 20451
rect 40681 20411 40739 20417
rect 41598 20408 41604 20460
rect 41656 20448 41662 20460
rect 41656 20420 41920 20448
rect 41656 20408 41662 20420
rect 41046 20380 41052 20392
rect 37875 20352 38056 20380
rect 38258 20352 41052 20380
rect 37875 20349 37887 20352
rect 37829 20343 37887 20349
rect 23753 20315 23811 20321
rect 23753 20281 23765 20315
rect 23799 20312 23811 20315
rect 31754 20312 31760 20324
rect 23799 20284 31760 20312
rect 23799 20281 23811 20284
rect 23753 20275 23811 20281
rect 31754 20272 31760 20284
rect 31812 20272 31818 20324
rect 36170 20272 36176 20324
rect 36228 20312 36234 20324
rect 37844 20312 37872 20343
rect 36228 20284 37872 20312
rect 36228 20272 36234 20284
rect 22281 20247 22339 20253
rect 22281 20244 22293 20247
rect 22066 20216 22293 20244
rect 14921 20207 14979 20213
rect 22281 20213 22293 20216
rect 22327 20244 22339 20247
rect 25406 20244 25412 20256
rect 22327 20216 25412 20244
rect 22327 20213 22339 20216
rect 22281 20207 22339 20213
rect 25406 20204 25412 20216
rect 25464 20244 25470 20256
rect 27709 20247 27767 20253
rect 27709 20244 27721 20247
rect 25464 20216 27721 20244
rect 25464 20204 25470 20216
rect 27709 20213 27721 20216
rect 27755 20244 27767 20247
rect 27890 20244 27896 20256
rect 27755 20216 27896 20244
rect 27755 20213 27767 20216
rect 27709 20207 27767 20213
rect 27890 20204 27896 20216
rect 27948 20204 27954 20256
rect 33962 20204 33968 20256
rect 34020 20204 34026 20256
rect 34422 20204 34428 20256
rect 34480 20244 34486 20256
rect 35161 20247 35219 20253
rect 35161 20244 35173 20247
rect 34480 20216 35173 20244
rect 34480 20204 34486 20216
rect 35161 20213 35173 20216
rect 35207 20213 35219 20247
rect 35161 20207 35219 20213
rect 36906 20204 36912 20256
rect 36964 20204 36970 20256
rect 36998 20204 37004 20256
rect 37056 20244 37062 20256
rect 38258 20244 38286 20352
rect 41046 20340 41052 20352
rect 41104 20380 41110 20392
rect 41233 20383 41291 20389
rect 41233 20380 41245 20383
rect 41104 20352 41245 20380
rect 41104 20340 41110 20352
rect 41233 20349 41245 20352
rect 41279 20380 41291 20383
rect 41506 20380 41512 20392
rect 41279 20352 41512 20380
rect 41279 20349 41291 20352
rect 41233 20343 41291 20349
rect 41506 20340 41512 20352
rect 41564 20340 41570 20392
rect 37056 20216 38286 20244
rect 37056 20204 37062 20216
rect 39482 20204 39488 20256
rect 39540 20244 39546 20256
rect 39850 20244 39856 20256
rect 39540 20216 39856 20244
rect 39540 20204 39546 20216
rect 39850 20204 39856 20216
rect 39908 20204 39914 20256
rect 39942 20204 39948 20256
rect 40000 20244 40006 20256
rect 41892 20253 41920 20420
rect 46658 20408 46664 20460
rect 46716 20408 46722 20460
rect 46768 20457 46796 20556
rect 47026 20544 47032 20556
rect 47084 20544 47090 20596
rect 52730 20584 52736 20596
rect 48148 20556 52736 20584
rect 47210 20476 47216 20528
rect 47268 20476 47274 20528
rect 46753 20451 46811 20457
rect 46753 20417 46765 20451
rect 46799 20417 46811 20451
rect 46753 20411 46811 20417
rect 47302 20408 47308 20460
rect 47360 20448 47366 20460
rect 48148 20457 48176 20556
rect 48682 20476 48688 20528
rect 48740 20516 48746 20528
rect 48740 20488 48898 20516
rect 48740 20476 48746 20488
rect 50540 20457 50568 20556
rect 52730 20544 52736 20556
rect 52788 20544 52794 20596
rect 55214 20584 55220 20596
rect 52932 20556 55220 20584
rect 50798 20476 50804 20528
rect 50856 20476 50862 20528
rect 52932 20516 52960 20556
rect 52026 20488 52960 20516
rect 53006 20476 53012 20528
rect 53064 20476 53070 20528
rect 53392 20516 53420 20556
rect 55214 20544 55220 20556
rect 55272 20544 55278 20596
rect 55950 20544 55956 20596
rect 56008 20584 56014 20596
rect 56008 20556 56548 20584
rect 56008 20544 56014 20556
rect 56520 20525 56548 20556
rect 56505 20519 56563 20525
rect 53392 20488 53498 20516
rect 56505 20485 56517 20519
rect 56551 20485 56563 20519
rect 56505 20479 56563 20485
rect 48133 20451 48191 20457
rect 48133 20448 48145 20451
rect 47360 20420 48145 20448
rect 47360 20408 47366 20420
rect 48133 20417 48145 20420
rect 48179 20417 48191 20451
rect 48133 20411 48191 20417
rect 50525 20451 50583 20457
rect 50525 20417 50537 20451
rect 50571 20417 50583 20451
rect 50525 20411 50583 20417
rect 52730 20408 52736 20460
rect 52788 20408 52794 20460
rect 54846 20408 54852 20460
rect 54904 20408 54910 20460
rect 55122 20408 55128 20460
rect 55180 20408 55186 20460
rect 55217 20451 55275 20457
rect 55217 20417 55229 20451
rect 55263 20448 55275 20451
rect 55490 20448 55496 20460
rect 55263 20420 55496 20448
rect 55263 20417 55275 20420
rect 55217 20411 55275 20417
rect 55490 20408 55496 20420
rect 55548 20408 55554 20460
rect 55769 20451 55827 20457
rect 55769 20448 55781 20451
rect 55600 20420 55781 20448
rect 45186 20340 45192 20392
rect 45244 20380 45250 20392
rect 46477 20383 46535 20389
rect 46477 20380 46489 20383
rect 45244 20352 46489 20380
rect 45244 20340 45250 20352
rect 46477 20349 46489 20352
rect 46523 20380 46535 20383
rect 47394 20380 47400 20392
rect 46523 20352 47400 20380
rect 46523 20349 46535 20352
rect 46477 20343 46535 20349
rect 47394 20340 47400 20352
rect 47452 20340 47458 20392
rect 48406 20340 48412 20392
rect 48464 20340 48470 20392
rect 52270 20340 52276 20392
rect 52328 20340 52334 20392
rect 54864 20380 54892 20408
rect 52840 20352 54892 20380
rect 42518 20272 42524 20324
rect 42576 20312 42582 20324
rect 43809 20315 43867 20321
rect 43809 20312 43821 20315
rect 42576 20284 43821 20312
rect 42576 20272 42582 20284
rect 43809 20281 43821 20284
rect 43855 20312 43867 20315
rect 44174 20312 44180 20324
rect 43855 20284 44180 20312
rect 43855 20281 43867 20284
rect 43809 20275 43867 20281
rect 44174 20272 44180 20284
rect 44232 20272 44238 20324
rect 52178 20272 52184 20324
rect 52236 20312 52242 20324
rect 52840 20312 52868 20352
rect 52236 20284 52868 20312
rect 52236 20272 52242 20284
rect 54202 20272 54208 20324
rect 54260 20312 54266 20324
rect 54481 20315 54539 20321
rect 54481 20312 54493 20315
rect 54260 20284 54493 20312
rect 54260 20272 54266 20284
rect 54481 20281 54493 20284
rect 54527 20281 54539 20315
rect 54481 20275 54539 20281
rect 55122 20272 55128 20324
rect 55180 20312 55186 20324
rect 55600 20321 55628 20420
rect 55769 20417 55781 20420
rect 55815 20417 55827 20451
rect 56781 20451 56839 20457
rect 56781 20448 56793 20451
rect 55769 20411 55827 20417
rect 56244 20420 56793 20448
rect 55585 20315 55643 20321
rect 55585 20312 55597 20315
rect 55180 20284 55597 20312
rect 55180 20272 55186 20284
rect 55585 20281 55597 20284
rect 55631 20281 55643 20315
rect 55585 20275 55643 20281
rect 40129 20247 40187 20253
rect 40129 20244 40141 20247
rect 40000 20216 40141 20244
rect 40000 20204 40006 20216
rect 40129 20213 40141 20216
rect 40175 20213 40187 20247
rect 40129 20207 40187 20213
rect 41877 20247 41935 20253
rect 41877 20213 41889 20247
rect 41923 20244 41935 20247
rect 44358 20244 44364 20256
rect 41923 20216 44364 20244
rect 41923 20213 41935 20216
rect 41877 20207 41935 20213
rect 44358 20204 44364 20216
rect 44416 20204 44422 20256
rect 47854 20204 47860 20256
rect 47912 20244 47918 20256
rect 48958 20244 48964 20256
rect 47912 20216 48964 20244
rect 47912 20204 47918 20216
rect 48958 20204 48964 20216
rect 49016 20204 49022 20256
rect 49510 20204 49516 20256
rect 49568 20244 49574 20256
rect 49881 20247 49939 20253
rect 49881 20244 49893 20247
rect 49568 20216 49893 20244
rect 49568 20204 49574 20216
rect 49881 20213 49893 20216
rect 49927 20213 49939 20247
rect 49881 20207 49939 20213
rect 53650 20204 53656 20256
rect 53708 20244 53714 20256
rect 54938 20244 54944 20256
rect 53708 20216 54944 20244
rect 53708 20204 53714 20216
rect 54938 20204 54944 20216
rect 54996 20204 55002 20256
rect 55398 20204 55404 20256
rect 55456 20204 55462 20256
rect 56042 20204 56048 20256
rect 56100 20244 56106 20256
rect 56244 20253 56272 20420
rect 56781 20417 56793 20420
rect 56827 20417 56839 20451
rect 56781 20411 56839 20417
rect 56229 20247 56287 20253
rect 56229 20244 56241 20247
rect 56100 20216 56241 20244
rect 56100 20204 56106 20216
rect 56229 20213 56241 20216
rect 56275 20213 56287 20247
rect 56229 20207 56287 20213
rect 56318 20204 56324 20256
rect 56376 20244 56382 20256
rect 56873 20247 56931 20253
rect 56873 20244 56885 20247
rect 56376 20216 56885 20244
rect 56376 20204 56382 20216
rect 56873 20213 56885 20216
rect 56919 20213 56931 20247
rect 56873 20207 56931 20213
rect 1104 20154 78844 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 78844 20154
rect 1104 20080 78844 20102
rect 7561 20043 7619 20049
rect 7561 20009 7573 20043
rect 7607 20040 7619 20043
rect 7650 20040 7656 20052
rect 7607 20012 7656 20040
rect 7607 20009 7619 20012
rect 7561 20003 7619 20009
rect 7374 19972 7380 19984
rect 6932 19944 7380 19972
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 6932 19836 6960 19944
rect 7374 19932 7380 19944
rect 7432 19932 7438 19984
rect 7006 19864 7012 19916
rect 7064 19904 7070 19916
rect 7064 19876 7236 19904
rect 7064 19864 7070 19876
rect 7208 19845 7236 19876
rect 7101 19839 7159 19845
rect 7101 19836 7113 19839
rect 6932 19808 7113 19836
rect 1673 19799 1731 19805
rect 7101 19805 7113 19808
rect 7147 19805 7159 19839
rect 7101 19799 7159 19805
rect 7193 19839 7251 19845
rect 7193 19805 7205 19839
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19836 7343 19839
rect 7576 19836 7604 20003
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 7745 20043 7803 20049
rect 7745 20009 7757 20043
rect 7791 20040 7803 20043
rect 7926 20040 7932 20052
rect 7791 20012 7932 20040
rect 7791 20009 7803 20012
rect 7745 20003 7803 20009
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 9858 20000 9864 20052
rect 9916 20000 9922 20052
rect 10042 20000 10048 20052
rect 10100 20000 10106 20052
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 10192 20012 11897 20040
rect 10192 20000 10198 20012
rect 11885 20009 11897 20012
rect 11931 20009 11943 20043
rect 11885 20003 11943 20009
rect 7834 19864 7840 19916
rect 7892 19904 7898 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 7892 19876 10149 19904
rect 7892 19864 7898 19876
rect 10137 19873 10149 19876
rect 10183 19904 10195 19907
rect 10962 19904 10968 19916
rect 10183 19876 10968 19904
rect 10183 19873 10195 19876
rect 10137 19867 10195 19873
rect 10962 19864 10968 19876
rect 11020 19864 11026 19916
rect 11900 19904 11928 20003
rect 27246 20000 27252 20052
rect 27304 20040 27310 20052
rect 28399 20043 28457 20049
rect 28399 20040 28411 20043
rect 27304 20012 28411 20040
rect 27304 20000 27310 20012
rect 28399 20009 28411 20012
rect 28445 20040 28457 20043
rect 30098 20040 30104 20052
rect 28445 20012 30104 20040
rect 28445 20009 28457 20012
rect 28399 20003 28457 20009
rect 30098 20000 30104 20012
rect 30156 20000 30162 20052
rect 31754 20000 31760 20052
rect 31812 20000 31818 20052
rect 32398 20000 32404 20052
rect 32456 20040 32462 20052
rect 33321 20043 33379 20049
rect 33321 20040 33333 20043
rect 32456 20012 33333 20040
rect 32456 20000 32462 20012
rect 33321 20009 33333 20012
rect 33367 20009 33379 20043
rect 33321 20003 33379 20009
rect 34054 20000 34060 20052
rect 34112 20000 34118 20052
rect 36262 20000 36268 20052
rect 36320 20040 36326 20052
rect 36633 20043 36691 20049
rect 36633 20040 36645 20043
rect 36320 20012 36645 20040
rect 36320 20000 36326 20012
rect 36633 20009 36645 20012
rect 36679 20040 36691 20043
rect 36814 20040 36820 20052
rect 36679 20012 36820 20040
rect 36679 20009 36691 20012
rect 36633 20003 36691 20009
rect 36814 20000 36820 20012
rect 36872 20000 36878 20052
rect 36906 20000 36912 20052
rect 36964 20040 36970 20052
rect 39206 20040 39212 20052
rect 36964 20012 39212 20040
rect 36964 20000 36970 20012
rect 39206 20000 39212 20012
rect 39264 20040 39270 20052
rect 39942 20040 39948 20052
rect 39264 20012 39948 20040
rect 39264 20000 39270 20012
rect 39942 20000 39948 20012
rect 40000 20000 40006 20052
rect 46477 20043 46535 20049
rect 46477 20009 46489 20043
rect 46523 20040 46535 20043
rect 47394 20040 47400 20052
rect 46523 20012 47400 20040
rect 46523 20009 46535 20012
rect 46477 20003 46535 20009
rect 47394 20000 47400 20012
rect 47452 20000 47458 20052
rect 47489 20043 47547 20049
rect 47489 20009 47501 20043
rect 47535 20009 47547 20043
rect 47489 20003 47547 20009
rect 34072 19972 34100 20000
rect 33244 19944 34100 19972
rect 12161 19907 12219 19913
rect 12161 19904 12173 19907
rect 11900 19876 12173 19904
rect 12161 19873 12173 19876
rect 12207 19873 12219 19907
rect 12161 19867 12219 19873
rect 12805 19907 12863 19913
rect 12805 19873 12817 19907
rect 12851 19904 12863 19907
rect 12851 19876 13124 19904
rect 12851 19873 12863 19876
rect 12805 19867 12863 19873
rect 7331 19808 7604 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 1688 19768 1716 19799
rect 8202 19796 8208 19848
rect 8260 19836 8266 19848
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 8260 19808 9413 19836
rect 8260 19796 8266 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 9490 19796 9496 19848
rect 9548 19796 9554 19848
rect 9861 19839 9919 19845
rect 9861 19805 9873 19839
rect 9907 19805 9919 19839
rect 9861 19799 9919 19805
rect 7834 19768 7840 19780
rect 1688 19740 7840 19768
rect 7834 19728 7840 19740
rect 7892 19768 7898 19780
rect 7929 19771 7987 19777
rect 7929 19768 7941 19771
rect 7892 19740 7941 19768
rect 7892 19728 7898 19740
rect 7929 19737 7941 19740
rect 7975 19768 7987 19771
rect 9876 19768 9904 19799
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 13096 19845 13124 19876
rect 14274 19864 14280 19916
rect 14332 19864 14338 19916
rect 14550 19864 14556 19916
rect 14608 19864 14614 19916
rect 12897 19839 12955 19845
rect 12897 19836 12909 19839
rect 12676 19808 12909 19836
rect 12676 19796 12682 19808
rect 12897 19805 12909 19808
rect 12943 19805 12955 19839
rect 12897 19799 12955 19805
rect 13081 19839 13139 19845
rect 13081 19805 13093 19839
rect 13127 19805 13139 19839
rect 13081 19799 13139 19805
rect 18506 19796 18512 19848
rect 18564 19796 18570 19848
rect 24578 19796 24584 19848
rect 24636 19836 24642 19848
rect 26602 19836 26608 19848
rect 24636 19808 26608 19836
rect 24636 19796 24642 19808
rect 26602 19796 26608 19808
rect 26660 19796 26666 19848
rect 26878 19796 26884 19848
rect 26936 19836 26942 19848
rect 33244 19845 33272 19944
rect 44542 19932 44548 19984
rect 44600 19972 44606 19984
rect 45465 19975 45523 19981
rect 45465 19972 45477 19975
rect 44600 19944 45477 19972
rect 44600 19932 44606 19944
rect 45465 19941 45477 19944
rect 45511 19941 45523 19975
rect 45465 19935 45523 19941
rect 46014 19932 46020 19984
rect 46072 19972 46078 19984
rect 46842 19972 46848 19984
rect 46072 19944 46848 19972
rect 46072 19932 46078 19944
rect 46842 19932 46848 19944
rect 46900 19972 46906 19984
rect 47504 19972 47532 20003
rect 48406 20000 48412 20052
rect 48464 20040 48470 20052
rect 48593 20043 48651 20049
rect 48593 20040 48605 20043
rect 48464 20012 48605 20040
rect 48464 20000 48470 20012
rect 48593 20009 48605 20012
rect 48639 20009 48651 20043
rect 48593 20003 48651 20009
rect 49053 20043 49111 20049
rect 49053 20009 49065 20043
rect 49099 20040 49111 20043
rect 49142 20040 49148 20052
rect 49099 20012 49148 20040
rect 49099 20009 49111 20012
rect 49053 20003 49111 20009
rect 49142 20000 49148 20012
rect 49200 20000 49206 20052
rect 50798 20040 50804 20052
rect 50356 20012 50804 20040
rect 46900 19944 47532 19972
rect 46900 19932 46906 19944
rect 48498 19932 48504 19984
rect 48556 19972 48562 19984
rect 50356 19972 50384 20012
rect 50798 20000 50804 20012
rect 50856 20000 50862 20052
rect 50890 20000 50896 20052
rect 50948 20000 50954 20052
rect 51169 20043 51227 20049
rect 51169 20009 51181 20043
rect 51215 20040 51227 20043
rect 51626 20040 51632 20052
rect 51215 20012 51632 20040
rect 51215 20009 51227 20012
rect 51169 20003 51227 20009
rect 51626 20000 51632 20012
rect 51684 20000 51690 20052
rect 52822 20000 52828 20052
rect 52880 20000 52886 20052
rect 54846 20000 54852 20052
rect 54904 20040 54910 20052
rect 55309 20043 55367 20049
rect 55309 20040 55321 20043
rect 54904 20012 55321 20040
rect 54904 20000 54910 20012
rect 55309 20009 55321 20012
rect 55355 20009 55367 20043
rect 55309 20003 55367 20009
rect 48556 19944 50384 19972
rect 48556 19932 48562 19944
rect 33686 19904 33692 19916
rect 33520 19876 33692 19904
rect 33520 19845 33548 19876
rect 33686 19864 33692 19876
rect 33744 19864 33750 19916
rect 33781 19907 33839 19913
rect 33781 19873 33793 19907
rect 33827 19904 33839 19907
rect 34422 19904 34428 19916
rect 33827 19876 34428 19904
rect 33827 19873 33839 19876
rect 33781 19867 33839 19873
rect 34422 19864 34428 19876
rect 34480 19864 34486 19916
rect 35434 19904 35440 19916
rect 34992 19876 35440 19904
rect 26973 19839 27031 19845
rect 26973 19836 26985 19839
rect 26936 19808 26985 19836
rect 26936 19796 26942 19808
rect 26973 19805 26985 19808
rect 27019 19805 27031 19839
rect 26973 19799 27031 19805
rect 33229 19839 33287 19845
rect 33229 19805 33241 19839
rect 33275 19805 33287 19839
rect 33229 19799 33287 19805
rect 33505 19839 33563 19845
rect 33505 19805 33517 19839
rect 33551 19805 33563 19839
rect 33505 19799 33563 19805
rect 33597 19839 33655 19845
rect 33597 19805 33609 19839
rect 33643 19805 33655 19839
rect 33597 19799 33655 19805
rect 33873 19839 33931 19845
rect 33873 19805 33885 19839
rect 33919 19836 33931 19839
rect 33962 19836 33968 19848
rect 33919 19808 33968 19836
rect 33919 19805 33931 19808
rect 33873 19799 33931 19805
rect 7975 19740 9904 19768
rect 7975 19737 7987 19740
rect 7929 19731 7987 19737
rect 10410 19728 10416 19780
rect 10468 19728 10474 19780
rect 28537 19771 28595 19777
rect 28537 19768 28549 19771
rect 10796 19740 10902 19768
rect 14936 19740 15042 19768
rect 28014 19740 28549 19768
rect 842 19660 848 19712
rect 900 19700 906 19712
rect 1489 19703 1547 19709
rect 1489 19700 1501 19703
rect 900 19672 1501 19700
rect 900 19660 906 19672
rect 1489 19669 1501 19672
rect 1535 19669 1547 19703
rect 1489 19663 1547 19669
rect 7466 19660 7472 19712
rect 7524 19660 7530 19712
rect 7742 19709 7748 19712
rect 7729 19703 7748 19709
rect 7729 19669 7741 19703
rect 7729 19663 7748 19669
rect 7742 19660 7748 19663
rect 7800 19660 7806 19712
rect 9674 19660 9680 19712
rect 9732 19700 9738 19712
rect 10796 19700 10824 19740
rect 14936 19712 14964 19740
rect 28537 19737 28549 19740
rect 28583 19768 28595 19771
rect 30282 19768 30288 19780
rect 28583 19740 30288 19768
rect 28583 19737 28595 19740
rect 28537 19731 28595 19737
rect 30282 19728 30288 19740
rect 30340 19728 30346 19780
rect 33612 19768 33640 19799
rect 33962 19796 33968 19808
rect 34020 19796 34026 19848
rect 34606 19796 34612 19848
rect 34664 19836 34670 19848
rect 34664 19808 34836 19836
rect 34664 19796 34670 19808
rect 34808 19768 34836 19808
rect 34882 19796 34888 19848
rect 34940 19796 34946 19848
rect 34992 19845 35020 19876
rect 35434 19864 35440 19876
rect 35492 19864 35498 19916
rect 38930 19864 38936 19916
rect 38988 19904 38994 19916
rect 39574 19904 39580 19916
rect 38988 19876 39580 19904
rect 38988 19864 38994 19876
rect 39574 19864 39580 19876
rect 39632 19904 39638 19916
rect 40678 19904 40684 19916
rect 39632 19876 40684 19904
rect 39632 19864 39638 19876
rect 40678 19864 40684 19876
rect 40736 19864 40742 19916
rect 42978 19904 42984 19916
rect 42076 19876 42984 19904
rect 34977 19839 35035 19845
rect 34977 19805 34989 19839
rect 35023 19805 35035 19839
rect 34977 19799 35035 19805
rect 35253 19839 35311 19845
rect 35253 19805 35265 19839
rect 35299 19836 35311 19839
rect 35342 19836 35348 19848
rect 35299 19808 35348 19836
rect 35299 19805 35311 19808
rect 35253 19799 35311 19805
rect 35342 19796 35348 19808
rect 35400 19796 35406 19848
rect 42076 19845 42104 19876
rect 42978 19864 42984 19876
rect 43036 19864 43042 19916
rect 45649 19907 45707 19913
rect 45649 19873 45661 19907
rect 45695 19904 45707 19907
rect 45695 19876 46796 19904
rect 45695 19873 45707 19876
rect 45649 19867 45707 19873
rect 42061 19839 42119 19845
rect 42061 19805 42073 19839
rect 42107 19805 42119 19839
rect 42061 19799 42119 19805
rect 42245 19839 42303 19845
rect 42245 19805 42257 19839
rect 42291 19836 42303 19839
rect 42702 19836 42708 19848
rect 42291 19808 42708 19836
rect 42291 19805 42303 19808
rect 42245 19799 42303 19805
rect 42702 19796 42708 19808
rect 42760 19796 42766 19848
rect 46658 19796 46664 19848
rect 46716 19796 46722 19848
rect 46768 19845 46796 19876
rect 46753 19839 46811 19845
rect 46753 19805 46765 19839
rect 46799 19836 46811 19839
rect 46934 19836 46940 19848
rect 46799 19808 46940 19836
rect 46799 19805 46811 19808
rect 46753 19799 46811 19805
rect 46934 19796 46940 19808
rect 46992 19836 46998 19848
rect 47762 19836 47768 19848
rect 46992 19808 47768 19836
rect 46992 19796 46998 19808
rect 47762 19796 47768 19808
rect 47820 19796 47826 19848
rect 48516 19836 48544 19932
rect 50246 19864 50252 19916
rect 50304 19904 50310 19916
rect 51074 19904 51080 19916
rect 50304 19876 51080 19904
rect 50304 19864 50310 19876
rect 48774 19836 48780 19848
rect 48516 19808 48780 19836
rect 48774 19796 48780 19808
rect 48832 19796 48838 19848
rect 48866 19796 48872 19848
rect 48924 19796 48930 19848
rect 49050 19796 49056 19848
rect 49108 19836 49114 19848
rect 49145 19839 49203 19845
rect 49145 19836 49157 19839
rect 49108 19808 49157 19836
rect 49108 19796 49114 19808
rect 49145 19805 49157 19808
rect 49191 19836 49203 19839
rect 49237 19839 49295 19845
rect 49237 19836 49249 19839
rect 49191 19808 49249 19836
rect 49191 19805 49203 19808
rect 49145 19799 49203 19805
rect 49237 19805 49249 19808
rect 49283 19836 49295 19839
rect 49510 19836 49516 19848
rect 49283 19808 49516 19836
rect 49283 19805 49295 19808
rect 49237 19799 49295 19805
rect 49510 19796 49516 19808
rect 49568 19836 49574 19848
rect 50157 19839 50215 19845
rect 50157 19836 50169 19839
rect 49568 19808 50169 19836
rect 49568 19796 49574 19808
rect 50157 19805 50169 19808
rect 50203 19805 50215 19839
rect 50157 19799 50215 19805
rect 50341 19839 50399 19845
rect 50341 19805 50353 19839
rect 50387 19836 50399 19839
rect 50430 19836 50436 19848
rect 50387 19808 50436 19836
rect 50387 19805 50399 19808
rect 50341 19799 50399 19805
rect 35069 19771 35127 19777
rect 35069 19768 35081 19771
rect 33612 19740 34744 19768
rect 34808 19740 35081 19768
rect 9732 19672 10824 19700
rect 9732 19660 9738 19672
rect 12986 19660 12992 19712
rect 13044 19660 13050 19712
rect 14918 19660 14924 19712
rect 14976 19660 14982 19712
rect 16025 19703 16083 19709
rect 16025 19669 16037 19703
rect 16071 19700 16083 19703
rect 17862 19700 17868 19712
rect 16071 19672 17868 19700
rect 16071 19669 16083 19672
rect 16025 19663 16083 19669
rect 17862 19660 17868 19672
rect 17920 19660 17926 19712
rect 17954 19660 17960 19712
rect 18012 19660 18018 19712
rect 28810 19660 28816 19712
rect 28868 19700 28874 19712
rect 30926 19700 30932 19712
rect 28868 19672 30932 19700
rect 28868 19660 28874 19672
rect 30926 19660 30932 19672
rect 30984 19660 30990 19712
rect 34716 19709 34744 19740
rect 35069 19737 35081 19740
rect 35115 19737 35127 19771
rect 35069 19731 35127 19737
rect 35158 19728 35164 19780
rect 35216 19768 35222 19780
rect 37918 19768 37924 19780
rect 35216 19740 37924 19768
rect 35216 19728 35222 19740
rect 37918 19728 37924 19740
rect 37976 19728 37982 19780
rect 40862 19768 40868 19780
rect 38488 19740 40868 19768
rect 38488 19712 38516 19740
rect 40862 19728 40868 19740
rect 40920 19728 40926 19780
rect 42429 19771 42487 19777
rect 42429 19737 42441 19771
rect 42475 19768 42487 19771
rect 44082 19768 44088 19780
rect 42475 19740 44088 19768
rect 42475 19737 42487 19740
rect 42429 19731 42487 19737
rect 44082 19728 44088 19740
rect 44140 19768 44146 19780
rect 44542 19768 44548 19780
rect 44140 19740 44548 19768
rect 44140 19728 44146 19740
rect 44542 19728 44548 19740
rect 44600 19768 44606 19780
rect 45189 19771 45247 19777
rect 45189 19768 45201 19771
rect 44600 19740 45201 19768
rect 44600 19728 44606 19740
rect 45189 19737 45201 19740
rect 45235 19737 45247 19771
rect 45189 19731 45247 19737
rect 47210 19728 47216 19780
rect 47268 19728 47274 19780
rect 47305 19771 47363 19777
rect 47305 19737 47317 19771
rect 47351 19768 47363 19771
rect 47394 19768 47400 19780
rect 47351 19740 47400 19768
rect 47351 19737 47363 19740
rect 47305 19731 47363 19737
rect 47394 19728 47400 19740
rect 47452 19728 47458 19780
rect 48590 19768 48596 19780
rect 47688 19740 48596 19768
rect 34701 19703 34759 19709
rect 34701 19669 34713 19703
rect 34747 19669 34759 19703
rect 34701 19663 34759 19669
rect 35986 19660 35992 19712
rect 36044 19700 36050 19712
rect 36722 19700 36728 19712
rect 36044 19672 36728 19700
rect 36044 19660 36050 19672
rect 36722 19660 36728 19672
rect 36780 19700 36786 19712
rect 36817 19703 36875 19709
rect 36817 19700 36829 19703
rect 36780 19672 36829 19700
rect 36780 19660 36786 19672
rect 36817 19669 36829 19672
rect 36863 19700 36875 19703
rect 36906 19700 36912 19712
rect 36863 19672 36912 19700
rect 36863 19669 36875 19672
rect 36817 19663 36875 19669
rect 36906 19660 36912 19672
rect 36964 19660 36970 19712
rect 38194 19660 38200 19712
rect 38252 19700 38258 19712
rect 38470 19700 38476 19712
rect 38252 19672 38476 19700
rect 38252 19660 38258 19672
rect 38470 19660 38476 19672
rect 38528 19660 38534 19712
rect 38838 19660 38844 19712
rect 38896 19700 38902 19712
rect 41877 19703 41935 19709
rect 41877 19700 41889 19703
rect 38896 19672 41889 19700
rect 38896 19660 38902 19672
rect 41877 19669 41889 19672
rect 41923 19669 41935 19703
rect 41877 19663 41935 19669
rect 42153 19703 42211 19709
rect 42153 19669 42165 19703
rect 42199 19700 42211 19703
rect 44266 19700 44272 19712
rect 42199 19672 44272 19700
rect 42199 19669 42211 19672
rect 42153 19663 42211 19669
rect 44266 19660 44272 19672
rect 44324 19660 44330 19712
rect 47026 19660 47032 19712
rect 47084 19700 47090 19712
rect 47688 19709 47716 19740
rect 48590 19728 48596 19740
rect 48648 19728 48654 19780
rect 50172 19768 50200 19799
rect 50430 19796 50436 19808
rect 50488 19796 50494 19848
rect 50522 19796 50528 19848
rect 50580 19796 50586 19848
rect 50724 19845 50752 19876
rect 51074 19864 51080 19876
rect 51132 19904 51138 19916
rect 51132 19876 52684 19904
rect 51132 19864 51138 19876
rect 50709 19839 50767 19845
rect 50709 19805 50721 19839
rect 50755 19805 50767 19839
rect 50709 19799 50767 19805
rect 50798 19796 50804 19848
rect 50856 19836 50862 19848
rect 50985 19839 51043 19845
rect 50985 19836 50997 19839
rect 50856 19808 50997 19836
rect 50856 19796 50862 19808
rect 50985 19805 50997 19808
rect 51031 19836 51043 19839
rect 51353 19839 51411 19845
rect 51353 19836 51365 19839
rect 51031 19808 51365 19836
rect 51031 19805 51043 19808
rect 50985 19799 51043 19805
rect 51353 19805 51365 19808
rect 51399 19805 51411 19839
rect 51353 19799 51411 19805
rect 52178 19796 52184 19848
rect 52236 19836 52242 19848
rect 52273 19839 52331 19845
rect 52273 19836 52285 19839
rect 52236 19808 52285 19836
rect 52236 19796 52242 19808
rect 52273 19805 52285 19808
rect 52319 19805 52331 19839
rect 52273 19799 52331 19805
rect 52362 19796 52368 19848
rect 52420 19836 52426 19848
rect 52656 19845 52684 19876
rect 55398 19864 55404 19916
rect 55456 19904 55462 19916
rect 56781 19907 56839 19913
rect 56781 19904 56793 19907
rect 55456 19876 56793 19904
rect 55456 19864 55462 19876
rect 56781 19873 56793 19876
rect 56827 19873 56839 19907
rect 56781 19867 56839 19873
rect 57054 19864 57060 19916
rect 57112 19864 57118 19916
rect 52549 19839 52607 19845
rect 52549 19836 52561 19839
rect 52420 19808 52561 19836
rect 52420 19796 52426 19808
rect 52549 19805 52561 19808
rect 52595 19805 52607 19839
rect 52549 19799 52607 19805
rect 52641 19839 52699 19845
rect 52641 19805 52653 19839
rect 52687 19836 52699 19839
rect 53098 19836 53104 19848
rect 52687 19808 53104 19836
rect 52687 19805 52699 19808
rect 52641 19799 52699 19805
rect 53098 19796 53104 19808
rect 53156 19796 53162 19848
rect 50617 19771 50675 19777
rect 50617 19768 50629 19771
rect 50172 19740 50629 19768
rect 50617 19737 50629 19740
rect 50663 19737 50675 19771
rect 52457 19771 52515 19777
rect 52457 19768 52469 19771
rect 50617 19731 50675 19737
rect 52380 19740 52469 19768
rect 52380 19712 52408 19740
rect 52457 19737 52469 19740
rect 52503 19768 52515 19771
rect 54570 19768 54576 19780
rect 52503 19740 54576 19768
rect 52503 19737 52515 19740
rect 52457 19731 52515 19737
rect 54570 19728 54576 19740
rect 54628 19728 54634 19780
rect 55214 19728 55220 19780
rect 55272 19768 55278 19780
rect 55272 19740 55614 19768
rect 55272 19728 55278 19740
rect 47505 19703 47563 19709
rect 47505 19700 47517 19703
rect 47084 19672 47517 19700
rect 47084 19660 47090 19672
rect 47505 19669 47517 19672
rect 47551 19669 47563 19703
rect 47505 19663 47563 19669
rect 47673 19703 47731 19709
rect 47673 19669 47685 19703
rect 47719 19669 47731 19703
rect 47673 19663 47731 19669
rect 50522 19660 50528 19712
rect 50580 19700 50586 19712
rect 52362 19700 52368 19712
rect 50580 19672 52368 19700
rect 50580 19660 50586 19672
rect 52362 19660 52368 19672
rect 52420 19660 52426 19712
rect 1104 19610 78844 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 66314 19610
rect 66366 19558 66378 19610
rect 66430 19558 66442 19610
rect 66494 19558 66506 19610
rect 66558 19558 66570 19610
rect 66622 19558 78844 19610
rect 1104 19536 78844 19558
rect 12066 19456 12072 19508
rect 12124 19456 12130 19508
rect 14461 19499 14519 19505
rect 14461 19465 14473 19499
rect 14507 19496 14519 19499
rect 15470 19496 15476 19508
rect 14507 19468 15476 19496
rect 14507 19465 14519 19468
rect 14461 19459 14519 19465
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 37093 19499 37151 19505
rect 25240 19468 28212 19496
rect 12986 19388 12992 19440
rect 13044 19388 13050 19440
rect 13998 19388 14004 19440
rect 14056 19388 14062 19440
rect 17856 19431 17914 19437
rect 17856 19397 17868 19431
rect 17902 19428 17914 19431
rect 17954 19428 17960 19440
rect 17902 19400 17960 19428
rect 17902 19397 17914 19400
rect 17856 19391 17914 19397
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 24946 19388 24952 19440
rect 25004 19428 25010 19440
rect 25240 19428 25268 19468
rect 25004 19400 25346 19428
rect 25004 19388 25010 19400
rect 26602 19388 26608 19440
rect 26660 19428 26666 19440
rect 28184 19428 28212 19468
rect 37093 19465 37105 19499
rect 37139 19496 37151 19499
rect 37139 19468 37596 19496
rect 37139 19465 37151 19468
rect 37093 19459 37151 19465
rect 28810 19428 28816 19440
rect 26660 19400 28120 19428
rect 28184 19400 28816 19428
rect 26660 19388 26666 19400
rect 7466 19320 7472 19372
rect 7524 19360 7530 19372
rect 7561 19363 7619 19369
rect 7561 19360 7573 19363
rect 7524 19332 7573 19360
rect 7524 19320 7530 19332
rect 7561 19329 7573 19332
rect 7607 19329 7619 19363
rect 7561 19323 7619 19329
rect 7742 19320 7748 19372
rect 7800 19320 7806 19372
rect 7834 19320 7840 19372
rect 7892 19320 7898 19372
rect 10594 19320 10600 19372
rect 10652 19320 10658 19372
rect 10781 19363 10839 19369
rect 10781 19329 10793 19363
rect 10827 19360 10839 19363
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 10827 19332 12173 19360
rect 10827 19329 10839 19332
rect 10781 19323 10839 19329
rect 12161 19329 12173 19332
rect 12207 19360 12219 19363
rect 12618 19360 12624 19372
rect 12207 19332 12624 19360
rect 12207 19329 12219 19332
rect 12161 19323 12219 19329
rect 9490 19252 9496 19304
rect 9548 19292 9554 19304
rect 9861 19295 9919 19301
rect 9861 19292 9873 19295
rect 9548 19264 9873 19292
rect 9548 19252 9554 19264
rect 9861 19261 9873 19264
rect 9907 19261 9919 19295
rect 9861 19255 9919 19261
rect 10042 19252 10048 19304
rect 10100 19292 10106 19304
rect 10796 19292 10824 19323
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 12710 19320 12716 19372
rect 12768 19320 12774 19372
rect 16574 19320 16580 19372
rect 16632 19360 16638 19372
rect 17589 19363 17647 19369
rect 17589 19360 17601 19363
rect 16632 19332 17601 19360
rect 16632 19320 16638 19332
rect 17589 19329 17601 19332
rect 17635 19329 17647 19363
rect 17589 19323 17647 19329
rect 24578 19320 24584 19372
rect 24636 19320 24642 19372
rect 26878 19320 26884 19372
rect 26936 19320 26942 19372
rect 26970 19320 26976 19372
rect 27028 19360 27034 19372
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 27028 19332 27169 19360
rect 27028 19320 27034 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 27246 19320 27252 19372
rect 27304 19320 27310 19372
rect 27338 19320 27344 19372
rect 27396 19320 27402 19372
rect 27522 19320 27528 19372
rect 27580 19320 27586 19372
rect 28092 19369 28120 19400
rect 28810 19388 28816 19400
rect 28868 19388 28874 19440
rect 30926 19388 30932 19440
rect 30984 19388 30990 19440
rect 35158 19428 35164 19440
rect 32784 19400 35164 19428
rect 28077 19363 28135 19369
rect 28077 19329 28089 19363
rect 28123 19329 28135 19363
rect 28077 19323 28135 19329
rect 29638 19320 29644 19372
rect 29696 19360 29702 19372
rect 32784 19369 32812 19400
rect 35158 19388 35164 19400
rect 35216 19388 35222 19440
rect 35434 19388 35440 19440
rect 35492 19428 35498 19440
rect 35492 19400 36584 19428
rect 35492 19388 35498 19400
rect 30193 19363 30251 19369
rect 30193 19360 30205 19363
rect 29696 19332 30205 19360
rect 29696 19320 29702 19332
rect 30193 19329 30205 19332
rect 30239 19329 30251 19363
rect 32769 19363 32827 19369
rect 32769 19360 32781 19363
rect 30193 19323 30251 19329
rect 31956 19332 32781 19360
rect 19242 19292 19248 19304
rect 10100 19264 10824 19292
rect 18984 19264 19248 19292
rect 10100 19252 10106 19264
rect 18984 19233 19012 19264
rect 19242 19252 19248 19264
rect 19300 19292 19306 19304
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 19300 19264 19625 19292
rect 19300 19252 19306 19264
rect 19613 19261 19625 19264
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 24854 19252 24860 19304
rect 24912 19252 24918 19304
rect 18969 19227 19027 19233
rect 18969 19193 18981 19227
rect 19015 19193 19027 19227
rect 26896 19224 26924 19320
rect 28350 19252 28356 19304
rect 28408 19252 28414 19304
rect 29822 19252 29828 19304
rect 29880 19252 29886 19304
rect 30469 19295 30527 19301
rect 30469 19261 30481 19295
rect 30515 19292 30527 19295
rect 31110 19292 31116 19304
rect 30515 19264 31116 19292
rect 30515 19261 30527 19264
rect 30469 19255 30527 19261
rect 31110 19252 31116 19264
rect 31168 19252 31174 19304
rect 31956 19301 31984 19332
rect 32769 19329 32781 19332
rect 32815 19329 32827 19363
rect 32769 19323 32827 19329
rect 32950 19320 32956 19372
rect 33008 19360 33014 19372
rect 33045 19363 33103 19369
rect 33045 19360 33057 19363
rect 33008 19332 33057 19360
rect 33008 19320 33014 19332
rect 33045 19329 33057 19332
rect 33091 19360 33103 19363
rect 34882 19360 34888 19372
rect 33091 19332 34888 19360
rect 33091 19329 33103 19332
rect 33045 19323 33103 19329
rect 34882 19320 34888 19332
rect 34940 19320 34946 19372
rect 35342 19320 35348 19372
rect 35400 19360 35406 19372
rect 35897 19363 35955 19369
rect 35897 19360 35909 19363
rect 35400 19332 35909 19360
rect 35400 19320 35406 19332
rect 35897 19329 35909 19332
rect 35943 19329 35955 19363
rect 35897 19323 35955 19329
rect 35986 19320 35992 19372
rect 36044 19360 36050 19372
rect 36081 19363 36139 19369
rect 36081 19360 36093 19363
rect 36044 19332 36093 19360
rect 36044 19320 36050 19332
rect 36081 19329 36093 19332
rect 36127 19329 36139 19363
rect 36081 19323 36139 19329
rect 36170 19320 36176 19372
rect 36228 19320 36234 19372
rect 36262 19320 36268 19372
rect 36320 19320 36326 19372
rect 36556 19369 36584 19400
rect 36541 19363 36599 19369
rect 36541 19329 36553 19363
rect 36587 19329 36599 19363
rect 36541 19323 36599 19329
rect 36722 19320 36728 19372
rect 36780 19320 36786 19372
rect 36814 19320 36820 19372
rect 36872 19320 36878 19372
rect 36909 19363 36967 19369
rect 36909 19329 36921 19363
rect 36955 19360 36967 19363
rect 37182 19360 37188 19372
rect 36955 19332 37188 19360
rect 36955 19329 36967 19332
rect 36909 19323 36967 19329
rect 37182 19320 37188 19332
rect 37240 19320 37246 19372
rect 37568 19369 37596 19468
rect 37642 19456 37648 19508
rect 37700 19496 37706 19508
rect 38010 19496 38016 19508
rect 37700 19468 38016 19496
rect 37700 19456 37706 19468
rect 38010 19456 38016 19468
rect 38068 19496 38074 19508
rect 38286 19496 38292 19508
rect 38068 19468 38292 19496
rect 38068 19456 38074 19468
rect 38286 19456 38292 19468
rect 38344 19456 38350 19508
rect 38378 19456 38384 19508
rect 38436 19456 38442 19508
rect 38470 19456 38476 19508
rect 38528 19496 38534 19508
rect 38528 19468 38654 19496
rect 38528 19456 38534 19468
rect 37660 19428 37688 19456
rect 37660 19400 37872 19428
rect 37844 19369 37872 19400
rect 37918 19388 37924 19440
rect 37976 19388 37982 19440
rect 38396 19428 38424 19456
rect 38120 19400 38424 19428
rect 38626 19428 38654 19468
rect 40034 19456 40040 19508
rect 40092 19456 40098 19508
rect 41417 19499 41475 19505
rect 41417 19465 41429 19499
rect 41463 19496 41475 19499
rect 42610 19496 42616 19508
rect 41463 19468 42616 19496
rect 41463 19465 41475 19468
rect 41417 19459 41475 19465
rect 42610 19456 42616 19468
rect 42668 19456 42674 19508
rect 43257 19499 43315 19505
rect 43257 19465 43269 19499
rect 43303 19496 43315 19499
rect 43438 19496 43444 19508
rect 43303 19468 43444 19496
rect 43303 19465 43315 19468
rect 43257 19459 43315 19465
rect 43438 19456 43444 19468
rect 43496 19456 43502 19508
rect 43533 19499 43591 19505
rect 43533 19465 43545 19499
rect 43579 19496 43591 19499
rect 43622 19496 43628 19508
rect 43579 19468 43628 19496
rect 43579 19465 43591 19468
rect 43533 19459 43591 19465
rect 43622 19456 43628 19468
rect 43680 19456 43686 19508
rect 44266 19456 44272 19508
rect 44324 19456 44330 19508
rect 44453 19499 44511 19505
rect 44453 19465 44465 19499
rect 44499 19496 44511 19499
rect 45186 19496 45192 19508
rect 44499 19468 45192 19496
rect 44499 19465 44511 19468
rect 44453 19459 44511 19465
rect 45186 19456 45192 19468
rect 45244 19456 45250 19508
rect 47118 19456 47124 19508
rect 47176 19496 47182 19508
rect 47305 19499 47363 19505
rect 47305 19496 47317 19499
rect 47176 19468 47317 19496
rect 47176 19456 47182 19468
rect 47305 19465 47317 19468
rect 47351 19465 47363 19499
rect 47305 19459 47363 19465
rect 47581 19499 47639 19505
rect 47581 19465 47593 19499
rect 47627 19496 47639 19499
rect 48498 19496 48504 19508
rect 47627 19468 48504 19496
rect 47627 19465 47639 19468
rect 47581 19459 47639 19465
rect 48498 19456 48504 19468
rect 48556 19456 48562 19508
rect 40497 19431 40555 19437
rect 38626 19400 39712 19428
rect 37553 19363 37611 19369
rect 37553 19329 37565 19363
rect 37599 19329 37611 19363
rect 37553 19323 37611 19329
rect 37701 19363 37759 19369
rect 37701 19329 37713 19363
rect 37747 19360 37759 19363
rect 37829 19363 37887 19369
rect 37747 19329 37780 19360
rect 37701 19323 37780 19329
rect 37829 19329 37841 19363
rect 37875 19329 37887 19363
rect 37829 19323 37887 19329
rect 31941 19295 31999 19301
rect 31941 19261 31953 19295
rect 31987 19261 31999 19295
rect 31941 19255 31999 19261
rect 32674 19252 32680 19304
rect 32732 19292 32738 19304
rect 33229 19295 33287 19301
rect 33229 19292 33241 19295
rect 32732 19264 33241 19292
rect 32732 19252 32738 19264
rect 33229 19261 33241 19264
rect 33275 19292 33287 19295
rect 36740 19292 36768 19320
rect 37366 19292 37372 19304
rect 33275 19264 36676 19292
rect 36740 19264 37372 19292
rect 33275 19261 33287 19264
rect 33229 19255 33287 19261
rect 26973 19227 27031 19233
rect 26973 19224 26985 19227
rect 26896 19196 26985 19224
rect 18969 19187 19027 19193
rect 26973 19193 26985 19196
rect 27019 19193 27031 19227
rect 36538 19224 36544 19236
rect 26973 19187 27031 19193
rect 31726 19196 36544 19224
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 7377 19159 7435 19165
rect 7377 19156 7389 19159
rect 7340 19128 7389 19156
rect 7340 19116 7346 19128
rect 7377 19125 7389 19128
rect 7423 19125 7435 19159
rect 7377 19119 7435 19125
rect 10226 19116 10232 19168
rect 10284 19156 10290 19168
rect 10505 19159 10563 19165
rect 10505 19156 10517 19159
rect 10284 19128 10517 19156
rect 10284 19116 10290 19128
rect 10505 19125 10517 19128
rect 10551 19125 10563 19159
rect 10505 19119 10563 19125
rect 10778 19116 10784 19168
rect 10836 19116 10842 19168
rect 19058 19116 19064 19168
rect 19116 19116 19122 19168
rect 26234 19116 26240 19168
rect 26292 19156 26298 19168
rect 26329 19159 26387 19165
rect 26329 19156 26341 19159
rect 26292 19128 26341 19156
rect 26292 19116 26298 19128
rect 26329 19125 26341 19128
rect 26375 19156 26387 19159
rect 31726 19156 31754 19196
rect 36538 19184 36544 19196
rect 36596 19184 36602 19236
rect 36648 19224 36676 19264
rect 37366 19252 37372 19264
rect 37424 19252 37430 19304
rect 37752 19292 37780 19323
rect 38010 19320 38016 19372
rect 38068 19369 38074 19372
rect 38068 19360 38076 19369
rect 38120 19360 38148 19400
rect 38930 19360 38936 19372
rect 38068 19332 38148 19360
rect 38212 19332 38936 19360
rect 38068 19323 38076 19332
rect 38068 19320 38074 19323
rect 38212 19292 38240 19332
rect 38930 19320 38936 19332
rect 38988 19320 38994 19372
rect 39485 19363 39543 19369
rect 39485 19329 39497 19363
rect 39531 19360 39543 19363
rect 39574 19360 39580 19372
rect 39531 19332 39580 19360
rect 39531 19329 39543 19332
rect 39485 19323 39543 19329
rect 39574 19320 39580 19332
rect 39632 19320 39638 19372
rect 39684 19369 39712 19400
rect 40497 19397 40509 19431
rect 40543 19428 40555 19431
rect 41601 19431 41659 19437
rect 41601 19428 41613 19431
rect 40543 19400 41613 19428
rect 40543 19397 40555 19400
rect 40497 19391 40555 19397
rect 41601 19397 41613 19400
rect 41647 19428 41659 19431
rect 42334 19428 42340 19440
rect 41647 19400 42340 19428
rect 41647 19397 41659 19400
rect 41601 19391 41659 19397
rect 42334 19388 42340 19400
rect 42392 19428 42398 19440
rect 42886 19428 42892 19440
rect 42392 19400 42892 19428
rect 42392 19388 42398 19400
rect 42886 19388 42892 19400
rect 42944 19388 42950 19440
rect 46842 19388 46848 19440
rect 46900 19428 46906 19440
rect 47857 19431 47915 19437
rect 47857 19428 47869 19431
rect 46900 19400 47869 19428
rect 46900 19388 46906 19400
rect 47857 19397 47869 19400
rect 47903 19397 47915 19431
rect 47857 19391 47915 19397
rect 47946 19388 47952 19440
rect 48004 19388 48010 19440
rect 48682 19388 48688 19440
rect 48740 19428 48746 19440
rect 56042 19428 56048 19440
rect 48740 19400 56048 19428
rect 48740 19388 48746 19400
rect 56042 19388 56048 19400
rect 56100 19388 56106 19440
rect 39669 19363 39727 19369
rect 39669 19329 39681 19363
rect 39715 19329 39727 19363
rect 39669 19323 39727 19329
rect 39761 19363 39819 19369
rect 39761 19329 39773 19363
rect 39807 19329 39819 19363
rect 39761 19323 39819 19329
rect 37752 19264 38240 19292
rect 38286 19252 38292 19304
rect 38344 19292 38350 19304
rect 38473 19295 38531 19301
rect 38473 19292 38485 19295
rect 38344 19264 38485 19292
rect 38344 19252 38350 19264
rect 38473 19261 38485 19264
rect 38519 19261 38531 19295
rect 38473 19255 38531 19261
rect 38746 19252 38752 19304
rect 38804 19292 38810 19304
rect 39022 19292 39028 19304
rect 38804 19264 39028 19292
rect 38804 19252 38810 19264
rect 39022 19252 39028 19264
rect 39080 19252 39086 19304
rect 39390 19252 39396 19304
rect 39448 19292 39454 19304
rect 39776 19292 39804 19323
rect 39850 19320 39856 19372
rect 39908 19360 39914 19372
rect 40218 19360 40224 19372
rect 39908 19332 40224 19360
rect 39908 19320 39914 19332
rect 40218 19320 40224 19332
rect 40276 19320 40282 19372
rect 40310 19320 40316 19372
rect 40368 19320 40374 19372
rect 40405 19363 40463 19369
rect 40405 19329 40417 19363
rect 40451 19329 40463 19363
rect 40405 19323 40463 19329
rect 39448 19264 39804 19292
rect 39448 19252 39454 19264
rect 40034 19252 40040 19304
rect 40092 19292 40098 19304
rect 40420 19292 40448 19323
rect 40678 19320 40684 19372
rect 40736 19320 40742 19372
rect 40770 19320 40776 19372
rect 40828 19366 40834 19372
rect 40865 19366 40923 19369
rect 40828 19363 40923 19366
rect 40828 19338 40877 19363
rect 40828 19320 40834 19338
rect 40865 19329 40877 19338
rect 40911 19329 40923 19363
rect 40865 19323 40923 19329
rect 40954 19320 40960 19372
rect 41012 19350 41018 19372
rect 41049 19363 41107 19369
rect 41049 19350 41061 19363
rect 41012 19329 41061 19350
rect 41095 19329 41107 19363
rect 41012 19323 41107 19329
rect 41141 19363 41199 19369
rect 41141 19329 41153 19363
rect 41187 19329 41199 19363
rect 41257 19363 41315 19369
rect 41257 19360 41269 19363
rect 41141 19323 41199 19329
rect 41248 19329 41269 19360
rect 41303 19329 41315 19363
rect 41248 19323 41315 19329
rect 43073 19363 43131 19369
rect 43073 19329 43085 19363
rect 43119 19329 43131 19363
rect 43073 19323 43131 19329
rect 41012 19322 41092 19323
rect 41012 19320 41018 19322
rect 41156 19292 41184 19323
rect 40092 19264 41184 19292
rect 40092 19252 40098 19264
rect 39114 19224 39120 19236
rect 36648 19196 39120 19224
rect 39114 19184 39120 19196
rect 39172 19184 39178 19236
rect 40310 19184 40316 19236
rect 40368 19224 40374 19236
rect 41248 19224 41276 19323
rect 40368 19196 41276 19224
rect 40368 19184 40374 19196
rect 26375 19128 31754 19156
rect 26375 19125 26387 19128
rect 26329 19119 26387 19125
rect 32122 19116 32128 19168
rect 32180 19116 32186 19168
rect 32858 19116 32864 19168
rect 32916 19116 32922 19168
rect 32950 19116 32956 19168
rect 33008 19156 33014 19168
rect 33410 19156 33416 19168
rect 33008 19128 33416 19156
rect 33008 19116 33014 19128
rect 33410 19116 33416 19128
rect 33468 19156 33474 19168
rect 34606 19156 34612 19168
rect 33468 19128 34612 19156
rect 33468 19116 33474 19128
rect 34606 19116 34612 19128
rect 34664 19116 34670 19168
rect 36449 19159 36507 19165
rect 36449 19125 36461 19159
rect 36495 19156 36507 19159
rect 37182 19156 37188 19168
rect 36495 19128 37188 19156
rect 36495 19125 36507 19128
rect 36449 19119 36507 19125
rect 37182 19116 37188 19128
rect 37240 19116 37246 19168
rect 38194 19116 38200 19168
rect 38252 19116 38258 19168
rect 38378 19116 38384 19168
rect 38436 19156 38442 19168
rect 39850 19156 39856 19168
rect 38436 19128 39856 19156
rect 38436 19116 38442 19128
rect 39850 19116 39856 19128
rect 39908 19116 39914 19168
rect 40126 19116 40132 19168
rect 40184 19116 40190 19168
rect 41506 19116 41512 19168
rect 41564 19156 41570 19168
rect 42429 19159 42487 19165
rect 42429 19156 42441 19159
rect 41564 19128 42441 19156
rect 41564 19116 41570 19128
rect 42429 19125 42441 19128
rect 42475 19125 42487 19159
rect 42429 19119 42487 19125
rect 42981 19159 43039 19165
rect 42981 19125 42993 19159
rect 43027 19156 43039 19159
rect 43088 19156 43116 19323
rect 43714 19320 43720 19372
rect 43772 19320 43778 19372
rect 44174 19320 44180 19372
rect 44232 19320 44238 19372
rect 44542 19320 44548 19372
rect 44600 19320 44606 19372
rect 47762 19320 47768 19372
rect 47820 19320 47826 19372
rect 48067 19363 48125 19369
rect 48067 19360 48079 19363
rect 47872 19332 48079 19360
rect 43254 19252 43260 19304
rect 43312 19292 43318 19304
rect 43809 19295 43867 19301
rect 43809 19292 43821 19295
rect 43312 19264 43821 19292
rect 43312 19252 43318 19264
rect 43809 19261 43821 19264
rect 43855 19261 43867 19295
rect 43809 19255 43867 19261
rect 44634 19252 44640 19304
rect 44692 19252 44698 19304
rect 47118 19252 47124 19304
rect 47176 19292 47182 19304
rect 47872 19292 47900 19332
rect 48067 19329 48079 19332
rect 48113 19329 48125 19363
rect 48067 19323 48125 19329
rect 49142 19320 49148 19372
rect 49200 19360 49206 19372
rect 50985 19363 51043 19369
rect 50985 19360 50997 19363
rect 49200 19332 50997 19360
rect 49200 19320 49206 19332
rect 50985 19329 50997 19332
rect 51031 19329 51043 19363
rect 50985 19323 51043 19329
rect 47176 19264 47900 19292
rect 47176 19252 47182 19264
rect 48222 19252 48228 19304
rect 48280 19252 48286 19304
rect 48130 19184 48136 19236
rect 48188 19224 48194 19236
rect 48866 19224 48872 19236
rect 48188 19196 48872 19224
rect 48188 19184 48194 19196
rect 48866 19184 48872 19196
rect 48924 19184 48930 19236
rect 43806 19156 43812 19168
rect 43027 19128 43812 19156
rect 43027 19125 43039 19128
rect 42981 19119 43039 19125
rect 43806 19116 43812 19128
rect 43864 19116 43870 19168
rect 44818 19116 44824 19168
rect 44876 19116 44882 19168
rect 51169 19159 51227 19165
rect 51169 19125 51181 19159
rect 51215 19156 51227 19159
rect 51350 19156 51356 19168
rect 51215 19128 51356 19156
rect 51215 19125 51227 19128
rect 51169 19119 51227 19125
rect 51350 19116 51356 19128
rect 51408 19116 51414 19168
rect 1104 19066 78844 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 78844 19066
rect 1104 18992 78844 19014
rect 7834 18912 7840 18964
rect 7892 18952 7898 18964
rect 8757 18955 8815 18961
rect 8757 18952 8769 18955
rect 7892 18924 8769 18952
rect 7892 18912 7898 18924
rect 8757 18921 8769 18924
rect 8803 18952 8815 18955
rect 8803 18924 9628 18952
rect 8803 18921 8815 18924
rect 8757 18915 8815 18921
rect 7009 18819 7067 18825
rect 7009 18785 7021 18819
rect 7055 18816 7067 18819
rect 9490 18816 9496 18828
rect 7055 18788 9496 18816
rect 7055 18785 7067 18788
rect 7009 18779 7067 18785
rect 9490 18776 9496 18788
rect 9548 18776 9554 18828
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18748 9459 18751
rect 9600 18748 9628 18924
rect 10778 18912 10784 18964
rect 10836 18952 10842 18964
rect 15914 18955 15972 18961
rect 15914 18952 15926 18955
rect 10836 18924 15926 18952
rect 10836 18912 10842 18924
rect 15914 18921 15926 18924
rect 15960 18921 15972 18955
rect 15914 18915 15972 18921
rect 18049 18955 18107 18961
rect 18049 18921 18061 18955
rect 18095 18952 18107 18955
rect 18506 18952 18512 18964
rect 18095 18924 18512 18952
rect 18095 18921 18107 18924
rect 18049 18915 18107 18921
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 28350 18912 28356 18964
rect 28408 18912 28414 18964
rect 29822 18912 29828 18964
rect 29880 18912 29886 18964
rect 31110 18912 31116 18964
rect 31168 18912 31174 18964
rect 31573 18955 31631 18961
rect 31573 18921 31585 18955
rect 31619 18952 31631 18955
rect 32398 18952 32404 18964
rect 31619 18924 32404 18952
rect 31619 18921 31631 18924
rect 31573 18915 31631 18921
rect 32398 18912 32404 18924
rect 32456 18912 32462 18964
rect 35434 18952 35440 18964
rect 32968 18924 35440 18952
rect 19521 18887 19579 18893
rect 19521 18884 19533 18887
rect 18524 18856 19533 18884
rect 15657 18819 15715 18825
rect 15657 18785 15669 18819
rect 15703 18816 15715 18819
rect 16482 18816 16488 18828
rect 15703 18788 16488 18816
rect 15703 18785 15715 18788
rect 15657 18779 15715 18785
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 17862 18776 17868 18828
rect 17920 18816 17926 18828
rect 18524 18825 18552 18856
rect 19521 18853 19533 18856
rect 19567 18853 19579 18887
rect 19521 18847 19579 18853
rect 18509 18819 18567 18825
rect 18509 18816 18521 18819
rect 17920 18788 18521 18816
rect 17920 18776 17926 18788
rect 18509 18785 18521 18788
rect 18555 18785 18567 18819
rect 18509 18779 18567 18785
rect 18598 18776 18604 18828
rect 18656 18776 18662 18828
rect 19242 18776 19248 18828
rect 19300 18776 19306 18828
rect 28997 18819 29055 18825
rect 28997 18785 29009 18819
rect 29043 18816 29055 18819
rect 29840 18816 29868 18912
rect 32858 18884 32864 18896
rect 31726 18856 32864 18884
rect 31726 18816 31754 18856
rect 32858 18844 32864 18856
rect 32916 18844 32922 18896
rect 32968 18816 32996 18924
rect 35434 18912 35440 18924
rect 35492 18912 35498 18964
rect 37274 18912 37280 18964
rect 37332 18912 37338 18964
rect 37734 18912 37740 18964
rect 37792 18952 37798 18964
rect 38102 18952 38108 18964
rect 37792 18924 38108 18952
rect 37792 18912 37798 18924
rect 38102 18912 38108 18924
rect 38160 18912 38166 18964
rect 38194 18912 38200 18964
rect 38252 18912 38258 18964
rect 38565 18955 38623 18961
rect 38565 18921 38577 18955
rect 38611 18952 38623 18955
rect 38746 18952 38752 18964
rect 38611 18924 38752 18952
rect 38611 18921 38623 18924
rect 38565 18915 38623 18921
rect 38746 18912 38752 18924
rect 38804 18912 38810 18964
rect 39040 18924 39896 18952
rect 33502 18844 33508 18896
rect 33560 18884 33566 18896
rect 34514 18884 34520 18896
rect 33560 18856 34520 18884
rect 33560 18844 33566 18856
rect 34514 18844 34520 18856
rect 34572 18884 34578 18896
rect 36817 18887 36875 18893
rect 34572 18856 36309 18884
rect 34572 18844 34578 18856
rect 29043 18788 29868 18816
rect 31404 18788 31754 18816
rect 32416 18788 32996 18816
rect 33060 18788 33640 18816
rect 29043 18785 29055 18788
rect 28997 18779 29055 18785
rect 9447 18720 9628 18748
rect 9447 18717 9459 18720
rect 9401 18711 9459 18717
rect 9766 18708 9772 18760
rect 9824 18748 9830 18760
rect 10042 18748 10048 18760
rect 9824 18720 10048 18748
rect 9824 18708 9830 18720
rect 10042 18708 10048 18720
rect 10100 18708 10106 18760
rect 10226 18708 10232 18760
rect 10284 18708 10290 18760
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 19058 18748 19064 18760
rect 18463 18720 19064 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 19058 18708 19064 18720
rect 19116 18708 19122 18760
rect 23293 18751 23351 18757
rect 23293 18717 23305 18751
rect 23339 18748 23351 18751
rect 23842 18748 23848 18760
rect 23339 18720 23848 18748
rect 23339 18717 23351 18720
rect 23293 18711 23351 18717
rect 23842 18708 23848 18720
rect 23900 18708 23906 18760
rect 27338 18708 27344 18760
rect 27396 18748 27402 18760
rect 28478 18751 28536 18757
rect 28478 18748 28490 18751
rect 27396 18720 28490 18748
rect 27396 18708 27402 18720
rect 28478 18717 28490 18720
rect 28524 18717 28536 18751
rect 28478 18711 28536 18717
rect 28905 18751 28963 18757
rect 28905 18717 28917 18751
rect 28951 18748 28963 18751
rect 28951 18720 29500 18748
rect 28951 18717 28963 18720
rect 28905 18711 28963 18717
rect 7282 18640 7288 18692
rect 7340 18640 7346 18692
rect 9306 18680 9312 18692
rect 8510 18652 9312 18680
rect 9306 18640 9312 18652
rect 9364 18640 9370 18692
rect 14918 18640 14924 18692
rect 14976 18680 14982 18692
rect 17954 18680 17960 18692
rect 14976 18652 16422 18680
rect 17328 18652 17960 18680
rect 14976 18640 14982 18652
rect 9858 18572 9864 18624
rect 9916 18612 9922 18624
rect 9953 18615 10011 18621
rect 9953 18612 9965 18615
rect 9916 18584 9965 18612
rect 9916 18572 9922 18584
rect 9953 18581 9965 18584
rect 9999 18581 10011 18615
rect 9953 18575 10011 18581
rect 10137 18615 10195 18621
rect 10137 18581 10149 18615
rect 10183 18612 10195 18615
rect 10686 18612 10692 18624
rect 10183 18584 10692 18612
rect 10183 18581 10195 18584
rect 10137 18575 10195 18581
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 16316 18612 16344 18652
rect 17328 18612 17356 18652
rect 17954 18640 17960 18652
rect 18012 18680 18018 18692
rect 18598 18680 18604 18692
rect 18012 18652 18604 18680
rect 18012 18640 18018 18652
rect 18598 18640 18604 18652
rect 18656 18640 18662 18692
rect 28074 18640 28080 18692
rect 28132 18680 28138 18692
rect 28261 18683 28319 18689
rect 28261 18680 28273 18683
rect 28132 18652 28273 18680
rect 28132 18640 28138 18652
rect 28261 18649 28273 18652
rect 28307 18680 28319 18683
rect 28626 18680 28632 18692
rect 28307 18652 28632 18680
rect 28307 18649 28319 18652
rect 28261 18643 28319 18649
rect 28626 18640 28632 18652
rect 28684 18640 28690 18692
rect 29178 18640 29184 18692
rect 29236 18640 29242 18692
rect 29472 18680 29500 18720
rect 29546 18708 29552 18760
rect 29604 18708 29610 18760
rect 31404 18757 31432 18788
rect 31297 18751 31355 18757
rect 31297 18717 31309 18751
rect 31343 18717 31355 18751
rect 31297 18711 31355 18717
rect 31389 18751 31447 18757
rect 31389 18717 31401 18751
rect 31435 18717 31447 18751
rect 31389 18711 31447 18717
rect 31665 18751 31723 18757
rect 31665 18717 31677 18751
rect 31711 18748 31723 18751
rect 32122 18748 32128 18760
rect 31711 18720 32128 18748
rect 31711 18717 31723 18720
rect 31665 18711 31723 18717
rect 31312 18680 31340 18711
rect 32122 18708 32128 18720
rect 32180 18708 32186 18760
rect 32416 18757 32444 18788
rect 32401 18751 32459 18757
rect 32401 18717 32413 18751
rect 32447 18717 32459 18751
rect 32401 18711 32459 18717
rect 32493 18751 32551 18757
rect 32493 18717 32505 18751
rect 32539 18748 32551 18751
rect 32582 18748 32588 18760
rect 32539 18720 32588 18748
rect 32539 18717 32551 18720
rect 32493 18711 32551 18717
rect 32582 18708 32588 18720
rect 32640 18748 32646 18760
rect 32766 18748 32772 18760
rect 32640 18720 32772 18748
rect 32640 18708 32646 18720
rect 32766 18708 32772 18720
rect 32824 18748 32830 18760
rect 33060 18748 33088 18788
rect 33612 18760 33640 18788
rect 34330 18776 34336 18828
rect 34388 18776 34394 18828
rect 32824 18720 33088 18748
rect 33229 18751 33287 18757
rect 32824 18708 32830 18720
rect 33229 18717 33241 18751
rect 33275 18748 33287 18751
rect 33318 18748 33324 18760
rect 33275 18720 33324 18748
rect 33275 18717 33287 18720
rect 33229 18711 33287 18717
rect 33318 18708 33324 18720
rect 33376 18708 33382 18760
rect 33410 18708 33416 18760
rect 33468 18708 33474 18760
rect 33502 18708 33508 18760
rect 33560 18708 33566 18760
rect 33594 18708 33600 18760
rect 33652 18757 33658 18760
rect 33652 18751 33679 18757
rect 33667 18717 33679 18751
rect 33652 18711 33679 18717
rect 33652 18708 33658 18711
rect 33778 18708 33784 18760
rect 33836 18748 33842 18760
rect 34054 18748 34060 18760
rect 33836 18720 34060 18748
rect 33836 18708 33842 18720
rect 34054 18708 34060 18720
rect 34112 18708 34118 18760
rect 34149 18751 34207 18757
rect 34149 18717 34161 18751
rect 34195 18717 34207 18751
rect 34149 18711 34207 18717
rect 34425 18751 34483 18757
rect 34425 18717 34437 18751
rect 34471 18748 34483 18751
rect 34885 18751 34943 18757
rect 34885 18748 34897 18751
rect 34471 18720 34897 18748
rect 34471 18717 34483 18720
rect 34425 18711 34483 18717
rect 34885 18717 34897 18720
rect 34931 18717 34943 18751
rect 34885 18711 34943 18717
rect 32030 18680 32036 18692
rect 29472 18652 29684 18680
rect 31312 18652 32036 18680
rect 16316 18584 17356 18612
rect 17405 18615 17463 18621
rect 17405 18581 17417 18615
rect 17451 18612 17463 18615
rect 18046 18612 18052 18624
rect 17451 18584 18052 18612
rect 17451 18581 17463 18584
rect 17405 18575 17463 18581
rect 18046 18572 18052 18584
rect 18104 18572 18110 18624
rect 19705 18615 19763 18621
rect 19705 18581 19717 18615
rect 19751 18612 19763 18615
rect 19794 18612 19800 18624
rect 19751 18584 19800 18612
rect 19751 18581 19763 18584
rect 19705 18575 19763 18581
rect 19794 18572 19800 18584
rect 19852 18572 19858 18624
rect 21266 18572 21272 18624
rect 21324 18612 21330 18624
rect 22649 18615 22707 18621
rect 22649 18612 22661 18615
rect 21324 18584 22661 18612
rect 21324 18572 21330 18584
rect 22649 18581 22661 18584
rect 22695 18581 22707 18615
rect 22649 18575 22707 18581
rect 28350 18572 28356 18624
rect 28408 18612 28414 18624
rect 28537 18615 28595 18621
rect 28537 18612 28549 18615
rect 28408 18584 28549 18612
rect 28408 18572 28414 18584
rect 28537 18581 28549 18584
rect 28583 18581 28595 18615
rect 28537 18575 28595 18581
rect 29270 18572 29276 18624
rect 29328 18572 29334 18624
rect 29656 18621 29684 18652
rect 32030 18640 32036 18652
rect 32088 18640 32094 18692
rect 32309 18683 32367 18689
rect 32309 18649 32321 18683
rect 32355 18680 32367 18683
rect 32950 18680 32956 18692
rect 32355 18652 32956 18680
rect 32355 18649 32367 18652
rect 32309 18643 32367 18649
rect 32950 18640 32956 18652
rect 33008 18640 33014 18692
rect 34164 18680 34192 18711
rect 35342 18708 35348 18760
rect 35400 18748 35406 18760
rect 35437 18751 35495 18757
rect 35437 18748 35449 18751
rect 35400 18720 35449 18748
rect 35400 18708 35406 18720
rect 35437 18717 35449 18720
rect 35483 18717 35495 18751
rect 35437 18711 35495 18717
rect 36170 18708 36176 18760
rect 36228 18708 36234 18760
rect 36281 18757 36309 18856
rect 36817 18853 36829 18887
rect 36863 18853 36875 18887
rect 36817 18847 36875 18853
rect 36832 18816 36860 18847
rect 36906 18844 36912 18896
rect 36964 18884 36970 18896
rect 37752 18884 37780 18912
rect 36964 18856 37780 18884
rect 38013 18887 38071 18893
rect 36964 18844 36970 18856
rect 38013 18853 38025 18887
rect 38059 18884 38071 18887
rect 38059 18856 38240 18884
rect 38059 18853 38071 18856
rect 38013 18847 38071 18853
rect 38212 18825 38240 18856
rect 38286 18844 38292 18896
rect 38344 18884 38350 18896
rect 38657 18887 38715 18893
rect 38657 18884 38669 18887
rect 38344 18856 38669 18884
rect 38344 18844 38350 18856
rect 38657 18853 38669 18856
rect 38703 18853 38715 18887
rect 38657 18847 38715 18853
rect 38197 18819 38255 18825
rect 36832 18788 38056 18816
rect 36266 18751 36324 18757
rect 36266 18717 36278 18751
rect 36312 18717 36324 18751
rect 36266 18711 36324 18717
rect 36446 18708 36452 18760
rect 36504 18708 36510 18760
rect 36538 18708 36544 18760
rect 36596 18708 36602 18760
rect 36679 18751 36737 18757
rect 36679 18717 36691 18751
rect 36725 18748 36737 18751
rect 36725 18720 37136 18748
rect 36725 18717 36737 18720
rect 36679 18711 36737 18717
rect 33796 18652 34192 18680
rect 36464 18680 36492 18708
rect 36998 18680 37004 18692
rect 36464 18652 37004 18680
rect 29641 18615 29699 18621
rect 29641 18581 29653 18615
rect 29687 18612 29699 18615
rect 30282 18612 30288 18624
rect 29687 18584 30288 18612
rect 29687 18581 29699 18584
rect 29641 18575 29699 18581
rect 30282 18572 30288 18584
rect 30340 18572 30346 18624
rect 32490 18572 32496 18624
rect 32548 18612 32554 18624
rect 33796 18621 33824 18652
rect 36998 18640 37004 18652
rect 37056 18640 37062 18692
rect 37108 18680 37136 18720
rect 37182 18708 37188 18760
rect 37240 18748 37246 18760
rect 37369 18751 37427 18757
rect 37369 18748 37381 18751
rect 37240 18720 37381 18748
rect 37240 18708 37246 18720
rect 37369 18717 37381 18720
rect 37415 18717 37427 18751
rect 37369 18711 37427 18717
rect 37458 18708 37464 18760
rect 37516 18708 37522 18760
rect 37642 18708 37648 18760
rect 37700 18708 37706 18760
rect 37826 18708 37832 18760
rect 37884 18757 37890 18760
rect 37884 18748 37892 18757
rect 37884 18720 37929 18748
rect 37884 18711 37892 18720
rect 37884 18708 37890 18711
rect 37737 18683 37795 18689
rect 37108 18652 37412 18680
rect 37384 18624 37412 18652
rect 37737 18649 37749 18683
rect 37783 18649 37795 18683
rect 38028 18680 38056 18788
rect 38197 18785 38209 18819
rect 38243 18785 38255 18819
rect 39040 18816 39068 18924
rect 39868 18893 39896 18924
rect 40126 18912 40132 18964
rect 40184 18912 40190 18964
rect 40405 18955 40463 18961
rect 40405 18921 40417 18955
rect 40451 18952 40463 18955
rect 40494 18952 40500 18964
rect 40451 18924 40500 18952
rect 40451 18921 40463 18924
rect 40405 18915 40463 18921
rect 39853 18887 39911 18893
rect 39853 18853 39865 18887
rect 39899 18853 39911 18887
rect 40420 18884 40448 18915
rect 40494 18912 40500 18924
rect 40552 18912 40558 18964
rect 41046 18912 41052 18964
rect 41104 18912 41110 18964
rect 48222 18912 48228 18964
rect 48280 18952 48286 18964
rect 51997 18955 52055 18961
rect 51997 18952 52009 18955
rect 48280 18924 52009 18952
rect 48280 18912 48286 18924
rect 51997 18921 52009 18924
rect 52043 18952 52055 18955
rect 52454 18952 52460 18964
rect 52043 18924 52460 18952
rect 52043 18921 52055 18924
rect 51997 18915 52055 18921
rect 52454 18912 52460 18924
rect 52512 18912 52518 18964
rect 55858 18952 55864 18964
rect 53024 18924 55864 18952
rect 39853 18847 39911 18853
rect 39960 18856 40448 18884
rect 39960 18816 39988 18856
rect 40678 18844 40684 18896
rect 40736 18884 40742 18896
rect 47210 18884 47216 18896
rect 40736 18856 47216 18884
rect 40736 18844 40742 18856
rect 47210 18844 47216 18856
rect 47268 18844 47274 18896
rect 47302 18844 47308 18896
rect 47360 18884 47366 18896
rect 48593 18887 48651 18893
rect 48593 18884 48605 18887
rect 47360 18856 48605 18884
rect 47360 18844 47366 18856
rect 48593 18853 48605 18856
rect 48639 18884 48651 18887
rect 49142 18884 49148 18896
rect 48639 18856 49148 18884
rect 48639 18853 48651 18856
rect 48593 18847 48651 18853
rect 49142 18844 49148 18856
rect 49200 18844 49206 18896
rect 52086 18884 52092 18896
rect 51552 18856 52092 18884
rect 38197 18779 38255 18785
rect 38304 18788 39068 18816
rect 39224 18788 39988 18816
rect 40129 18819 40187 18825
rect 38105 18751 38163 18757
rect 38105 18717 38117 18751
rect 38151 18748 38163 18751
rect 38304 18748 38332 18788
rect 38151 18720 38332 18748
rect 38381 18751 38439 18757
rect 38151 18717 38163 18720
rect 38105 18711 38163 18717
rect 38381 18717 38393 18751
rect 38427 18717 38439 18751
rect 38381 18711 38439 18717
rect 38396 18680 38424 18711
rect 38838 18708 38844 18760
rect 38896 18708 38902 18760
rect 39022 18757 39028 18760
rect 38989 18751 39028 18757
rect 38989 18717 39001 18751
rect 38989 18711 39028 18717
rect 39022 18708 39028 18711
rect 39080 18708 39086 18760
rect 39117 18751 39175 18757
rect 39117 18717 39129 18751
rect 39163 18748 39175 18751
rect 39224 18748 39252 18788
rect 40129 18785 40141 18819
rect 40175 18816 40187 18819
rect 47228 18816 47256 18844
rect 49694 18816 49700 18828
rect 40175 18788 40816 18816
rect 47228 18788 49700 18816
rect 40175 18785 40187 18788
rect 40129 18779 40187 18785
rect 39163 18720 39252 18748
rect 39347 18751 39405 18757
rect 39163 18717 39175 18720
rect 39117 18711 39175 18717
rect 39347 18717 39359 18751
rect 39393 18748 39405 18751
rect 39574 18748 39580 18760
rect 39393 18720 39580 18748
rect 39393 18717 39405 18720
rect 39347 18711 39405 18717
rect 39574 18708 39580 18720
rect 39632 18708 39638 18760
rect 40221 18751 40279 18757
rect 40221 18717 40233 18751
rect 40267 18717 40279 18751
rect 40221 18711 40279 18717
rect 38028 18652 38424 18680
rect 37737 18643 37795 18649
rect 32677 18615 32735 18621
rect 32677 18612 32689 18615
rect 32548 18584 32689 18612
rect 32548 18572 32554 18584
rect 32677 18581 32689 18584
rect 32723 18581 32735 18615
rect 32677 18575 32735 18581
rect 33781 18615 33839 18621
rect 33781 18581 33793 18615
rect 33827 18581 33839 18615
rect 33781 18575 33839 18581
rect 33870 18572 33876 18624
rect 33928 18572 33934 18624
rect 36722 18572 36728 18624
rect 36780 18612 36786 18624
rect 37274 18612 37280 18624
rect 36780 18584 37280 18612
rect 36780 18572 36786 18584
rect 37274 18572 37280 18584
rect 37332 18572 37338 18624
rect 37366 18572 37372 18624
rect 37424 18572 37430 18624
rect 37752 18612 37780 18643
rect 39206 18640 39212 18692
rect 39264 18640 39270 18692
rect 40236 18680 40264 18711
rect 39500 18652 40264 18680
rect 39390 18612 39396 18624
rect 37752 18584 39396 18612
rect 39390 18572 39396 18584
rect 39448 18572 39454 18624
rect 39500 18621 39528 18652
rect 39485 18615 39543 18621
rect 39485 18581 39497 18615
rect 39531 18581 39543 18615
rect 40788 18612 40816 18788
rect 49694 18776 49700 18788
rect 49752 18776 49758 18828
rect 50249 18819 50307 18825
rect 50249 18785 50261 18819
rect 50295 18816 50307 18819
rect 51258 18816 51264 18828
rect 50295 18788 51264 18816
rect 50295 18785 50307 18788
rect 50249 18779 50307 18785
rect 51258 18776 51264 18788
rect 51316 18816 51322 18828
rect 51552 18816 51580 18856
rect 52086 18844 52092 18856
rect 52144 18844 52150 18896
rect 52181 18887 52239 18893
rect 52181 18853 52193 18887
rect 52227 18884 52239 18887
rect 53024 18884 53052 18924
rect 55858 18912 55864 18924
rect 55916 18912 55922 18964
rect 52227 18856 53052 18884
rect 52227 18853 52239 18856
rect 52181 18847 52239 18853
rect 51316 18788 51580 18816
rect 51316 18776 51322 18788
rect 41046 18708 41052 18760
rect 41104 18748 41110 18760
rect 41233 18751 41291 18757
rect 41233 18748 41245 18751
rect 41104 18720 41245 18748
rect 41104 18708 41110 18720
rect 41233 18717 41245 18720
rect 41279 18717 41291 18751
rect 41233 18711 41291 18717
rect 41616 18720 43484 18748
rect 40862 18640 40868 18692
rect 40920 18640 40926 18692
rect 41616 18612 41644 18720
rect 43254 18640 43260 18692
rect 43312 18640 43318 18692
rect 43456 18680 43484 18720
rect 43530 18708 43536 18760
rect 43588 18708 43594 18760
rect 43714 18708 43720 18760
rect 43772 18748 43778 18760
rect 43809 18751 43867 18757
rect 43809 18748 43821 18751
rect 43772 18720 43821 18748
rect 43772 18708 43778 18720
rect 43809 18717 43821 18720
rect 43855 18748 43867 18751
rect 45186 18748 45192 18760
rect 43855 18720 45192 18748
rect 43855 18717 43867 18720
rect 43809 18711 43867 18717
rect 45186 18708 45192 18720
rect 45244 18708 45250 18760
rect 48406 18708 48412 18760
rect 48464 18708 48470 18760
rect 48685 18751 48743 18757
rect 48685 18717 48697 18751
rect 48731 18748 48743 18751
rect 49329 18751 49387 18757
rect 49329 18748 49341 18751
rect 48731 18720 49341 18748
rect 48731 18717 48743 18720
rect 48685 18711 48743 18717
rect 49329 18717 49341 18720
rect 49375 18717 49387 18751
rect 49329 18711 49387 18717
rect 49970 18708 49976 18760
rect 50028 18708 50034 18760
rect 52196 18748 52224 18847
rect 54478 18844 54484 18896
rect 54536 18884 54542 18896
rect 54938 18884 54944 18896
rect 54536 18856 54944 18884
rect 54536 18844 54542 18856
rect 54938 18844 54944 18856
rect 54996 18844 55002 18896
rect 52270 18776 52276 18828
rect 52328 18816 52334 18828
rect 54297 18819 54355 18825
rect 54297 18816 54309 18819
rect 52328 18788 54309 18816
rect 52328 18776 52334 18788
rect 54297 18785 54309 18788
rect 54343 18816 54355 18819
rect 56410 18816 56416 18828
rect 54343 18788 56416 18816
rect 54343 18785 54355 18788
rect 54297 18779 54355 18785
rect 56410 18776 56416 18788
rect 56468 18776 56474 18828
rect 51658 18720 52224 18748
rect 54386 18708 54392 18760
rect 54444 18708 54450 18760
rect 54662 18708 54668 18760
rect 54720 18708 54726 18760
rect 44634 18680 44640 18692
rect 43456 18652 44640 18680
rect 44634 18640 44640 18652
rect 44692 18640 44698 18692
rect 50522 18640 50528 18692
rect 50580 18640 50586 18692
rect 51902 18640 51908 18692
rect 51960 18680 51966 18692
rect 51960 18652 52854 18680
rect 51960 18640 51966 18652
rect 54018 18640 54024 18692
rect 54076 18640 54082 18692
rect 40788 18584 41644 18612
rect 39485 18575 39543 18581
rect 41690 18572 41696 18624
rect 41748 18612 41754 18624
rect 42242 18612 42248 18624
rect 41748 18584 42248 18612
rect 41748 18572 41754 18584
rect 42242 18572 42248 18584
rect 42300 18612 42306 18624
rect 42521 18615 42579 18621
rect 42521 18612 42533 18615
rect 42300 18584 42533 18612
rect 42300 18572 42306 18584
rect 42521 18581 42533 18584
rect 42567 18581 42579 18615
rect 42521 18575 42579 18581
rect 43162 18572 43168 18624
rect 43220 18572 43226 18624
rect 43346 18572 43352 18624
rect 43404 18612 43410 18624
rect 48130 18612 48136 18624
rect 43404 18584 48136 18612
rect 43404 18572 43410 18584
rect 48130 18572 48136 18584
rect 48188 18572 48194 18624
rect 48225 18615 48283 18621
rect 48225 18581 48237 18615
rect 48271 18612 48283 18615
rect 48314 18612 48320 18624
rect 48271 18584 48320 18612
rect 48271 18581 48283 18584
rect 48225 18575 48283 18581
rect 48314 18572 48320 18584
rect 48372 18572 48378 18624
rect 51442 18572 51448 18624
rect 51500 18612 51506 18624
rect 52549 18615 52607 18621
rect 52549 18612 52561 18615
rect 51500 18584 52561 18612
rect 51500 18572 51506 18584
rect 52549 18581 52561 18584
rect 52595 18612 52607 18615
rect 53006 18612 53012 18624
rect 52595 18584 53012 18612
rect 52595 18581 52607 18584
rect 52549 18575 52607 18581
rect 53006 18572 53012 18584
rect 53064 18572 53070 18624
rect 54849 18615 54907 18621
rect 54849 18581 54861 18615
rect 54895 18612 54907 18615
rect 56134 18612 56140 18624
rect 54895 18584 56140 18612
rect 54895 18581 54907 18584
rect 54849 18575 54907 18581
rect 56134 18572 56140 18584
rect 56192 18572 56198 18624
rect 1104 18522 78844 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 66314 18522
rect 66366 18470 66378 18522
rect 66430 18470 66442 18522
rect 66494 18470 66506 18522
rect 66558 18470 66570 18522
rect 66622 18470 78844 18522
rect 1104 18448 78844 18470
rect 20346 18368 20352 18420
rect 20404 18408 20410 18420
rect 20441 18411 20499 18417
rect 20441 18408 20453 18411
rect 20404 18380 20453 18408
rect 20404 18368 20410 18380
rect 20441 18377 20453 18380
rect 20487 18377 20499 18411
rect 20441 18371 20499 18377
rect 21637 18411 21695 18417
rect 21637 18377 21649 18411
rect 21683 18377 21695 18411
rect 21637 18371 21695 18377
rect 21652 18340 21680 18371
rect 23842 18368 23848 18420
rect 23900 18368 23906 18420
rect 24854 18368 24860 18420
rect 24912 18408 24918 18420
rect 25041 18411 25099 18417
rect 25041 18408 25053 18411
rect 24912 18380 25053 18408
rect 24912 18368 24918 18380
rect 25041 18377 25053 18380
rect 25087 18377 25099 18411
rect 25041 18371 25099 18377
rect 25777 18411 25835 18417
rect 25777 18377 25789 18411
rect 25823 18408 25835 18411
rect 26053 18411 26111 18417
rect 25823 18380 26004 18408
rect 25823 18377 25835 18380
rect 25777 18371 25835 18377
rect 22373 18343 22431 18349
rect 22373 18340 22385 18343
rect 21652 18312 22385 18340
rect 22373 18309 22385 18312
rect 22419 18309 22431 18343
rect 22373 18303 22431 18309
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18272 9735 18275
rect 9766 18272 9772 18284
rect 9723 18244 9772 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 9858 18232 9864 18284
rect 9916 18232 9922 18284
rect 17862 18232 17868 18284
rect 17920 18272 17926 18284
rect 18815 18275 18873 18281
rect 18815 18272 18827 18275
rect 17920 18244 18827 18272
rect 17920 18232 17926 18244
rect 18815 18241 18827 18244
rect 18861 18241 18873 18275
rect 18815 18235 18873 18241
rect 18969 18275 19027 18281
rect 18969 18241 18981 18275
rect 19015 18272 19027 18275
rect 19242 18272 19248 18284
rect 19015 18244 19248 18272
rect 19015 18241 19027 18244
rect 18969 18235 19027 18241
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 20070 18232 20076 18284
rect 20128 18232 20134 18284
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18272 20315 18275
rect 20438 18272 20444 18284
rect 20303 18244 20444 18272
rect 20303 18241 20315 18244
rect 20257 18235 20315 18241
rect 20438 18232 20444 18244
rect 20496 18232 20502 18284
rect 20530 18232 20536 18284
rect 20588 18272 20594 18284
rect 20625 18275 20683 18281
rect 20625 18272 20637 18275
rect 20588 18244 20637 18272
rect 20588 18232 20594 18244
rect 20625 18241 20637 18244
rect 20671 18241 20683 18275
rect 20625 18235 20683 18241
rect 21266 18232 21272 18284
rect 21324 18232 21330 18284
rect 23860 18272 23888 18368
rect 25976 18340 26004 18380
rect 26053 18377 26065 18411
rect 26099 18408 26111 18411
rect 27522 18408 27528 18420
rect 26099 18380 27528 18408
rect 26099 18377 26111 18380
rect 26053 18371 26111 18377
rect 27522 18368 27528 18380
rect 27580 18368 27586 18420
rect 28350 18368 28356 18420
rect 28408 18368 28414 18420
rect 28626 18368 28632 18420
rect 28684 18408 28690 18420
rect 28905 18411 28963 18417
rect 28905 18408 28917 18411
rect 28684 18380 28917 18408
rect 28684 18368 28690 18380
rect 28905 18377 28917 18380
rect 28951 18408 28963 18411
rect 30742 18408 30748 18420
rect 28951 18380 30748 18408
rect 28951 18377 28963 18380
rect 28905 18371 28963 18377
rect 30742 18368 30748 18380
rect 30800 18368 30806 18420
rect 33318 18368 33324 18420
rect 33376 18408 33382 18420
rect 34790 18408 34796 18420
rect 33376 18380 34796 18408
rect 33376 18368 33382 18380
rect 34790 18368 34796 18380
rect 34848 18368 34854 18420
rect 34882 18368 34888 18420
rect 34940 18408 34946 18420
rect 34940 18380 36124 18408
rect 34940 18368 34946 18380
rect 27430 18340 27436 18352
rect 25424 18312 25820 18340
rect 25976 18312 27436 18340
rect 24305 18275 24363 18281
rect 24305 18272 24317 18275
rect 14274 18164 14280 18216
rect 14332 18164 14338 18216
rect 21361 18207 21419 18213
rect 21361 18173 21373 18207
rect 21407 18204 21419 18207
rect 21450 18204 21456 18216
rect 21407 18176 21456 18204
rect 21407 18173 21419 18176
rect 21361 18167 21419 18173
rect 21450 18164 21456 18176
rect 21508 18164 21514 18216
rect 22094 18164 22100 18216
rect 22152 18164 22158 18216
rect 18598 18096 18604 18148
rect 18656 18096 18662 18148
rect 23492 18136 23520 18258
rect 23860 18244 24317 18272
rect 24305 18241 24317 18244
rect 24351 18241 24363 18275
rect 24305 18235 24363 18241
rect 24486 18232 24492 18284
rect 24544 18232 24550 18284
rect 25225 18275 25283 18281
rect 25225 18241 25237 18275
rect 25271 18272 25283 18275
rect 25424 18272 25452 18312
rect 25271 18244 25452 18272
rect 25501 18275 25559 18281
rect 25271 18241 25283 18244
rect 25225 18235 25283 18241
rect 25501 18241 25513 18275
rect 25547 18272 25559 18275
rect 25590 18272 25596 18284
rect 25547 18244 25596 18272
rect 25547 18241 25559 18244
rect 25501 18235 25559 18241
rect 25590 18232 25596 18244
rect 25648 18232 25654 18284
rect 25682 18232 25688 18284
rect 25740 18232 25746 18284
rect 25792 18272 25820 18312
rect 27430 18300 27436 18312
rect 27488 18300 27494 18352
rect 28445 18343 28503 18349
rect 28445 18340 28457 18343
rect 27816 18312 28457 18340
rect 27816 18284 27844 18312
rect 28445 18309 28457 18312
rect 28491 18309 28503 18343
rect 29270 18340 29276 18352
rect 28445 18303 28503 18309
rect 29104 18312 29276 18340
rect 25958 18272 25964 18284
rect 25792 18244 25964 18272
rect 25958 18232 25964 18244
rect 26016 18232 26022 18284
rect 26421 18275 26479 18281
rect 26421 18241 26433 18275
rect 26467 18272 26479 18275
rect 27798 18272 27804 18284
rect 26467 18244 27804 18272
rect 26467 18241 26479 18244
rect 26421 18235 26479 18241
rect 27798 18232 27804 18244
rect 27856 18232 27862 18284
rect 28074 18232 28080 18284
rect 28132 18232 28138 18284
rect 28166 18232 28172 18284
rect 28224 18232 28230 18284
rect 28261 18275 28319 18281
rect 28261 18241 28273 18275
rect 28307 18241 28319 18275
rect 28261 18235 28319 18241
rect 28537 18275 28595 18281
rect 28537 18241 28549 18275
rect 28583 18241 28595 18275
rect 28537 18235 28595 18241
rect 24397 18207 24455 18213
rect 24397 18173 24409 18207
rect 24443 18204 24455 18207
rect 26237 18207 26295 18213
rect 26237 18204 26249 18207
rect 24443 18176 26249 18204
rect 24443 18173 24455 18176
rect 24397 18167 24455 18173
rect 26237 18173 26249 18176
rect 26283 18173 26295 18207
rect 26237 18167 26295 18173
rect 26326 18164 26332 18216
rect 26384 18164 26390 18216
rect 26510 18164 26516 18216
rect 26568 18164 26574 18216
rect 27614 18164 27620 18216
rect 27672 18204 27678 18216
rect 28276 18204 28304 18235
rect 27672 18176 28304 18204
rect 28552 18204 28580 18235
rect 28626 18232 28632 18284
rect 28684 18232 28690 18284
rect 29104 18281 29132 18312
rect 29270 18300 29276 18312
rect 29328 18340 29334 18352
rect 32214 18340 32220 18352
rect 29328 18312 32220 18340
rect 29328 18300 29334 18312
rect 32214 18300 32220 18312
rect 32272 18300 32278 18352
rect 33778 18340 33784 18352
rect 32324 18312 33784 18340
rect 29089 18275 29147 18281
rect 29089 18241 29101 18275
rect 29135 18241 29147 18275
rect 29089 18235 29147 18241
rect 30653 18275 30711 18281
rect 30653 18241 30665 18275
rect 30699 18272 30711 18275
rect 30742 18272 30748 18284
rect 30699 18244 30748 18272
rect 30699 18241 30711 18244
rect 30653 18235 30711 18241
rect 30742 18232 30748 18244
rect 30800 18232 30806 18284
rect 32030 18232 32036 18284
rect 32088 18272 32094 18284
rect 32324 18281 32352 18312
rect 33778 18300 33784 18312
rect 33836 18300 33842 18352
rect 33870 18300 33876 18352
rect 33928 18300 33934 18352
rect 35434 18300 35440 18352
rect 35492 18340 35498 18352
rect 35989 18343 36047 18349
rect 35989 18340 36001 18343
rect 35492 18312 36001 18340
rect 35492 18300 35498 18312
rect 35989 18309 36001 18312
rect 36035 18309 36047 18343
rect 36096 18340 36124 18380
rect 36170 18368 36176 18420
rect 36228 18408 36234 18420
rect 36265 18411 36323 18417
rect 36265 18408 36277 18411
rect 36228 18380 36277 18408
rect 36228 18368 36234 18380
rect 36265 18377 36277 18380
rect 36311 18377 36323 18411
rect 36265 18371 36323 18377
rect 36446 18368 36452 18420
rect 36504 18408 36510 18420
rect 36541 18411 36599 18417
rect 36541 18408 36553 18411
rect 36504 18380 36553 18408
rect 36504 18368 36510 18380
rect 36541 18377 36553 18380
rect 36587 18408 36599 18411
rect 36722 18408 36728 18420
rect 36587 18380 36728 18408
rect 36587 18377 36599 18380
rect 36541 18371 36599 18377
rect 36722 18368 36728 18380
rect 36780 18368 36786 18420
rect 36817 18411 36875 18417
rect 36817 18377 36829 18411
rect 36863 18408 36875 18411
rect 37274 18408 37280 18420
rect 36863 18380 37280 18408
rect 36863 18377 36875 18380
rect 36817 18371 36875 18377
rect 37274 18368 37280 18380
rect 37332 18368 37338 18420
rect 37461 18411 37519 18417
rect 37461 18377 37473 18411
rect 37507 18408 37519 18411
rect 37550 18408 37556 18420
rect 37507 18380 37556 18408
rect 37507 18377 37519 18380
rect 37461 18371 37519 18377
rect 37550 18368 37556 18380
rect 37608 18368 37614 18420
rect 39390 18368 39396 18420
rect 39448 18408 39454 18420
rect 40497 18411 40555 18417
rect 40497 18408 40509 18411
rect 39448 18380 40509 18408
rect 39448 18368 39454 18380
rect 40497 18377 40509 18380
rect 40543 18377 40555 18411
rect 42613 18411 42671 18417
rect 40497 18371 40555 18377
rect 40604 18380 42564 18408
rect 37645 18343 37703 18349
rect 37645 18340 37657 18343
rect 36096 18312 37657 18340
rect 35989 18303 36047 18309
rect 32309 18275 32367 18281
rect 32309 18272 32321 18275
rect 32088 18244 32321 18272
rect 32088 18232 32094 18244
rect 32309 18241 32321 18244
rect 32355 18241 32367 18275
rect 32309 18235 32367 18241
rect 32401 18275 32459 18281
rect 32401 18241 32413 18275
rect 32447 18272 32459 18275
rect 32490 18272 32496 18284
rect 32447 18244 32496 18272
rect 32447 18241 32459 18244
rect 32401 18235 32459 18241
rect 32490 18232 32496 18244
rect 32548 18232 32554 18284
rect 32674 18232 32680 18284
rect 32732 18232 32738 18284
rect 35526 18272 35532 18284
rect 35006 18244 35532 18272
rect 35526 18232 35532 18244
rect 35584 18232 35590 18284
rect 35713 18275 35771 18281
rect 35713 18241 35725 18275
rect 35759 18241 35771 18275
rect 35713 18235 35771 18241
rect 35897 18275 35955 18281
rect 35897 18241 35909 18275
rect 35943 18241 35955 18275
rect 35897 18235 35955 18241
rect 29454 18204 29460 18216
rect 28552 18176 29460 18204
rect 27672 18164 27678 18176
rect 29454 18164 29460 18176
rect 29512 18164 29518 18216
rect 33597 18207 33655 18213
rect 33597 18173 33609 18207
rect 33643 18204 33655 18207
rect 33870 18204 33876 18216
rect 33643 18176 33876 18204
rect 33643 18173 33655 18176
rect 33597 18167 33655 18173
rect 33870 18164 33876 18176
rect 33928 18164 33934 18216
rect 34882 18164 34888 18216
rect 34940 18204 34946 18216
rect 35728 18204 35756 18235
rect 34940 18176 35756 18204
rect 35912 18204 35940 18235
rect 36078 18232 36084 18284
rect 36136 18232 36142 18284
rect 36633 18275 36691 18281
rect 36633 18241 36645 18275
rect 36679 18272 36691 18275
rect 36814 18272 36820 18284
rect 36679 18244 36820 18272
rect 36679 18241 36691 18244
rect 36633 18235 36691 18241
rect 36262 18204 36268 18216
rect 35912 18176 36268 18204
rect 34940 18164 34946 18176
rect 36262 18164 36268 18176
rect 36320 18204 36326 18216
rect 36446 18204 36452 18216
rect 36320 18176 36452 18204
rect 36320 18164 36326 18176
rect 36446 18164 36452 18176
rect 36504 18164 36510 18216
rect 24854 18136 24860 18148
rect 23492 18108 24860 18136
rect 24854 18096 24860 18108
rect 24912 18096 24918 18148
rect 24946 18096 24952 18148
rect 25004 18136 25010 18148
rect 25317 18139 25375 18145
rect 25317 18136 25329 18139
rect 25004 18108 25329 18136
rect 25004 18096 25010 18108
rect 25317 18105 25329 18108
rect 25363 18105 25375 18139
rect 25317 18099 25375 18105
rect 25409 18139 25467 18145
rect 25409 18105 25421 18139
rect 25455 18136 25467 18139
rect 25498 18136 25504 18148
rect 25455 18108 25504 18136
rect 25455 18105 25467 18108
rect 25409 18099 25467 18105
rect 25498 18096 25504 18108
rect 25556 18096 25562 18148
rect 25961 18139 26019 18145
rect 25961 18105 25973 18139
rect 26007 18136 26019 18139
rect 27338 18136 27344 18148
rect 26007 18108 27344 18136
rect 26007 18105 26019 18108
rect 25961 18099 26019 18105
rect 27338 18096 27344 18108
rect 27396 18096 27402 18148
rect 35621 18139 35679 18145
rect 35621 18136 35633 18139
rect 34900 18108 35633 18136
rect 9674 18028 9680 18080
rect 9732 18028 9738 18080
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 13633 18071 13691 18077
rect 13633 18068 13645 18071
rect 13320 18040 13645 18068
rect 13320 18028 13326 18040
rect 13633 18037 13645 18040
rect 13679 18037 13691 18071
rect 13633 18031 13691 18037
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 20165 18071 20223 18077
rect 20165 18068 20177 18071
rect 20036 18040 20177 18068
rect 20036 18028 20042 18040
rect 20165 18037 20177 18040
rect 20211 18037 20223 18071
rect 20165 18031 20223 18037
rect 23014 18028 23020 18080
rect 23072 18068 23078 18080
rect 25682 18068 25688 18080
rect 23072 18040 25688 18068
rect 23072 18028 23078 18040
rect 25682 18028 25688 18040
rect 25740 18028 25746 18080
rect 27893 18071 27951 18077
rect 27893 18037 27905 18071
rect 27939 18068 27951 18071
rect 28258 18068 28264 18080
rect 27939 18040 28264 18068
rect 27939 18037 27951 18040
rect 27893 18031 27951 18037
rect 28258 18028 28264 18040
rect 28316 18028 28322 18080
rect 30469 18071 30527 18077
rect 30469 18037 30481 18071
rect 30515 18068 30527 18071
rect 30650 18068 30656 18080
rect 30515 18040 30656 18068
rect 30515 18037 30527 18040
rect 30469 18031 30527 18037
rect 30650 18028 30656 18040
rect 30708 18028 30714 18080
rect 30742 18028 30748 18080
rect 30800 18028 30806 18080
rect 32122 18028 32128 18080
rect 32180 18028 32186 18080
rect 32398 18028 32404 18080
rect 32456 18068 32462 18080
rect 32585 18071 32643 18077
rect 32585 18068 32597 18071
rect 32456 18040 32597 18068
rect 32456 18028 32462 18040
rect 32585 18037 32597 18040
rect 32631 18068 32643 18071
rect 33410 18068 33416 18080
rect 32631 18040 33416 18068
rect 32631 18037 32643 18040
rect 32585 18031 32643 18037
rect 33410 18028 33416 18040
rect 33468 18028 33474 18080
rect 34514 18028 34520 18080
rect 34572 18068 34578 18080
rect 34900 18068 34928 18108
rect 35621 18105 35633 18108
rect 35667 18136 35679 18139
rect 36648 18136 36676 18235
rect 36814 18232 36820 18244
rect 36872 18232 36878 18284
rect 37292 18281 37320 18312
rect 37645 18309 37657 18312
rect 37691 18309 37703 18343
rect 37645 18303 37703 18309
rect 37826 18300 37832 18352
rect 37884 18340 37890 18352
rect 38102 18340 38108 18352
rect 37884 18312 38108 18340
rect 37884 18300 37890 18312
rect 38102 18300 38108 18312
rect 38160 18340 38166 18352
rect 40604 18340 40632 18380
rect 38160 18312 40632 18340
rect 38160 18300 38166 18312
rect 41506 18300 41512 18352
rect 41564 18300 41570 18352
rect 42536 18340 42564 18380
rect 42613 18377 42625 18411
rect 42659 18408 42671 18411
rect 42978 18408 42984 18420
rect 42659 18380 42984 18408
rect 42659 18377 42671 18380
rect 42613 18371 42671 18377
rect 42978 18368 42984 18380
rect 43036 18368 43042 18420
rect 46842 18408 46848 18420
rect 45388 18380 46848 18408
rect 43346 18340 43352 18352
rect 42536 18312 43352 18340
rect 43346 18300 43352 18312
rect 43404 18300 43410 18352
rect 44358 18340 44364 18352
rect 44298 18312 44364 18340
rect 44358 18300 44364 18312
rect 44416 18300 44422 18352
rect 45388 18340 45416 18380
rect 46842 18368 46848 18380
rect 46900 18408 46906 18420
rect 49789 18411 49847 18417
rect 46900 18380 48084 18408
rect 46900 18368 46906 18380
rect 45296 18312 45416 18340
rect 37277 18275 37335 18281
rect 37277 18241 37289 18275
rect 37323 18241 37335 18275
rect 37734 18272 37740 18284
rect 37277 18235 37335 18241
rect 37384 18244 37740 18272
rect 36998 18164 37004 18216
rect 37056 18204 37062 18216
rect 37384 18204 37412 18244
rect 37734 18232 37740 18244
rect 37792 18272 37798 18284
rect 40678 18272 40684 18284
rect 37792 18244 40684 18272
rect 37792 18232 37798 18244
rect 40678 18232 40684 18244
rect 40736 18232 40742 18284
rect 42429 18275 42487 18281
rect 42429 18241 42441 18275
rect 42475 18272 42487 18275
rect 42702 18272 42708 18284
rect 42475 18244 42708 18272
rect 42475 18241 42487 18244
rect 42429 18235 42487 18241
rect 42702 18232 42708 18244
rect 42760 18232 42766 18284
rect 45296 18281 45324 18312
rect 48056 18281 48084 18380
rect 49789 18377 49801 18411
rect 49835 18408 49847 18411
rect 49970 18408 49976 18420
rect 49835 18380 49976 18408
rect 49835 18377 49847 18380
rect 49789 18371 49847 18377
rect 49970 18368 49976 18380
rect 50028 18408 50034 18420
rect 50028 18380 50385 18408
rect 50028 18368 50034 18380
rect 48314 18300 48320 18352
rect 48372 18300 48378 18352
rect 45281 18275 45339 18281
rect 45281 18241 45293 18275
rect 45327 18241 45339 18275
rect 48041 18275 48099 18281
rect 45281 18235 45339 18241
rect 37056 18176 37412 18204
rect 37056 18164 37062 18176
rect 37458 18164 37464 18216
rect 37516 18204 37522 18216
rect 39761 18207 39819 18213
rect 39761 18204 39773 18207
rect 37516 18176 39773 18204
rect 37516 18164 37522 18176
rect 39761 18173 39773 18176
rect 39807 18204 39819 18207
rect 40218 18204 40224 18216
rect 39807 18176 40224 18204
rect 39807 18173 39819 18176
rect 39761 18167 39819 18173
rect 40218 18164 40224 18176
rect 40276 18164 40282 18216
rect 41969 18207 42027 18213
rect 41969 18173 41981 18207
rect 42015 18204 42027 18207
rect 42015 18176 42196 18204
rect 42015 18173 42027 18176
rect 41969 18167 42027 18173
rect 35667 18108 36676 18136
rect 37093 18139 37151 18145
rect 35667 18105 35679 18108
rect 35621 18099 35679 18105
rect 37093 18105 37105 18139
rect 37139 18136 37151 18139
rect 37366 18136 37372 18148
rect 37139 18108 37372 18136
rect 37139 18105 37151 18108
rect 37093 18099 37151 18105
rect 37366 18096 37372 18108
rect 37424 18136 37430 18148
rect 38286 18136 38292 18148
rect 37424 18108 38292 18136
rect 37424 18096 37430 18108
rect 38286 18096 38292 18108
rect 38344 18136 38350 18148
rect 39298 18136 39304 18148
rect 38344 18108 39304 18136
rect 38344 18096 38350 18108
rect 39298 18096 39304 18108
rect 39356 18096 39362 18148
rect 34572 18040 34928 18068
rect 34572 18028 34578 18040
rect 35342 18028 35348 18080
rect 35400 18028 35406 18080
rect 36078 18028 36084 18080
rect 36136 18068 36142 18080
rect 37829 18071 37887 18077
rect 37829 18068 37841 18071
rect 36136 18040 37841 18068
rect 36136 18028 36142 18040
rect 37829 18037 37841 18040
rect 37875 18068 37887 18071
rect 38378 18068 38384 18080
rect 37875 18040 38384 18068
rect 37875 18037 37887 18040
rect 37829 18031 37887 18037
rect 38378 18028 38384 18040
rect 38436 18028 38442 18080
rect 38746 18028 38752 18080
rect 38804 18068 38810 18080
rect 39209 18071 39267 18077
rect 39209 18068 39221 18071
rect 38804 18040 39221 18068
rect 38804 18028 38810 18040
rect 39209 18037 39221 18040
rect 39255 18037 39267 18071
rect 42168 18068 42196 18176
rect 42242 18164 42248 18216
rect 42300 18204 42306 18216
rect 42794 18204 42800 18216
rect 42300 18176 42800 18204
rect 42300 18164 42306 18176
rect 42794 18164 42800 18176
rect 42852 18164 42858 18216
rect 43070 18164 43076 18216
rect 43128 18164 43134 18216
rect 45554 18164 45560 18216
rect 45612 18164 45618 18216
rect 46676 18204 46704 18258
rect 48041 18241 48053 18275
rect 48087 18241 48099 18275
rect 48041 18235 48099 18241
rect 48314 18204 48320 18216
rect 46676 18176 48320 18204
rect 48314 18164 48320 18176
rect 48372 18204 48378 18216
rect 49436 18204 49464 18258
rect 50246 18232 50252 18284
rect 50304 18232 50310 18284
rect 50357 18281 50385 18380
rect 50522 18368 50528 18420
rect 50580 18408 50586 18420
rect 50985 18411 51043 18417
rect 50985 18408 50997 18411
rect 50580 18380 50997 18408
rect 50580 18368 50586 18380
rect 50985 18377 50997 18380
rect 51031 18377 51043 18411
rect 50985 18371 51043 18377
rect 54018 18368 54024 18420
rect 54076 18408 54082 18420
rect 54205 18411 54263 18417
rect 54205 18408 54217 18411
rect 54076 18380 54217 18408
rect 54076 18368 54082 18380
rect 54205 18377 54217 18380
rect 54251 18377 54263 18411
rect 56597 18411 56655 18417
rect 56597 18408 56609 18411
rect 54205 18371 54263 18377
rect 55876 18380 56609 18408
rect 55876 18352 55904 18380
rect 56597 18377 56609 18380
rect 56643 18377 56655 18411
rect 56597 18371 56655 18377
rect 50617 18343 50675 18349
rect 50617 18309 50629 18343
rect 50663 18340 50675 18343
rect 51442 18340 51448 18352
rect 50663 18312 51448 18340
rect 50663 18309 50675 18312
rect 50617 18303 50675 18309
rect 51442 18300 51448 18312
rect 51500 18300 51506 18352
rect 54110 18340 54116 18352
rect 53024 18312 54116 18340
rect 53024 18284 53052 18312
rect 54110 18300 54116 18312
rect 54168 18300 54174 18352
rect 55858 18340 55864 18352
rect 55706 18312 55864 18340
rect 55858 18300 55864 18312
rect 55916 18300 55922 18352
rect 56134 18300 56140 18352
rect 56192 18300 56198 18352
rect 50342 18275 50400 18281
rect 50342 18241 50354 18275
rect 50388 18241 50400 18275
rect 50342 18235 50400 18241
rect 48372 18176 49464 18204
rect 50357 18204 50385 18235
rect 50430 18232 50436 18284
rect 50488 18272 50494 18284
rect 50798 18281 50804 18284
rect 50525 18275 50583 18281
rect 50525 18272 50537 18275
rect 50488 18244 50537 18272
rect 50488 18232 50494 18244
rect 50525 18241 50537 18244
rect 50571 18241 50583 18275
rect 50525 18235 50583 18241
rect 50755 18275 50804 18281
rect 50755 18241 50767 18275
rect 50801 18241 50804 18275
rect 50755 18235 50804 18241
rect 50798 18232 50804 18235
rect 50856 18232 50862 18284
rect 51169 18275 51227 18281
rect 51169 18272 51181 18275
rect 50908 18244 51181 18272
rect 50614 18204 50620 18216
rect 50357 18176 50620 18204
rect 48372 18164 48378 18176
rect 42886 18068 42892 18080
rect 42168 18040 42892 18068
rect 39209 18031 39267 18037
rect 42886 18028 42892 18040
rect 42944 18028 42950 18080
rect 44542 18028 44548 18080
rect 44600 18028 44606 18080
rect 47026 18028 47032 18080
rect 47084 18028 47090 18080
rect 49436 18068 49464 18176
rect 50614 18164 50620 18176
rect 50672 18164 50678 18216
rect 50908 18145 50936 18244
rect 51169 18241 51181 18244
rect 51215 18241 51227 18275
rect 51169 18235 51227 18241
rect 52454 18232 52460 18284
rect 52512 18232 52518 18284
rect 53006 18232 53012 18284
rect 53064 18232 53070 18284
rect 54018 18232 54024 18284
rect 54076 18232 54082 18284
rect 56410 18232 56416 18284
rect 56468 18232 56474 18284
rect 51445 18207 51503 18213
rect 51445 18173 51457 18207
rect 51491 18204 51503 18207
rect 51813 18207 51871 18213
rect 51813 18204 51825 18207
rect 51491 18176 51825 18204
rect 51491 18173 51503 18176
rect 51445 18167 51503 18173
rect 51813 18173 51825 18176
rect 51859 18173 51871 18207
rect 51813 18167 51871 18173
rect 53653 18207 53711 18213
rect 53653 18173 53665 18207
rect 53699 18204 53711 18207
rect 53745 18207 53803 18213
rect 53745 18204 53757 18207
rect 53699 18176 53757 18204
rect 53699 18173 53711 18176
rect 53653 18167 53711 18173
rect 53745 18173 53757 18176
rect 53791 18173 53803 18207
rect 53745 18167 53803 18173
rect 53837 18207 53895 18213
rect 53837 18173 53849 18207
rect 53883 18204 53895 18207
rect 54478 18204 54484 18216
rect 53883 18176 54484 18204
rect 53883 18173 53895 18176
rect 53837 18167 53895 18173
rect 50893 18139 50951 18145
rect 50893 18105 50905 18139
rect 50939 18105 50951 18139
rect 51902 18136 51908 18148
rect 50893 18099 50951 18105
rect 51046 18108 51908 18136
rect 51046 18068 51074 18108
rect 51902 18096 51908 18108
rect 51960 18096 51966 18148
rect 49436 18040 51074 18068
rect 51350 18028 51356 18080
rect 51408 18068 51414 18080
rect 53852 18068 53880 18167
rect 54478 18164 54484 18176
rect 54536 18164 54542 18216
rect 51408 18040 53880 18068
rect 51408 18028 51414 18040
rect 53926 18028 53932 18080
rect 53984 18068 53990 18080
rect 54386 18068 54392 18080
rect 53984 18040 54392 18068
rect 53984 18028 53990 18040
rect 54386 18028 54392 18040
rect 54444 18068 54450 18080
rect 54665 18071 54723 18077
rect 54665 18068 54677 18071
rect 54444 18040 54677 18068
rect 54444 18028 54450 18040
rect 54665 18037 54677 18040
rect 54711 18037 54723 18071
rect 54665 18031 54723 18037
rect 1104 17978 78844 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 78844 17978
rect 1104 17904 78844 17926
rect 22094 17864 22100 17876
rect 18248 17836 22100 17864
rect 16206 17756 16212 17808
rect 16264 17796 16270 17808
rect 16264 17768 16436 17796
rect 16264 17756 16270 17768
rect 10686 17688 10692 17740
rect 10744 17688 10750 17740
rect 13262 17688 13268 17740
rect 13320 17688 13326 17740
rect 13449 17731 13507 17737
rect 13449 17697 13461 17731
rect 13495 17728 13507 17731
rect 15102 17728 15108 17740
rect 13495 17700 15108 17728
rect 13495 17697 13507 17700
rect 13449 17691 13507 17697
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 9490 17620 9496 17672
rect 9548 17660 9554 17672
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 9548 17632 10425 17660
rect 9548 17620 9554 17632
rect 10413 17629 10425 17632
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 12710 17620 12716 17672
rect 12768 17660 12774 17672
rect 14461 17663 14519 17669
rect 14461 17660 14473 17663
rect 12768 17632 14473 17660
rect 12768 17620 12774 17632
rect 14461 17629 14473 17632
rect 14507 17629 14519 17663
rect 16408 17660 16436 17768
rect 16482 17688 16488 17740
rect 16540 17728 16546 17740
rect 18248 17737 18276 17836
rect 22094 17824 22100 17836
rect 22152 17824 22158 17876
rect 26510 17824 26516 17876
rect 26568 17864 26574 17876
rect 27065 17867 27123 17873
rect 27065 17864 27077 17867
rect 26568 17836 27077 17864
rect 26568 17824 26574 17836
rect 27065 17833 27077 17836
rect 27111 17833 27123 17867
rect 27065 17827 27123 17833
rect 29730 17824 29736 17876
rect 29788 17864 29794 17876
rect 30101 17867 30159 17873
rect 30101 17864 30113 17867
rect 29788 17836 30113 17864
rect 29788 17824 29794 17836
rect 30101 17833 30113 17836
rect 30147 17833 30159 17867
rect 30101 17827 30159 17833
rect 30561 17867 30619 17873
rect 30561 17833 30573 17867
rect 30607 17864 30619 17867
rect 30742 17864 30748 17876
rect 30607 17836 30748 17864
rect 30607 17833 30619 17836
rect 30561 17827 30619 17833
rect 30742 17824 30748 17836
rect 30800 17864 30806 17876
rect 31386 17864 31392 17876
rect 30800 17836 31392 17864
rect 30800 17824 30806 17836
rect 31386 17824 31392 17836
rect 31444 17824 31450 17876
rect 32674 17824 32680 17876
rect 32732 17864 32738 17876
rect 32861 17867 32919 17873
rect 32861 17864 32873 17867
rect 32732 17836 32873 17864
rect 32732 17824 32738 17836
rect 32861 17833 32873 17836
rect 32907 17864 32919 17867
rect 32950 17864 32956 17876
rect 32907 17836 32956 17864
rect 32907 17833 32919 17836
rect 32861 17827 32919 17833
rect 32950 17824 32956 17836
rect 33008 17824 33014 17876
rect 33042 17824 33048 17876
rect 33100 17864 33106 17876
rect 33505 17867 33563 17873
rect 33505 17864 33517 17867
rect 33100 17836 33517 17864
rect 33100 17824 33106 17836
rect 33505 17833 33517 17836
rect 33551 17833 33563 17867
rect 33505 17827 33563 17833
rect 19334 17796 19340 17808
rect 18340 17768 19340 17796
rect 18233 17731 18291 17737
rect 18233 17728 18245 17731
rect 16540 17700 18245 17728
rect 16540 17688 16546 17700
rect 18233 17697 18245 17700
rect 18279 17697 18291 17731
rect 18233 17691 18291 17697
rect 16853 17663 16911 17669
rect 16853 17660 16865 17663
rect 16408 17632 16865 17660
rect 14461 17623 14519 17629
rect 16853 17629 16865 17632
rect 16899 17629 16911 17663
rect 16853 17623 16911 17629
rect 17494 17620 17500 17672
rect 17552 17660 17558 17672
rect 18340 17660 18368 17768
rect 19334 17756 19340 17768
rect 19392 17756 19398 17808
rect 20530 17756 20536 17808
rect 20588 17756 20594 17808
rect 20625 17799 20683 17805
rect 20625 17765 20637 17799
rect 20671 17765 20683 17799
rect 20625 17759 20683 17765
rect 18414 17688 18420 17740
rect 18472 17728 18478 17740
rect 18693 17731 18751 17737
rect 18693 17728 18705 17731
rect 18472 17700 18705 17728
rect 18472 17688 18478 17700
rect 18693 17697 18705 17700
rect 18739 17697 18751 17731
rect 18693 17691 18751 17697
rect 19978 17688 19984 17740
rect 20036 17728 20042 17740
rect 20640 17728 20668 17759
rect 21450 17756 21456 17808
rect 21508 17756 21514 17808
rect 25590 17756 25596 17808
rect 25648 17796 25654 17808
rect 25685 17799 25743 17805
rect 25685 17796 25697 17799
rect 25648 17768 25697 17796
rect 25648 17756 25654 17768
rect 25685 17765 25697 17768
rect 25731 17765 25743 17799
rect 31018 17796 31024 17808
rect 25685 17759 25743 17765
rect 28092 17768 31024 17796
rect 20036 17700 20668 17728
rect 20717 17731 20775 17737
rect 20036 17688 20042 17700
rect 20717 17697 20729 17731
rect 20763 17697 20775 17731
rect 20717 17691 20775 17697
rect 26973 17731 27031 17737
rect 26973 17697 26985 17731
rect 27019 17728 27031 17731
rect 27019 17700 27384 17728
rect 27019 17697 27031 17700
rect 26973 17691 27031 17697
rect 17552 17632 18368 17660
rect 18509 17663 18567 17669
rect 17552 17620 17558 17632
rect 18509 17629 18521 17663
rect 18555 17660 18567 17663
rect 18598 17660 18604 17672
rect 18555 17632 18604 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 11146 17552 11152 17604
rect 11204 17552 11210 17604
rect 13173 17595 13231 17601
rect 13173 17592 13185 17595
rect 12176 17564 13185 17592
rect 12176 17533 12204 17564
rect 13173 17561 13185 17564
rect 13219 17592 13231 17595
rect 14182 17592 14188 17604
rect 13219 17564 14188 17592
rect 13219 17561 13231 17564
rect 13173 17555 13231 17561
rect 14182 17552 14188 17564
rect 14240 17552 14246 17604
rect 14734 17552 14740 17604
rect 14792 17552 14798 17604
rect 14936 17564 15226 17592
rect 14936 17536 14964 17564
rect 18138 17552 18144 17604
rect 18196 17592 18202 17604
rect 18524 17592 18552 17623
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 20165 17663 20223 17669
rect 20165 17660 20177 17663
rect 20128 17632 20177 17660
rect 20128 17620 20134 17632
rect 20165 17629 20177 17632
rect 20211 17660 20223 17663
rect 20622 17660 20628 17672
rect 20211 17632 20628 17660
rect 20211 17629 20223 17632
rect 20165 17623 20223 17629
rect 20622 17620 20628 17632
rect 20680 17620 20686 17672
rect 18196 17564 18552 17592
rect 18196 17552 18202 17564
rect 20438 17552 20444 17604
rect 20496 17592 20502 17604
rect 20732 17592 20760 17691
rect 21637 17663 21695 17669
rect 21637 17629 21649 17663
rect 21683 17660 21695 17663
rect 22094 17660 22100 17672
rect 21683 17632 22100 17660
rect 21683 17629 21695 17632
rect 21637 17623 21695 17629
rect 22094 17620 22100 17632
rect 22152 17620 22158 17672
rect 25958 17620 25964 17672
rect 26016 17620 26022 17672
rect 26053 17663 26111 17669
rect 26053 17629 26065 17663
rect 26099 17660 26111 17663
rect 26234 17660 26240 17672
rect 26099 17632 26240 17660
rect 26099 17629 26111 17632
rect 26053 17623 26111 17629
rect 26234 17620 26240 17632
rect 26292 17620 26298 17672
rect 27246 17620 27252 17672
rect 27304 17620 27310 17672
rect 27356 17669 27384 17700
rect 27341 17663 27399 17669
rect 27341 17629 27353 17663
rect 27387 17629 27399 17663
rect 27341 17623 27399 17629
rect 20496 17564 20760 17592
rect 21821 17595 21879 17601
rect 20496 17552 20502 17564
rect 21821 17561 21833 17595
rect 21867 17561 21879 17595
rect 25976 17592 26004 17620
rect 26970 17592 26976 17604
rect 25976 17564 26976 17592
rect 21821 17555 21879 17561
rect 12161 17527 12219 17533
rect 12161 17493 12173 17527
rect 12207 17493 12219 17527
rect 12161 17487 12219 17493
rect 12434 17484 12440 17536
rect 12492 17524 12498 17536
rect 12805 17527 12863 17533
rect 12805 17524 12817 17527
rect 12492 17496 12817 17524
rect 12492 17484 12498 17496
rect 12805 17493 12817 17496
rect 12851 17493 12863 17527
rect 12805 17487 12863 17493
rect 14918 17484 14924 17536
rect 14976 17484 14982 17536
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 16301 17527 16359 17533
rect 16301 17524 16313 17527
rect 15620 17496 16313 17524
rect 15620 17484 15626 17496
rect 16301 17493 16313 17496
rect 16347 17493 16359 17527
rect 16301 17487 16359 17493
rect 20990 17484 20996 17536
rect 21048 17524 21054 17536
rect 21836 17524 21864 17555
rect 26970 17552 26976 17564
rect 27028 17552 27034 17604
rect 27356 17592 27384 17623
rect 27430 17620 27436 17672
rect 27488 17660 27494 17672
rect 28092 17669 28120 17768
rect 31018 17756 31024 17768
rect 31076 17756 31082 17808
rect 28534 17728 28540 17740
rect 28184 17700 28540 17728
rect 27525 17663 27583 17669
rect 27525 17660 27537 17663
rect 27488 17632 27537 17660
rect 27488 17620 27494 17632
rect 27525 17629 27537 17632
rect 27571 17629 27583 17663
rect 27525 17623 27583 17629
rect 27617 17663 27675 17669
rect 27617 17629 27629 17663
rect 27663 17660 27675 17663
rect 27801 17663 27859 17669
rect 27801 17660 27813 17663
rect 27663 17632 27813 17660
rect 27663 17629 27675 17632
rect 27617 17623 27675 17629
rect 27801 17629 27813 17632
rect 27847 17629 27859 17663
rect 27801 17623 27859 17629
rect 27985 17663 28043 17669
rect 27985 17629 27997 17663
rect 28031 17629 28043 17663
rect 27985 17623 28043 17629
rect 28077 17663 28135 17669
rect 28077 17629 28089 17663
rect 28123 17629 28135 17663
rect 28077 17623 28135 17629
rect 27706 17592 27712 17604
rect 27356 17564 27712 17592
rect 27706 17552 27712 17564
rect 27764 17552 27770 17604
rect 28000 17592 28028 17623
rect 28184 17592 28212 17700
rect 28534 17688 28540 17700
rect 28592 17688 28598 17740
rect 30650 17728 30656 17740
rect 29932 17700 30656 17728
rect 28258 17620 28264 17672
rect 28316 17620 28322 17672
rect 28350 17620 28356 17672
rect 28408 17620 28414 17672
rect 29932 17669 29960 17700
rect 30650 17688 30656 17700
rect 30708 17688 30714 17740
rect 31110 17688 31116 17740
rect 31168 17688 31174 17740
rect 31389 17731 31447 17737
rect 31389 17697 31401 17731
rect 31435 17728 31447 17731
rect 32122 17728 32128 17740
rect 31435 17700 32128 17728
rect 31435 17697 31447 17700
rect 31389 17691 31447 17697
rect 32122 17688 32128 17700
rect 32180 17688 32186 17740
rect 29641 17663 29699 17669
rect 29641 17629 29653 17663
rect 29687 17629 29699 17663
rect 29641 17623 29699 17629
rect 29917 17663 29975 17669
rect 29917 17629 29929 17663
rect 29963 17629 29975 17663
rect 29917 17623 29975 17629
rect 28000 17564 28212 17592
rect 28276 17592 28304 17620
rect 28902 17592 28908 17604
rect 28276 17564 28908 17592
rect 28902 17552 28908 17564
rect 28960 17552 28966 17604
rect 21048 17496 21864 17524
rect 21048 17484 21054 17496
rect 27246 17484 27252 17536
rect 27304 17524 27310 17536
rect 29656 17524 29684 17623
rect 30926 17620 30932 17672
rect 30984 17660 30990 17672
rect 33321 17663 33379 17669
rect 30984 17632 31156 17660
rect 30984 17620 30990 17632
rect 31128 17604 31156 17632
rect 33321 17629 33333 17663
rect 33367 17660 33379 17663
rect 33367 17632 33456 17660
rect 33367 17629 33379 17632
rect 33321 17623 33379 17629
rect 30653 17595 30711 17601
rect 30653 17561 30665 17595
rect 30699 17592 30711 17595
rect 31018 17592 31024 17604
rect 30699 17564 31024 17592
rect 30699 17561 30711 17564
rect 30653 17555 30711 17561
rect 31018 17552 31024 17564
rect 31076 17552 31082 17604
rect 31110 17552 31116 17604
rect 31168 17592 31174 17604
rect 33045 17595 33103 17601
rect 33045 17592 33057 17595
rect 31168 17564 31878 17592
rect 32692 17564 33057 17592
rect 31168 17552 31174 17564
rect 27304 17496 29684 17524
rect 29733 17527 29791 17533
rect 27304 17484 27310 17496
rect 29733 17493 29745 17527
rect 29779 17524 29791 17527
rect 29822 17524 29828 17536
rect 29779 17496 29828 17524
rect 29779 17493 29791 17496
rect 29733 17487 29791 17493
rect 29822 17484 29828 17496
rect 29880 17524 29886 17536
rect 30193 17527 30251 17533
rect 30193 17524 30205 17527
rect 29880 17496 30205 17524
rect 29880 17484 29886 17496
rect 30193 17493 30205 17496
rect 30239 17493 30251 17527
rect 30193 17487 30251 17493
rect 30742 17484 30748 17536
rect 30800 17524 30806 17536
rect 32692 17524 32720 17564
rect 33045 17561 33057 17564
rect 33091 17561 33103 17595
rect 33045 17555 33103 17561
rect 30800 17496 32720 17524
rect 30800 17484 30806 17496
rect 33134 17484 33140 17536
rect 33192 17484 33198 17536
rect 33318 17484 33324 17536
rect 33376 17524 33382 17536
rect 33428 17524 33456 17632
rect 33520 17592 33548 17827
rect 33778 17824 33784 17876
rect 33836 17864 33842 17876
rect 34422 17864 34428 17876
rect 33836 17836 34428 17864
rect 33836 17824 33842 17836
rect 34422 17824 34428 17836
rect 34480 17824 34486 17876
rect 37550 17864 37556 17876
rect 36648 17836 37556 17864
rect 36446 17756 36452 17808
rect 36504 17756 36510 17808
rect 35342 17728 35348 17740
rect 34992 17700 35348 17728
rect 33594 17620 33600 17672
rect 33652 17660 33658 17672
rect 34992 17669 35020 17700
rect 35342 17688 35348 17700
rect 35400 17688 35406 17740
rect 34885 17663 34943 17669
rect 34885 17660 34897 17663
rect 33652 17632 34897 17660
rect 33652 17620 33658 17632
rect 34885 17629 34897 17632
rect 34931 17629 34943 17663
rect 34885 17623 34943 17629
rect 34977 17663 35035 17669
rect 34977 17629 34989 17663
rect 35023 17629 35035 17663
rect 34977 17623 35035 17629
rect 35253 17663 35311 17669
rect 35253 17629 35265 17663
rect 35299 17660 35311 17663
rect 35434 17660 35440 17672
rect 35299 17632 35440 17660
rect 35299 17629 35311 17632
rect 35253 17623 35311 17629
rect 35434 17620 35440 17632
rect 35492 17620 35498 17672
rect 36648 17669 36676 17836
rect 37550 17824 37556 17836
rect 37608 17824 37614 17876
rect 38838 17824 38844 17876
rect 38896 17864 38902 17876
rect 40862 17864 40868 17876
rect 38896 17836 40868 17864
rect 38896 17824 38902 17836
rect 40862 17824 40868 17836
rect 40920 17824 40926 17876
rect 41322 17824 41328 17876
rect 41380 17864 41386 17876
rect 42242 17864 42248 17876
rect 41380 17836 42248 17864
rect 41380 17824 41386 17836
rect 42242 17824 42248 17836
rect 42300 17824 42306 17876
rect 43438 17824 43444 17876
rect 43496 17864 43502 17876
rect 43625 17867 43683 17873
rect 43625 17864 43637 17867
rect 43496 17836 43637 17864
rect 43496 17824 43502 17836
rect 43625 17833 43637 17836
rect 43671 17833 43683 17867
rect 43625 17827 43683 17833
rect 45554 17824 45560 17876
rect 45612 17864 45618 17876
rect 45833 17867 45891 17873
rect 45833 17864 45845 17867
rect 45612 17836 45845 17864
rect 45612 17824 45618 17836
rect 45833 17833 45845 17836
rect 45879 17833 45891 17867
rect 45833 17827 45891 17833
rect 46124 17836 47440 17864
rect 37274 17796 37280 17808
rect 36924 17768 37280 17796
rect 36633 17663 36691 17669
rect 36633 17629 36645 17663
rect 36679 17629 36691 17663
rect 36633 17623 36691 17629
rect 36817 17663 36875 17669
rect 36817 17629 36829 17663
rect 36863 17660 36875 17663
rect 36924 17660 36952 17768
rect 37274 17756 37280 17768
rect 37332 17796 37338 17808
rect 38470 17796 38476 17808
rect 37332 17768 38476 17796
rect 37332 17756 37338 17768
rect 38470 17756 38476 17768
rect 38528 17756 38534 17808
rect 39390 17756 39396 17808
rect 39448 17796 39454 17808
rect 39448 17768 41736 17796
rect 39448 17756 39454 17768
rect 37458 17728 37464 17740
rect 37016 17700 37464 17728
rect 37016 17669 37044 17700
rect 37458 17688 37464 17700
rect 37516 17688 37522 17740
rect 38562 17688 38568 17740
rect 38620 17728 38626 17740
rect 40862 17728 40868 17740
rect 38620 17700 40868 17728
rect 38620 17688 38626 17700
rect 40862 17688 40868 17700
rect 40920 17728 40926 17740
rect 41322 17728 41328 17740
rect 40920 17700 41328 17728
rect 40920 17688 40926 17700
rect 41322 17688 41328 17700
rect 41380 17688 41386 17740
rect 36863 17632 36952 17660
rect 37001 17663 37059 17669
rect 36863 17629 36875 17632
rect 36817 17623 36875 17629
rect 37001 17629 37013 17663
rect 37047 17629 37059 17663
rect 37001 17623 37059 17629
rect 37093 17663 37151 17669
rect 37093 17629 37105 17663
rect 37139 17660 37151 17663
rect 37366 17660 37372 17672
rect 37139 17632 37372 17660
rect 37139 17629 37151 17632
rect 37093 17623 37151 17629
rect 35069 17595 35127 17601
rect 35069 17592 35081 17595
rect 33520 17564 35081 17592
rect 35069 17561 35081 17564
rect 35115 17561 35127 17595
rect 35069 17555 35127 17561
rect 36538 17552 36544 17604
rect 36596 17592 36602 17604
rect 36725 17595 36783 17601
rect 36725 17592 36737 17595
rect 36596 17564 36737 17592
rect 36596 17552 36602 17564
rect 36725 17561 36737 17564
rect 36771 17561 36783 17595
rect 36725 17555 36783 17561
rect 33778 17524 33784 17536
rect 33376 17496 33784 17524
rect 33376 17484 33382 17496
rect 33778 17484 33784 17496
rect 33836 17484 33842 17536
rect 34514 17484 34520 17536
rect 34572 17524 34578 17536
rect 34701 17527 34759 17533
rect 34701 17524 34713 17527
rect 34572 17496 34713 17524
rect 34572 17484 34578 17496
rect 34701 17493 34713 17496
rect 34747 17493 34759 17527
rect 34701 17487 34759 17493
rect 35342 17484 35348 17536
rect 35400 17524 35406 17536
rect 35437 17527 35495 17533
rect 35437 17524 35449 17527
rect 35400 17496 35449 17524
rect 35400 17484 35406 17496
rect 35437 17493 35449 17496
rect 35483 17524 35495 17527
rect 35526 17524 35532 17536
rect 35483 17496 35532 17524
rect 35483 17493 35495 17496
rect 35437 17487 35495 17493
rect 35526 17484 35532 17496
rect 35584 17484 35590 17536
rect 36354 17484 36360 17536
rect 36412 17524 36418 17536
rect 37108 17524 37136 17623
rect 37366 17620 37372 17632
rect 37424 17620 37430 17672
rect 38933 17663 38991 17669
rect 38933 17629 38945 17663
rect 38979 17660 38991 17663
rect 39022 17660 39028 17672
rect 38979 17632 39028 17660
rect 38979 17629 38991 17632
rect 38933 17623 38991 17629
rect 39022 17620 39028 17632
rect 39080 17620 39086 17672
rect 40034 17669 40040 17672
rect 39209 17663 39267 17669
rect 39209 17629 39221 17663
rect 39255 17629 39267 17663
rect 39209 17623 39267 17629
rect 39853 17663 39911 17669
rect 39853 17629 39865 17663
rect 39899 17629 39911 17663
rect 39853 17623 39911 17629
rect 40001 17663 40040 17669
rect 40001 17629 40013 17663
rect 40001 17623 40040 17629
rect 38194 17552 38200 17604
rect 38252 17592 38258 17604
rect 39224 17592 39252 17623
rect 39666 17592 39672 17604
rect 38252 17564 39672 17592
rect 38252 17552 38258 17564
rect 39666 17552 39672 17564
rect 39724 17552 39730 17604
rect 36412 17496 37136 17524
rect 36412 17484 36418 17496
rect 37274 17484 37280 17536
rect 37332 17484 37338 17536
rect 37366 17484 37372 17536
rect 37424 17524 37430 17536
rect 37461 17527 37519 17533
rect 37461 17524 37473 17527
rect 37424 17496 37473 17524
rect 37424 17484 37430 17496
rect 37461 17493 37473 17496
rect 37507 17493 37519 17527
rect 37461 17487 37519 17493
rect 39022 17484 39028 17536
rect 39080 17524 39086 17536
rect 39868 17524 39896 17623
rect 40034 17620 40040 17623
rect 40092 17620 40098 17672
rect 40218 17620 40224 17672
rect 40276 17620 40282 17672
rect 40310 17620 40316 17672
rect 40368 17669 40374 17672
rect 40368 17660 40376 17669
rect 40954 17660 40960 17672
rect 40368 17632 40413 17660
rect 40512 17632 40960 17660
rect 40368 17623 40376 17632
rect 40368 17620 40374 17623
rect 40129 17595 40187 17601
rect 40129 17561 40141 17595
rect 40175 17592 40187 17595
rect 40512 17592 40540 17632
rect 40954 17620 40960 17632
rect 41012 17620 41018 17672
rect 41708 17669 41736 17768
rect 42426 17688 42432 17740
rect 42484 17688 42490 17740
rect 42518 17688 42524 17740
rect 42576 17728 42582 17740
rect 42576 17700 42748 17728
rect 42576 17688 42582 17700
rect 41693 17663 41751 17669
rect 41693 17629 41705 17663
rect 41739 17629 41751 17663
rect 41693 17623 41751 17629
rect 42245 17663 42303 17669
rect 42245 17629 42257 17663
rect 42291 17660 42303 17663
rect 42337 17663 42395 17669
rect 42337 17660 42349 17663
rect 42291 17632 42349 17660
rect 42291 17629 42303 17632
rect 42245 17623 42303 17629
rect 42337 17629 42349 17632
rect 42383 17629 42395 17663
rect 42337 17623 42395 17629
rect 40175 17564 40540 17592
rect 40175 17561 40187 17564
rect 40129 17555 40187 17561
rect 40586 17552 40592 17604
rect 40644 17592 40650 17604
rect 41414 17592 41420 17604
rect 40644 17564 41420 17592
rect 40644 17552 40650 17564
rect 41414 17552 41420 17564
rect 41472 17552 41478 17604
rect 41708 17592 41736 17623
rect 42610 17620 42616 17672
rect 42668 17620 42674 17672
rect 42720 17669 42748 17700
rect 42886 17688 42892 17740
rect 42944 17688 42950 17740
rect 44542 17688 44548 17740
rect 44600 17728 44606 17740
rect 44729 17731 44787 17737
rect 44729 17728 44741 17731
rect 44600 17700 44741 17728
rect 44600 17688 44606 17700
rect 44729 17697 44741 17700
rect 44775 17697 44787 17731
rect 44729 17691 44787 17697
rect 45741 17731 45799 17737
rect 45741 17697 45753 17731
rect 45787 17728 45799 17731
rect 46124 17728 46152 17836
rect 46290 17756 46296 17808
rect 46348 17796 46354 17808
rect 47302 17796 47308 17808
rect 46348 17768 47308 17796
rect 46348 17756 46354 17768
rect 47302 17756 47308 17768
rect 47360 17756 47366 17808
rect 47412 17796 47440 17836
rect 47578 17824 47584 17876
rect 47636 17864 47642 17876
rect 47854 17864 47860 17876
rect 47636 17836 47860 17864
rect 47636 17824 47642 17836
rect 47854 17824 47860 17836
rect 47912 17824 47918 17876
rect 48406 17824 48412 17876
rect 48464 17824 48470 17876
rect 50798 17824 50804 17876
rect 50856 17864 50862 17876
rect 51074 17864 51080 17876
rect 50856 17836 51080 17864
rect 50856 17824 50862 17836
rect 51074 17824 51080 17836
rect 51132 17864 51138 17876
rect 51721 17867 51779 17873
rect 51721 17864 51733 17867
rect 51132 17836 51733 17864
rect 51132 17824 51138 17836
rect 51721 17833 51733 17836
rect 51767 17864 51779 17867
rect 52546 17864 52552 17876
rect 51767 17836 52552 17864
rect 51767 17833 51779 17836
rect 51721 17827 51779 17833
rect 52546 17824 52552 17836
rect 52604 17864 52610 17876
rect 53190 17864 53196 17876
rect 52604 17836 53196 17864
rect 52604 17824 52610 17836
rect 53190 17824 53196 17836
rect 53248 17824 53254 17876
rect 53377 17867 53435 17873
rect 53377 17833 53389 17867
rect 53423 17864 53435 17867
rect 54018 17864 54024 17876
rect 53423 17836 54024 17864
rect 53423 17833 53435 17836
rect 53377 17827 53435 17833
rect 54018 17824 54024 17836
rect 54076 17824 54082 17876
rect 54573 17867 54631 17873
rect 54573 17833 54585 17867
rect 54619 17864 54631 17867
rect 54662 17864 54668 17876
rect 54619 17836 54668 17864
rect 54619 17833 54631 17836
rect 54573 17827 54631 17833
rect 54662 17824 54668 17836
rect 54720 17824 54726 17876
rect 48774 17796 48780 17808
rect 47412 17768 48780 17796
rect 48774 17756 48780 17768
rect 48832 17756 48838 17808
rect 50246 17756 50252 17808
rect 50304 17796 50310 17808
rect 50304 17768 51672 17796
rect 50304 17756 50310 17768
rect 45787 17700 46152 17728
rect 45787 17697 45799 17700
rect 45741 17691 45799 17697
rect 46032 17672 46060 17700
rect 47026 17688 47032 17740
rect 47084 17728 47090 17740
rect 47397 17731 47455 17737
rect 47397 17728 47409 17731
rect 47084 17700 47409 17728
rect 47084 17688 47090 17700
rect 47397 17697 47409 17700
rect 47443 17728 47455 17731
rect 47443 17700 47900 17728
rect 47443 17697 47455 17700
rect 47397 17691 47455 17697
rect 47872 17672 47900 17700
rect 47946 17688 47952 17740
rect 48004 17728 48010 17740
rect 48004 17700 48360 17728
rect 48004 17688 48010 17700
rect 42705 17663 42763 17669
rect 42705 17629 42717 17663
rect 42751 17629 42763 17663
rect 42705 17623 42763 17629
rect 42981 17663 43039 17669
rect 42981 17629 42993 17663
rect 43027 17629 43039 17663
rect 42981 17623 43039 17629
rect 42996 17592 43024 17623
rect 43162 17620 43168 17672
rect 43220 17620 43226 17672
rect 43346 17620 43352 17672
rect 43404 17660 43410 17672
rect 43404 17620 43416 17660
rect 46014 17620 46020 17672
rect 46072 17620 46078 17672
rect 46106 17620 46112 17672
rect 46164 17620 46170 17672
rect 46385 17663 46443 17669
rect 46385 17629 46397 17663
rect 46431 17660 46443 17663
rect 46753 17663 46811 17669
rect 46753 17660 46765 17663
rect 46431 17632 46765 17660
rect 46431 17629 46443 17632
rect 46385 17623 46443 17629
rect 46753 17629 46765 17632
rect 46799 17629 46811 17663
rect 46753 17623 46811 17629
rect 47762 17620 47768 17672
rect 47820 17620 47826 17672
rect 47854 17620 47860 17672
rect 47912 17660 47918 17672
rect 47912 17632 47957 17660
rect 47912 17620 47918 17632
rect 48130 17620 48136 17672
rect 48188 17620 48194 17672
rect 48230 17663 48288 17669
rect 48230 17629 48242 17663
rect 48276 17660 48288 17663
rect 48332 17660 48360 17700
rect 49510 17688 49516 17740
rect 49568 17728 49574 17740
rect 50982 17728 50988 17740
rect 49568 17700 50988 17728
rect 49568 17688 49574 17700
rect 50982 17688 50988 17700
rect 51040 17688 51046 17740
rect 51353 17663 51411 17669
rect 51353 17660 51365 17663
rect 48276 17632 51365 17660
rect 48276 17629 48288 17632
rect 48230 17623 48288 17629
rect 51353 17629 51365 17632
rect 51399 17660 51411 17663
rect 51537 17663 51595 17669
rect 51537 17660 51549 17663
rect 51399 17632 51549 17660
rect 51399 17629 51411 17632
rect 51353 17623 51411 17629
rect 51537 17629 51549 17632
rect 51583 17629 51595 17663
rect 51644 17660 51672 17768
rect 52385 17768 53972 17796
rect 51902 17660 51908 17672
rect 51644 17632 51908 17660
rect 51537 17623 51595 17629
rect 51902 17620 51908 17632
rect 51960 17660 51966 17672
rect 52385 17660 52413 17768
rect 52454 17688 52460 17740
rect 52512 17728 52518 17740
rect 52512 17700 52868 17728
rect 52512 17688 52518 17700
rect 52840 17669 52868 17700
rect 52733 17663 52791 17669
rect 52733 17660 52745 17663
rect 51960 17632 52745 17660
rect 51960 17620 51966 17632
rect 52733 17629 52745 17632
rect 52779 17629 52791 17663
rect 52733 17623 52791 17629
rect 52826 17663 52884 17669
rect 52826 17629 52838 17663
rect 52872 17629 52884 17663
rect 53101 17663 53159 17669
rect 53101 17660 53113 17663
rect 52826 17623 52884 17629
rect 52932 17632 53113 17660
rect 43257 17595 43315 17601
rect 43257 17592 43269 17595
rect 41708 17564 43024 17592
rect 43180 17564 43269 17592
rect 43180 17536 43208 17564
rect 43257 17561 43269 17564
rect 43303 17561 43315 17595
rect 43388 17592 43416 17620
rect 43388 17564 45876 17592
rect 43257 17555 43315 17561
rect 39080 17496 39896 17524
rect 40497 17527 40555 17533
rect 39080 17484 39086 17496
rect 40497 17493 40509 17527
rect 40543 17524 40555 17527
rect 41322 17524 41328 17536
rect 40543 17496 41328 17524
rect 40543 17493 40555 17496
rect 40497 17487 40555 17493
rect 41322 17484 41328 17496
rect 41380 17484 41386 17536
rect 43162 17484 43168 17536
rect 43220 17484 43226 17536
rect 43438 17484 43444 17536
rect 43496 17524 43502 17536
rect 43533 17527 43591 17533
rect 43533 17524 43545 17527
rect 43496 17496 43545 17524
rect 43496 17484 43502 17496
rect 43533 17493 43545 17496
rect 43579 17493 43591 17527
rect 43533 17487 43591 17493
rect 43714 17484 43720 17536
rect 43772 17524 43778 17536
rect 44177 17527 44235 17533
rect 44177 17524 44189 17527
rect 43772 17496 44189 17524
rect 43772 17484 43778 17496
rect 44177 17493 44189 17496
rect 44223 17493 44235 17527
rect 45848 17524 45876 17564
rect 45922 17552 45928 17604
rect 45980 17592 45986 17604
rect 48041 17595 48099 17601
rect 48041 17592 48053 17595
rect 45980 17564 48053 17592
rect 45980 17552 45986 17564
rect 48041 17561 48053 17564
rect 48087 17592 48099 17595
rect 50338 17592 50344 17604
rect 48087 17564 50344 17592
rect 48087 17561 48099 17564
rect 48041 17555 48099 17561
rect 50338 17552 50344 17564
rect 50396 17552 50402 17604
rect 51074 17552 51080 17604
rect 51132 17592 51138 17604
rect 52932 17592 52960 17632
rect 53101 17629 53113 17632
rect 53147 17629 53159 17663
rect 53101 17623 53159 17629
rect 53190 17620 53196 17672
rect 53248 17669 53254 17672
rect 53944 17669 53972 17768
rect 54110 17756 54116 17808
rect 54168 17756 54174 17808
rect 54128 17728 54156 17756
rect 54037 17700 54156 17728
rect 54037 17669 54065 17700
rect 53248 17660 53256 17669
rect 53929 17663 53987 17669
rect 53248 17632 53293 17660
rect 53248 17623 53256 17632
rect 53929 17629 53941 17663
rect 53975 17629 53987 17663
rect 53929 17623 53987 17629
rect 54022 17663 54080 17669
rect 54022 17629 54034 17663
rect 54068 17629 54080 17663
rect 54022 17623 54080 17629
rect 53248 17620 53254 17623
rect 54110 17620 54116 17672
rect 54168 17660 54174 17672
rect 54394 17663 54452 17669
rect 54394 17660 54406 17663
rect 54168 17632 54406 17660
rect 54168 17620 54174 17632
rect 54394 17629 54406 17632
rect 54440 17660 54452 17663
rect 54570 17660 54576 17672
rect 54440 17632 54576 17660
rect 54440 17629 54452 17632
rect 54394 17623 54452 17629
rect 54570 17620 54576 17632
rect 54628 17620 54634 17672
rect 51132 17564 52960 17592
rect 51132 17552 51138 17564
rect 46198 17524 46204 17536
rect 45848 17496 46204 17524
rect 44177 17487 44235 17493
rect 46198 17484 46204 17496
rect 46256 17524 46262 17536
rect 47578 17524 47584 17536
rect 46256 17496 47584 17524
rect 46256 17484 46262 17496
rect 47578 17484 47584 17496
rect 47636 17484 47642 17536
rect 47762 17484 47768 17536
rect 47820 17524 47826 17536
rect 50246 17524 50252 17536
rect 47820 17496 50252 17524
rect 47820 17484 47826 17496
rect 50246 17484 50252 17496
rect 50304 17484 50310 17536
rect 52932 17524 52960 17564
rect 53006 17552 53012 17604
rect 53064 17592 53070 17604
rect 54205 17595 54263 17601
rect 54205 17592 54217 17595
rect 53064 17564 54217 17592
rect 53064 17552 53070 17564
rect 54128 17536 54156 17564
rect 54205 17561 54217 17564
rect 54251 17561 54263 17595
rect 54205 17555 54263 17561
rect 54297 17595 54355 17601
rect 54297 17561 54309 17595
rect 54343 17592 54355 17595
rect 55030 17592 55036 17604
rect 54343 17564 55036 17592
rect 54343 17561 54355 17564
rect 54297 17555 54355 17561
rect 55030 17552 55036 17564
rect 55088 17552 55094 17604
rect 53926 17524 53932 17536
rect 52932 17496 53932 17524
rect 53926 17484 53932 17496
rect 53984 17484 53990 17536
rect 54110 17484 54116 17536
rect 54168 17484 54174 17536
rect 1104 17434 78844 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 66314 17434
rect 66366 17382 66378 17434
rect 66430 17382 66442 17434
rect 66494 17382 66506 17434
rect 66558 17382 66570 17434
rect 66622 17382 78844 17434
rect 1104 17360 78844 17382
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 9548 17292 12204 17320
rect 9548 17280 9554 17292
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 9769 17255 9827 17261
rect 9769 17252 9781 17255
rect 9732 17224 9781 17252
rect 9732 17212 9738 17224
rect 9769 17221 9781 17224
rect 9815 17221 9827 17255
rect 9769 17215 9827 17221
rect 12176 17252 12204 17292
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 15105 17323 15163 17329
rect 15105 17320 15117 17323
rect 14792 17292 15117 17320
rect 14792 17280 14798 17292
rect 15105 17289 15117 17292
rect 15151 17289 15163 17323
rect 15105 17283 15163 17289
rect 15470 17280 15476 17332
rect 15528 17280 15534 17332
rect 15562 17280 15568 17332
rect 15620 17280 15626 17332
rect 20530 17320 20536 17332
rect 16132 17292 20536 17320
rect 12710 17252 12716 17264
rect 12176 17224 12716 17252
rect 9490 17144 9496 17196
rect 9548 17144 9554 17196
rect 11146 17184 11152 17196
rect 10902 17170 11152 17184
rect 10888 17156 11152 17170
rect 9306 17076 9312 17128
rect 9364 17116 9370 17128
rect 10778 17116 10784 17128
rect 9364 17088 10784 17116
rect 9364 17076 9370 17088
rect 10778 17076 10784 17088
rect 10836 17116 10842 17128
rect 10888 17116 10916 17156
rect 11146 17144 11152 17156
rect 11204 17144 11210 17196
rect 12176 17193 12204 17224
rect 12710 17212 12716 17224
rect 12768 17212 12774 17264
rect 13998 17252 14004 17264
rect 13662 17224 14004 17252
rect 13998 17212 14004 17224
rect 14056 17212 14062 17264
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 14182 17144 14188 17196
rect 14240 17184 14246 17196
rect 15488 17184 15516 17280
rect 16132 17193 16160 17292
rect 20530 17280 20536 17292
rect 20588 17280 20594 17332
rect 23661 17323 23719 17329
rect 23661 17289 23673 17323
rect 23707 17320 23719 17323
rect 29178 17320 29184 17332
rect 23707 17292 29184 17320
rect 23707 17289 23719 17292
rect 23661 17283 23719 17289
rect 29178 17280 29184 17292
rect 29236 17280 29242 17332
rect 29730 17280 29736 17332
rect 29788 17320 29794 17332
rect 30653 17323 30711 17329
rect 29788 17292 30604 17320
rect 29788 17280 29794 17292
rect 17954 17212 17960 17264
rect 18012 17212 18018 17264
rect 28350 17252 28356 17264
rect 28092 17224 28356 17252
rect 16117 17187 16175 17193
rect 16117 17184 16129 17187
rect 14240 17156 14780 17184
rect 15488 17156 16129 17184
rect 14240 17144 14246 17156
rect 10836 17088 10916 17116
rect 10836 17076 10842 17088
rect 11164 17048 11192 17144
rect 12434 17076 12440 17128
rect 12492 17076 12498 17128
rect 13909 17119 13967 17125
rect 13909 17085 13921 17119
rect 13955 17116 13967 17119
rect 14274 17116 14280 17128
rect 13955 17088 14280 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 14274 17076 14280 17088
rect 14332 17076 14338 17128
rect 14752 17048 14780 17156
rect 16117 17153 16129 17156
rect 16163 17153 16175 17187
rect 18877 17187 18935 17193
rect 18877 17184 18889 17187
rect 16117 17147 16175 17153
rect 18524 17156 18889 17184
rect 15010 17076 15016 17128
rect 15068 17116 15074 17128
rect 15657 17119 15715 17125
rect 15657 17116 15669 17119
rect 15068 17088 15669 17116
rect 15068 17076 15074 17088
rect 15657 17085 15669 17088
rect 15703 17085 15715 17119
rect 15657 17079 15715 17085
rect 16206 17076 16212 17128
rect 16264 17076 16270 17128
rect 16482 17076 16488 17128
rect 16540 17116 16546 17128
rect 17037 17119 17095 17125
rect 17037 17116 17049 17119
rect 16540 17088 17049 17116
rect 16540 17076 16546 17088
rect 17037 17085 17049 17088
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 17310 17076 17316 17128
rect 17368 17076 17374 17128
rect 18322 17076 18328 17128
rect 18380 17116 18386 17128
rect 18524 17116 18552 17156
rect 18877 17153 18889 17156
rect 18923 17153 18935 17187
rect 18877 17147 18935 17153
rect 23106 17144 23112 17196
rect 23164 17144 23170 17196
rect 23290 17144 23296 17196
rect 23348 17184 23354 17196
rect 23569 17187 23627 17193
rect 23569 17184 23581 17187
rect 23348 17156 23581 17184
rect 23348 17144 23354 17156
rect 23569 17153 23581 17156
rect 23615 17153 23627 17187
rect 23569 17147 23627 17153
rect 23753 17187 23811 17193
rect 23753 17153 23765 17187
rect 23799 17184 23811 17187
rect 24026 17184 24032 17196
rect 23799 17156 24032 17184
rect 23799 17153 23811 17156
rect 23753 17147 23811 17153
rect 24026 17144 24032 17156
rect 24084 17144 24090 17196
rect 27798 17144 27804 17196
rect 27856 17144 27862 17196
rect 28092 17193 28120 17224
rect 28350 17212 28356 17224
rect 28408 17212 28414 17264
rect 28810 17212 28816 17264
rect 28868 17252 28874 17264
rect 28868 17224 30144 17252
rect 28868 17212 28874 17224
rect 28077 17187 28135 17193
rect 28077 17153 28089 17187
rect 28123 17153 28135 17187
rect 28077 17147 28135 17153
rect 28258 17144 28264 17196
rect 28316 17184 28322 17196
rect 28316 17156 28396 17184
rect 28316 17144 28322 17156
rect 18380 17088 18552 17116
rect 18785 17119 18843 17125
rect 18380 17076 18386 17088
rect 18785 17085 18797 17119
rect 18831 17116 18843 17119
rect 18966 17116 18972 17128
rect 18831 17088 18972 17116
rect 18831 17085 18843 17088
rect 18785 17079 18843 17085
rect 18966 17076 18972 17088
rect 19024 17116 19030 17128
rect 19429 17119 19487 17125
rect 19429 17116 19441 17119
rect 19024 17088 19441 17116
rect 19024 17076 19030 17088
rect 19429 17085 19441 17088
rect 19475 17085 19487 17119
rect 20438 17116 20444 17128
rect 19429 17079 19487 17085
rect 20272 17088 20444 17116
rect 11164 17020 12296 17048
rect 14752 17020 17172 17048
rect 11241 16983 11299 16989
rect 11241 16949 11253 16983
rect 11287 16980 11299 16983
rect 12158 16980 12164 16992
rect 11287 16952 12164 16980
rect 11287 16949 11299 16952
rect 11241 16943 11299 16949
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 12268 16980 12296 17020
rect 13998 16980 14004 16992
rect 12268 16952 14004 16980
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 14458 16940 14464 16992
rect 14516 16940 14522 16992
rect 16393 16983 16451 16989
rect 16393 16949 16405 16983
rect 16439 16980 16451 16983
rect 17034 16980 17040 16992
rect 16439 16952 17040 16980
rect 16439 16949 16451 16952
rect 16393 16943 16451 16949
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 17144 16980 17172 17020
rect 19978 17008 19984 17060
rect 20036 17048 20042 17060
rect 20165 17051 20223 17057
rect 20165 17048 20177 17051
rect 20036 17020 20177 17048
rect 20036 17008 20042 17020
rect 20165 17017 20177 17020
rect 20211 17017 20223 17051
rect 20165 17011 20223 17017
rect 20070 16980 20076 16992
rect 17144 16952 20076 16980
rect 20070 16940 20076 16952
rect 20128 16980 20134 16992
rect 20272 16980 20300 17088
rect 20438 17076 20444 17088
rect 20496 17116 20502 17128
rect 20717 17119 20775 17125
rect 20717 17116 20729 17119
rect 20496 17088 20729 17116
rect 20496 17076 20502 17088
rect 20717 17085 20729 17088
rect 20763 17085 20775 17119
rect 20717 17079 20775 17085
rect 27430 17076 27436 17128
rect 27488 17116 27494 17128
rect 27709 17119 27767 17125
rect 27709 17116 27721 17119
rect 27488 17088 27721 17116
rect 27488 17076 27494 17088
rect 27709 17085 27721 17088
rect 27755 17085 27767 17119
rect 28368 17116 28396 17156
rect 28534 17144 28540 17196
rect 28592 17144 28598 17196
rect 28902 17144 28908 17196
rect 28960 17184 28966 17196
rect 29273 17187 29331 17193
rect 29273 17184 29285 17187
rect 28960 17156 29285 17184
rect 28960 17144 28966 17156
rect 29273 17153 29285 17156
rect 29319 17153 29331 17187
rect 29273 17147 29331 17153
rect 29362 17144 29368 17196
rect 29420 17184 29426 17196
rect 29457 17187 29515 17193
rect 29457 17184 29469 17187
rect 29420 17156 29469 17184
rect 29420 17144 29426 17156
rect 29457 17153 29469 17156
rect 29503 17184 29515 17187
rect 29822 17184 29828 17196
rect 29503 17156 29828 17184
rect 29503 17153 29515 17156
rect 29457 17147 29515 17153
rect 29822 17144 29828 17156
rect 29880 17144 29886 17196
rect 30006 17144 30012 17196
rect 30064 17144 30070 17196
rect 30116 17184 30144 17224
rect 30190 17212 30196 17264
rect 30248 17212 30254 17264
rect 30576 17252 30604 17292
rect 30653 17289 30665 17323
rect 30699 17320 30711 17323
rect 30742 17320 30748 17332
rect 30699 17292 30748 17320
rect 30699 17289 30711 17292
rect 30653 17283 30711 17289
rect 30742 17280 30748 17292
rect 30800 17280 30806 17332
rect 31018 17280 31024 17332
rect 31076 17280 31082 17332
rect 31481 17323 31539 17329
rect 31481 17289 31493 17323
rect 31527 17320 31539 17323
rect 32030 17320 32036 17332
rect 31527 17292 32036 17320
rect 31527 17289 31539 17292
rect 31481 17283 31539 17289
rect 32030 17280 32036 17292
rect 32088 17280 32094 17332
rect 32217 17323 32275 17329
rect 32217 17289 32229 17323
rect 32263 17320 32275 17323
rect 33134 17320 33140 17332
rect 32263 17292 33140 17320
rect 32263 17289 32275 17292
rect 32217 17283 32275 17289
rect 30576 17224 30788 17252
rect 30285 17187 30343 17193
rect 30285 17184 30297 17187
rect 30116 17156 30297 17184
rect 30285 17153 30297 17156
rect 30331 17153 30343 17187
rect 30285 17147 30343 17153
rect 30469 17187 30527 17193
rect 30469 17153 30481 17187
rect 30515 17184 30527 17187
rect 30650 17184 30656 17196
rect 30515 17156 30656 17184
rect 30515 17153 30527 17156
rect 30469 17147 30527 17153
rect 30650 17144 30656 17156
rect 30708 17144 30714 17196
rect 30760 17193 30788 17224
rect 30745 17187 30803 17193
rect 30745 17153 30757 17187
rect 30791 17153 30803 17187
rect 30745 17147 30803 17153
rect 31297 17187 31355 17193
rect 31297 17153 31309 17187
rect 31343 17153 31355 17187
rect 31297 17147 31355 17153
rect 31941 17187 31999 17193
rect 31941 17153 31953 17187
rect 31987 17184 31999 17187
rect 32232 17184 32260 17283
rect 33134 17280 33140 17292
rect 33192 17320 33198 17332
rect 33192 17292 41414 17320
rect 33192 17280 33198 17292
rect 32677 17255 32735 17261
rect 32677 17221 32689 17255
rect 32723 17252 32735 17255
rect 32723 17224 34836 17252
rect 32723 17221 32735 17224
rect 32677 17215 32735 17221
rect 34808 17196 34836 17224
rect 36446 17212 36452 17264
rect 36504 17252 36510 17264
rect 38746 17252 38752 17264
rect 36504 17224 36768 17252
rect 36504 17212 36510 17224
rect 31987 17156 32260 17184
rect 31987 17153 31999 17156
rect 31941 17147 31999 17153
rect 29178 17116 29184 17128
rect 28368 17088 29184 17116
rect 27709 17079 27767 17085
rect 29178 17076 29184 17088
rect 29236 17076 29242 17128
rect 29730 17076 29736 17128
rect 29788 17076 29794 17128
rect 30024 17116 30052 17144
rect 31018 17116 31024 17128
rect 30024 17088 31024 17116
rect 31018 17076 31024 17088
rect 31076 17076 31082 17128
rect 20530 17008 20536 17060
rect 20588 17008 20594 17060
rect 23385 17051 23443 17057
rect 23385 17017 23397 17051
rect 23431 17017 23443 17051
rect 23385 17011 23443 17017
rect 20128 16952 20300 16980
rect 20128 16940 20134 16952
rect 20438 16940 20444 16992
rect 20496 16980 20502 16992
rect 20548 16980 20576 17008
rect 20496 16952 20576 16980
rect 20496 16940 20502 16952
rect 20622 16940 20628 16992
rect 20680 16940 20686 16992
rect 20806 16940 20812 16992
rect 20864 16940 20870 16992
rect 23400 16980 23428 17011
rect 28166 17008 28172 17060
rect 28224 17048 28230 17060
rect 28810 17048 28816 17060
rect 28224 17020 28816 17048
rect 28224 17008 28230 17020
rect 28810 17008 28816 17020
rect 28868 17008 28874 17060
rect 29086 17048 29092 17060
rect 28966 17020 29092 17048
rect 27706 16980 27712 16992
rect 23400 16952 27712 16980
rect 27706 16940 27712 16952
rect 27764 16980 27770 16992
rect 28626 16980 28632 16992
rect 27764 16952 28632 16980
rect 27764 16940 27770 16952
rect 28626 16940 28632 16952
rect 28684 16980 28690 16992
rect 28966 16980 28994 17020
rect 29086 17008 29092 17020
rect 29144 17008 29150 17060
rect 28684 16952 28994 16980
rect 28684 16940 28690 16952
rect 29178 16940 29184 16992
rect 29236 16980 29242 16992
rect 29641 16983 29699 16989
rect 29641 16980 29653 16983
rect 29236 16952 29653 16980
rect 29236 16940 29242 16952
rect 29641 16949 29653 16952
rect 29687 16980 29699 16983
rect 29825 16983 29883 16989
rect 29825 16980 29837 16983
rect 29687 16952 29837 16980
rect 29687 16949 29699 16952
rect 29641 16943 29699 16949
rect 29825 16949 29837 16952
rect 29871 16980 29883 16983
rect 30837 16983 30895 16989
rect 30837 16980 30849 16983
rect 29871 16952 30849 16980
rect 29871 16949 29883 16952
rect 29825 16943 29883 16949
rect 30837 16949 30849 16952
rect 30883 16949 30895 16983
rect 30837 16943 30895 16949
rect 31205 16983 31263 16989
rect 31205 16949 31217 16983
rect 31251 16980 31263 16983
rect 31312 16980 31340 17147
rect 32582 17144 32588 17196
rect 32640 17144 32646 17196
rect 32769 17187 32827 17193
rect 32769 17153 32781 17187
rect 32815 17184 32827 17187
rect 32858 17184 32864 17196
rect 32815 17156 32864 17184
rect 32815 17153 32827 17156
rect 32769 17147 32827 17153
rect 32858 17144 32864 17156
rect 32916 17144 32922 17196
rect 32950 17144 32956 17196
rect 33008 17144 33014 17196
rect 33137 17187 33195 17193
rect 33137 17153 33149 17187
rect 33183 17184 33195 17187
rect 33226 17184 33232 17196
rect 33183 17156 33232 17184
rect 33183 17153 33195 17156
rect 33137 17147 33195 17153
rect 33226 17144 33232 17156
rect 33284 17184 33290 17196
rect 33284 17156 33364 17184
rect 33284 17144 33290 17156
rect 33336 17048 33364 17156
rect 33594 17144 33600 17196
rect 33652 17144 33658 17196
rect 34054 17144 34060 17196
rect 34112 17184 34118 17196
rect 34425 17187 34483 17193
rect 34425 17184 34437 17187
rect 34112 17156 34437 17184
rect 34112 17144 34118 17156
rect 34425 17153 34437 17156
rect 34471 17153 34483 17187
rect 34425 17147 34483 17153
rect 34514 17144 34520 17196
rect 34572 17144 34578 17196
rect 34790 17144 34796 17196
rect 34848 17144 34854 17196
rect 36740 17193 36768 17224
rect 38028 17224 38752 17252
rect 36633 17187 36691 17193
rect 36633 17153 36645 17187
rect 36679 17153 36691 17187
rect 36633 17147 36691 17153
rect 36725 17187 36783 17193
rect 36725 17153 36737 17187
rect 36771 17153 36783 17187
rect 36725 17147 36783 17153
rect 33410 17076 33416 17128
rect 33468 17116 33474 17128
rect 34330 17116 34336 17128
rect 33468 17088 34336 17116
rect 33468 17076 33474 17088
rect 34330 17076 34336 17088
rect 34388 17116 34394 17128
rect 34701 17119 34759 17125
rect 34701 17116 34713 17119
rect 34388 17088 34713 17116
rect 34388 17076 34394 17088
rect 34701 17085 34713 17088
rect 34747 17085 34759 17119
rect 34701 17079 34759 17085
rect 33336 17020 33824 17048
rect 31754 16980 31760 16992
rect 31251 16952 31760 16980
rect 31251 16949 31263 16952
rect 31205 16943 31263 16949
rect 31754 16940 31760 16952
rect 31812 16940 31818 16992
rect 32398 16940 32404 16992
rect 32456 16940 32462 16992
rect 33796 16989 33824 17020
rect 34054 17008 34060 17060
rect 34112 17048 34118 17060
rect 36648 17048 36676 17147
rect 36998 17144 37004 17196
rect 37056 17144 37062 17196
rect 38028 17193 38056 17224
rect 38746 17212 38752 17224
rect 38804 17212 38810 17264
rect 41230 17252 41236 17264
rect 40066 17224 41236 17252
rect 41230 17212 41236 17224
rect 41288 17212 41294 17264
rect 41386 17252 41414 17292
rect 43070 17280 43076 17332
rect 43128 17320 43134 17332
rect 43165 17323 43223 17329
rect 43165 17320 43177 17323
rect 43128 17292 43177 17320
rect 43128 17280 43134 17292
rect 43165 17289 43177 17292
rect 43211 17289 43223 17323
rect 45646 17320 45652 17332
rect 43165 17283 43223 17289
rect 43272 17292 45652 17320
rect 42521 17255 42579 17261
rect 42521 17252 42533 17255
rect 41386 17224 42533 17252
rect 42521 17221 42533 17224
rect 42567 17252 42579 17255
rect 42702 17252 42708 17264
rect 42567 17224 42708 17252
rect 42567 17221 42579 17224
rect 42521 17215 42579 17221
rect 42702 17212 42708 17224
rect 42760 17252 42766 17264
rect 43272 17252 43300 17292
rect 45646 17280 45652 17292
rect 45704 17280 45710 17332
rect 46106 17280 46112 17332
rect 46164 17320 46170 17332
rect 46293 17323 46351 17329
rect 46293 17320 46305 17323
rect 46164 17292 46305 17320
rect 46164 17280 46170 17292
rect 46293 17289 46305 17292
rect 46339 17289 46351 17323
rect 46293 17283 46351 17289
rect 50065 17323 50123 17329
rect 50065 17289 50077 17323
rect 50111 17320 50123 17323
rect 50522 17320 50528 17332
rect 50111 17292 50528 17320
rect 50111 17289 50123 17292
rect 50065 17283 50123 17289
rect 50522 17280 50528 17292
rect 50580 17320 50586 17332
rect 50706 17320 50712 17332
rect 50580 17292 50712 17320
rect 50580 17280 50586 17292
rect 50706 17280 50712 17292
rect 50764 17280 50770 17332
rect 52362 17280 52368 17332
rect 52420 17320 52426 17332
rect 53006 17320 53012 17332
rect 52420 17292 53012 17320
rect 52420 17280 52426 17292
rect 53006 17280 53012 17292
rect 53064 17280 53070 17332
rect 44913 17255 44971 17261
rect 44913 17252 44925 17255
rect 42760 17224 43300 17252
rect 43364 17224 44925 17252
rect 42760 17212 42766 17224
rect 38013 17187 38071 17193
rect 38013 17153 38025 17187
rect 38059 17153 38071 17187
rect 38013 17147 38071 17153
rect 38289 17187 38347 17193
rect 38289 17153 38301 17187
rect 38335 17184 38347 17187
rect 38378 17184 38384 17196
rect 38335 17156 38384 17184
rect 38335 17153 38347 17156
rect 38289 17147 38347 17153
rect 38378 17144 38384 17156
rect 38436 17144 38442 17196
rect 38562 17144 38568 17196
rect 38620 17144 38626 17196
rect 41046 17184 41052 17196
rect 40052 17156 41052 17184
rect 38473 17119 38531 17125
rect 38473 17085 38485 17119
rect 38519 17116 38531 17119
rect 38841 17119 38899 17125
rect 38841 17116 38853 17119
rect 38519 17088 38853 17116
rect 38519 17085 38531 17088
rect 38473 17079 38531 17085
rect 38841 17085 38853 17088
rect 38887 17085 38899 17119
rect 38841 17079 38899 17085
rect 38930 17076 38936 17128
rect 38988 17116 38994 17128
rect 40052 17116 40080 17156
rect 41046 17144 41052 17156
rect 41104 17144 41110 17196
rect 41322 17144 41328 17196
rect 41380 17144 41386 17196
rect 41414 17144 41420 17196
rect 41472 17184 41478 17196
rect 41690 17184 41696 17196
rect 41472 17156 41696 17184
rect 41472 17144 41478 17156
rect 41690 17144 41696 17156
rect 41748 17144 41754 17196
rect 42978 17144 42984 17196
rect 43036 17184 43042 17196
rect 43364 17193 43392 17224
rect 44913 17221 44925 17224
rect 44959 17252 44971 17255
rect 44959 17224 45876 17252
rect 44959 17221 44971 17224
rect 44913 17215 44971 17221
rect 43073 17187 43131 17193
rect 43073 17184 43085 17187
rect 43036 17156 43085 17184
rect 43036 17144 43042 17156
rect 43073 17153 43085 17156
rect 43119 17184 43131 17187
rect 43349 17187 43407 17193
rect 43349 17184 43361 17187
rect 43119 17156 43361 17184
rect 43119 17153 43131 17156
rect 43073 17147 43131 17153
rect 43349 17153 43361 17156
rect 43395 17153 43407 17187
rect 43349 17147 43407 17153
rect 43438 17144 43444 17196
rect 43496 17144 43502 17196
rect 43714 17144 43720 17196
rect 43772 17144 43778 17196
rect 45204 17193 45232 17224
rect 45189 17187 45247 17193
rect 45189 17153 45201 17187
rect 45235 17153 45247 17187
rect 45189 17147 45247 17153
rect 45281 17187 45339 17193
rect 45281 17153 45293 17187
rect 45327 17184 45339 17187
rect 45462 17184 45468 17196
rect 45327 17156 45468 17184
rect 45327 17153 45339 17156
rect 45281 17147 45339 17153
rect 45462 17144 45468 17156
rect 45520 17144 45526 17196
rect 45554 17144 45560 17196
rect 45612 17144 45618 17196
rect 45738 17144 45744 17196
rect 45796 17144 45802 17196
rect 45848 17184 45876 17224
rect 45922 17212 45928 17264
rect 45980 17212 45986 17264
rect 46017 17255 46075 17261
rect 46017 17221 46029 17255
rect 46063 17252 46075 17255
rect 50614 17252 50620 17264
rect 46063 17224 50620 17252
rect 46063 17221 46075 17224
rect 46017 17215 46075 17221
rect 50614 17212 50620 17224
rect 50672 17212 50678 17264
rect 54110 17212 54116 17264
rect 54168 17252 54174 17264
rect 54478 17252 54484 17264
rect 54168 17224 54484 17252
rect 54168 17212 54174 17224
rect 54478 17212 54484 17224
rect 54536 17212 54542 17264
rect 46109 17187 46167 17193
rect 45848 17156 46060 17184
rect 46032 17128 46060 17156
rect 46109 17153 46121 17187
rect 46155 17184 46167 17187
rect 46198 17184 46204 17196
rect 46155 17156 46204 17184
rect 46155 17153 46167 17156
rect 46109 17147 46167 17153
rect 46198 17144 46204 17156
rect 46256 17184 46262 17196
rect 46385 17187 46443 17193
rect 46385 17184 46397 17187
rect 46256 17156 46397 17184
rect 46256 17144 46262 17156
rect 46385 17153 46397 17156
rect 46431 17153 46443 17187
rect 46385 17147 46443 17153
rect 48038 17144 48044 17196
rect 48096 17184 48102 17196
rect 48317 17187 48375 17193
rect 48317 17184 48329 17187
rect 48096 17156 48329 17184
rect 48096 17144 48102 17156
rect 48317 17153 48329 17156
rect 48363 17184 48375 17187
rect 49050 17184 49056 17196
rect 48363 17156 49056 17184
rect 48363 17153 48375 17156
rect 48317 17147 48375 17153
rect 49050 17144 49056 17156
rect 49108 17144 49114 17196
rect 50338 17144 50344 17196
rect 50396 17184 50402 17196
rect 52181 17187 52239 17193
rect 52181 17184 52193 17187
rect 50396 17156 52193 17184
rect 50396 17144 50402 17156
rect 52181 17153 52193 17156
rect 52227 17153 52239 17187
rect 52181 17147 52239 17153
rect 53837 17187 53895 17193
rect 53837 17153 53849 17187
rect 53883 17153 53895 17187
rect 53837 17147 53895 17153
rect 38988 17088 40080 17116
rect 38988 17076 38994 17088
rect 40218 17076 40224 17128
rect 40276 17116 40282 17128
rect 40313 17119 40371 17125
rect 40313 17116 40325 17119
rect 40276 17088 40325 17116
rect 40276 17076 40282 17088
rect 40313 17085 40325 17088
rect 40359 17085 40371 17119
rect 40313 17079 40371 17085
rect 41141 17119 41199 17125
rect 41141 17085 41153 17119
rect 41187 17116 41199 17119
rect 42426 17116 42432 17128
rect 41187 17088 42432 17116
rect 41187 17085 41199 17088
rect 41141 17079 41199 17085
rect 34112 17020 36676 17048
rect 34112 17008 34118 17020
rect 33781 16983 33839 16989
rect 33781 16949 33793 16983
rect 33827 16980 33839 16983
rect 33965 16983 34023 16989
rect 33965 16980 33977 16983
rect 33827 16952 33977 16980
rect 33827 16949 33839 16952
rect 33781 16943 33839 16949
rect 33965 16949 33977 16952
rect 34011 16980 34023 16983
rect 34146 16980 34152 16992
rect 34011 16952 34152 16980
rect 34011 16949 34023 16952
rect 33965 16943 34023 16949
rect 34146 16940 34152 16952
rect 34204 16940 34210 16992
rect 34238 16940 34244 16992
rect 34296 16940 34302 16992
rect 36446 16940 36452 16992
rect 36504 16940 36510 16992
rect 36909 16983 36967 16989
rect 36909 16949 36921 16983
rect 36955 16980 36967 16983
rect 37274 16980 37280 16992
rect 36955 16952 37280 16980
rect 36955 16949 36967 16952
rect 36909 16943 36967 16949
rect 37274 16940 37280 16952
rect 37332 16980 37338 16992
rect 38105 16983 38163 16989
rect 38105 16980 38117 16983
rect 37332 16952 38117 16980
rect 37332 16940 37338 16952
rect 38105 16949 38117 16952
rect 38151 16980 38163 16983
rect 39942 16980 39948 16992
rect 38151 16952 39948 16980
rect 38151 16949 38163 16952
rect 38105 16943 38163 16949
rect 39942 16940 39948 16952
rect 40000 16980 40006 16992
rect 41156 16980 41184 17079
rect 42426 17076 42432 17088
rect 42484 17076 42490 17128
rect 45002 17076 45008 17128
rect 45060 17076 45066 17128
rect 46014 17076 46020 17128
rect 46072 17076 46078 17128
rect 49694 17076 49700 17128
rect 49752 17116 49758 17128
rect 50525 17119 50583 17125
rect 50525 17116 50537 17119
rect 49752 17088 50537 17116
rect 49752 17076 49758 17088
rect 41414 17008 41420 17060
rect 41472 17048 41478 17060
rect 41472 17020 41644 17048
rect 41472 17008 41478 17020
rect 40000 16952 41184 16980
rect 40000 16940 40006 16952
rect 41322 16940 41328 16992
rect 41380 16980 41386 16992
rect 41509 16983 41567 16989
rect 41509 16980 41521 16983
rect 41380 16952 41521 16980
rect 41380 16940 41386 16952
rect 41509 16949 41521 16952
rect 41555 16949 41567 16983
rect 41616 16980 41644 17020
rect 41690 17008 41696 17060
rect 41748 17048 41754 17060
rect 45830 17048 45836 17060
rect 41748 17020 45836 17048
rect 41748 17008 41754 17020
rect 45830 17008 45836 17020
rect 45888 17008 45894 17060
rect 49881 17051 49939 17057
rect 49881 17017 49893 17051
rect 49927 17048 49939 17051
rect 50062 17048 50068 17060
rect 49927 17020 50068 17048
rect 49927 17017 49939 17020
rect 49881 17011 49939 17017
rect 50062 17008 50068 17020
rect 50120 17008 50126 17060
rect 42245 16983 42303 16989
rect 42245 16980 42257 16983
rect 41616 16952 42257 16980
rect 41509 16943 41567 16949
rect 42245 16949 42257 16952
rect 42291 16980 42303 16983
rect 42334 16980 42340 16992
rect 42291 16952 42340 16980
rect 42291 16949 42303 16952
rect 42245 16943 42303 16949
rect 42334 16940 42340 16952
rect 42392 16940 42398 16992
rect 43622 16940 43628 16992
rect 43680 16980 43686 16992
rect 45465 16983 45523 16989
rect 45465 16980 45477 16983
rect 43680 16952 45477 16980
rect 43680 16940 43686 16952
rect 45465 16949 45477 16952
rect 45511 16980 45523 16983
rect 46290 16980 46296 16992
rect 45511 16952 46296 16980
rect 45511 16949 45523 16952
rect 45465 16943 45523 16949
rect 46290 16940 46296 16952
rect 46348 16940 46354 16992
rect 48593 16983 48651 16989
rect 48593 16949 48605 16983
rect 48639 16980 48651 16983
rect 48866 16980 48872 16992
rect 48639 16952 48872 16980
rect 48639 16949 48651 16952
rect 48593 16943 48651 16949
rect 48866 16940 48872 16952
rect 48924 16940 48930 16992
rect 50172 16980 50200 17088
rect 50525 17085 50537 17088
rect 50571 17085 50583 17119
rect 50525 17079 50583 17085
rect 51258 16980 51264 16992
rect 50172 16952 51264 16980
rect 51258 16940 51264 16952
rect 51316 16940 51322 16992
rect 53745 16983 53803 16989
rect 53745 16949 53757 16983
rect 53791 16980 53803 16983
rect 53852 16980 53880 17147
rect 53926 17144 53932 17196
rect 53984 17184 53990 17196
rect 53984 17156 54029 17184
rect 53984 17144 53990 17156
rect 54202 17144 54208 17196
rect 54260 17144 54266 17196
rect 54343 17187 54401 17193
rect 54343 17153 54355 17187
rect 54389 17184 54401 17187
rect 54570 17184 54576 17196
rect 54389 17156 54576 17184
rect 54389 17153 54401 17156
rect 54343 17147 54401 17153
rect 54570 17144 54576 17156
rect 54628 17144 54634 17196
rect 77846 17144 77852 17196
rect 77904 17184 77910 17196
rect 78033 17187 78091 17193
rect 78033 17184 78045 17187
rect 77904 17156 78045 17184
rect 77904 17144 77910 17156
rect 78033 17153 78045 17156
rect 78079 17153 78091 17187
rect 78033 17147 78091 17153
rect 78214 17008 78220 17060
rect 78272 17008 78278 17060
rect 54110 16980 54116 16992
rect 53791 16952 54116 16980
rect 53791 16949 53803 16952
rect 53745 16943 53803 16949
rect 54110 16940 54116 16952
rect 54168 16940 54174 16992
rect 54481 16983 54539 16989
rect 54481 16949 54493 16983
rect 54527 16980 54539 16983
rect 54754 16980 54760 16992
rect 54527 16952 54760 16980
rect 54527 16949 54539 16952
rect 54481 16943 54539 16949
rect 54754 16940 54760 16952
rect 54812 16940 54818 16992
rect 77846 16940 77852 16992
rect 77904 16940 77910 16992
rect 1104 16890 78844 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 78844 16890
rect 1104 16816 78844 16838
rect 12805 16779 12863 16785
rect 12805 16745 12817 16779
rect 12851 16776 12863 16779
rect 14090 16776 14096 16788
rect 12851 16748 14096 16776
rect 12851 16745 12863 16748
rect 12805 16739 12863 16745
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 20438 16736 20444 16788
rect 20496 16736 20502 16788
rect 20622 16776 20628 16788
rect 20548 16748 20628 16776
rect 11701 16711 11759 16717
rect 11701 16708 11713 16711
rect 11624 16680 11713 16708
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16572 10655 16575
rect 11624 16572 11652 16680
rect 11701 16677 11713 16680
rect 11747 16708 11759 16711
rect 17494 16708 17500 16720
rect 11747 16680 17500 16708
rect 11747 16677 11759 16680
rect 11701 16671 11759 16677
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 20548 16717 20576 16748
rect 20622 16736 20628 16748
rect 20680 16736 20686 16788
rect 20990 16736 20996 16788
rect 21048 16776 21054 16788
rect 25409 16779 25467 16785
rect 21048 16748 23980 16776
rect 21048 16736 21054 16748
rect 20533 16711 20591 16717
rect 20533 16708 20545 16711
rect 17604 16680 20545 16708
rect 12618 16600 12624 16652
rect 12676 16600 12682 16652
rect 10643 16544 11652 16572
rect 10643 16541 10655 16544
rect 10597 16535 10655 16541
rect 12158 16532 12164 16584
rect 12216 16572 12222 16584
rect 12529 16575 12587 16581
rect 12529 16572 12541 16575
rect 12216 16544 12541 16572
rect 12216 16532 12222 16544
rect 12529 16541 12541 16544
rect 12575 16572 12587 16575
rect 17604 16572 17632 16680
rect 20533 16677 20545 16680
rect 20579 16677 20591 16711
rect 20533 16671 20591 16677
rect 22925 16711 22983 16717
rect 22925 16677 22937 16711
rect 22971 16708 22983 16711
rect 23474 16708 23480 16720
rect 22971 16680 23480 16708
rect 22971 16677 22983 16680
rect 22925 16671 22983 16677
rect 23474 16668 23480 16680
rect 23532 16708 23538 16720
rect 23532 16680 23888 16708
rect 23532 16668 23538 16680
rect 18325 16643 18383 16649
rect 18325 16609 18337 16643
rect 18371 16640 18383 16643
rect 18414 16640 18420 16652
rect 18371 16612 18420 16640
rect 18371 16609 18383 16612
rect 18325 16603 18383 16609
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 18966 16600 18972 16652
rect 19024 16600 19030 16652
rect 20625 16643 20683 16649
rect 20625 16640 20637 16643
rect 19996 16612 20637 16640
rect 19996 16584 20024 16612
rect 20625 16609 20637 16612
rect 20671 16609 20683 16643
rect 20625 16603 20683 16609
rect 22094 16600 22100 16652
rect 22152 16640 22158 16652
rect 23106 16640 23112 16652
rect 22152 16612 23112 16640
rect 22152 16600 22158 16612
rect 12575 16544 17632 16572
rect 12575 16541 12587 16544
rect 12529 16535 12587 16541
rect 18046 16532 18052 16584
rect 18104 16572 18110 16584
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 18104 16544 18889 16572
rect 18104 16532 18110 16544
rect 18877 16541 18889 16544
rect 18923 16572 18935 16575
rect 19978 16572 19984 16584
rect 18923 16544 19984 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19978 16532 19984 16544
rect 20036 16532 20042 16584
rect 20070 16532 20076 16584
rect 20128 16532 20134 16584
rect 21450 16532 21456 16584
rect 21508 16572 21514 16584
rect 23032 16581 23060 16612
rect 23106 16600 23112 16612
rect 23164 16640 23170 16652
rect 23164 16612 23336 16640
rect 23164 16600 23170 16612
rect 22741 16575 22799 16581
rect 22741 16572 22753 16575
rect 21508 16544 22753 16572
rect 21508 16532 21514 16544
rect 22741 16541 22753 16544
rect 22787 16541 22799 16575
rect 22741 16535 22799 16541
rect 22925 16575 22983 16581
rect 22925 16541 22937 16575
rect 22971 16541 22983 16575
rect 22925 16535 22983 16541
rect 23017 16575 23075 16581
rect 23017 16541 23029 16575
rect 23063 16541 23075 16575
rect 23198 16572 23204 16584
rect 23017 16535 23075 16541
rect 23124 16544 23204 16572
rect 11425 16507 11483 16513
rect 11425 16473 11437 16507
rect 11471 16504 11483 16507
rect 11514 16504 11520 16516
rect 11471 16476 11520 16504
rect 11471 16473 11483 16476
rect 11425 16467 11483 16473
rect 11514 16464 11520 16476
rect 11572 16504 11578 16516
rect 12710 16504 12716 16516
rect 11572 16476 12716 16504
rect 11572 16464 11578 16476
rect 12710 16464 12716 16476
rect 12768 16504 12774 16516
rect 13630 16504 13636 16516
rect 12768 16476 13636 16504
rect 12768 16464 12774 16476
rect 13630 16464 13636 16476
rect 13688 16464 13694 16516
rect 18141 16507 18199 16513
rect 18141 16473 18153 16507
rect 18187 16504 18199 16507
rect 18322 16504 18328 16516
rect 18187 16476 18328 16504
rect 18187 16473 18199 16476
rect 18141 16467 18199 16473
rect 18322 16464 18328 16476
rect 18380 16464 18386 16516
rect 20806 16464 20812 16516
rect 20864 16504 20870 16516
rect 22940 16504 22968 16535
rect 23124 16504 23152 16544
rect 23198 16532 23204 16544
rect 23256 16532 23262 16584
rect 23308 16572 23336 16612
rect 23477 16575 23535 16581
rect 23477 16572 23489 16575
rect 23308 16544 23489 16572
rect 23477 16541 23489 16544
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16541 23719 16575
rect 23661 16535 23719 16541
rect 23676 16504 23704 16535
rect 20864 16476 23152 16504
rect 23216 16476 23704 16504
rect 23860 16504 23888 16680
rect 23952 16581 23980 16748
rect 25409 16745 25421 16779
rect 25455 16776 25467 16779
rect 25498 16776 25504 16788
rect 25455 16748 25504 16776
rect 25455 16745 25467 16748
rect 25409 16739 25467 16745
rect 25498 16736 25504 16748
rect 25556 16736 25562 16788
rect 25685 16779 25743 16785
rect 25685 16745 25697 16779
rect 25731 16776 25743 16779
rect 28166 16776 28172 16788
rect 25731 16748 28172 16776
rect 25731 16745 25743 16748
rect 25685 16739 25743 16745
rect 28166 16736 28172 16748
rect 28224 16736 28230 16788
rect 28258 16736 28264 16788
rect 28316 16736 28322 16788
rect 28534 16736 28540 16788
rect 28592 16776 28598 16788
rect 29730 16776 29736 16788
rect 28592 16748 29736 16776
rect 28592 16736 28598 16748
rect 29730 16736 29736 16748
rect 29788 16736 29794 16788
rect 32582 16776 32588 16788
rect 31680 16748 32588 16776
rect 25777 16711 25835 16717
rect 25777 16677 25789 16711
rect 25823 16708 25835 16711
rect 26237 16711 26295 16717
rect 26237 16708 26249 16711
rect 25823 16680 26249 16708
rect 25823 16677 25835 16680
rect 25777 16671 25835 16677
rect 26237 16677 26249 16680
rect 26283 16677 26295 16711
rect 26237 16671 26295 16677
rect 27801 16711 27859 16717
rect 27801 16677 27813 16711
rect 27847 16708 27859 16711
rect 28350 16708 28356 16720
rect 27847 16680 28356 16708
rect 27847 16677 27859 16680
rect 27801 16671 27859 16677
rect 24762 16600 24768 16652
rect 24820 16640 24826 16652
rect 28276 16649 28304 16680
rect 28350 16668 28356 16680
rect 28408 16668 28414 16720
rect 28902 16668 28908 16720
rect 28960 16708 28966 16720
rect 31680 16708 31708 16748
rect 32582 16736 32588 16748
rect 32640 16736 32646 16788
rect 36538 16736 36544 16788
rect 36596 16776 36602 16788
rect 38013 16779 38071 16785
rect 38013 16776 38025 16779
rect 36596 16748 38025 16776
rect 36596 16736 36602 16748
rect 38013 16745 38025 16748
rect 38059 16776 38071 16779
rect 38194 16776 38200 16788
rect 38059 16748 38200 16776
rect 38059 16745 38071 16748
rect 38013 16739 38071 16745
rect 38194 16736 38200 16748
rect 38252 16736 38258 16788
rect 38378 16736 38384 16788
rect 38436 16736 38442 16788
rect 41046 16736 41052 16788
rect 41104 16776 41110 16788
rect 42797 16779 42855 16785
rect 42797 16776 42809 16779
rect 41104 16748 42809 16776
rect 41104 16736 41110 16748
rect 42797 16745 42809 16748
rect 42843 16776 42855 16779
rect 43162 16776 43168 16788
rect 42843 16748 43168 16776
rect 42843 16745 42855 16748
rect 42797 16739 42855 16745
rect 43162 16736 43168 16748
rect 43220 16736 43226 16788
rect 45554 16736 45560 16788
rect 45612 16776 45618 16788
rect 45833 16779 45891 16785
rect 45833 16776 45845 16779
rect 45612 16748 45845 16776
rect 45612 16736 45618 16748
rect 45833 16745 45845 16748
rect 45879 16745 45891 16779
rect 45833 16739 45891 16745
rect 46014 16736 46020 16788
rect 46072 16736 46078 16788
rect 46290 16736 46296 16788
rect 46348 16736 46354 16788
rect 47670 16736 47676 16788
rect 47728 16776 47734 16788
rect 47728 16748 48176 16776
rect 47728 16736 47734 16748
rect 28960 16680 31708 16708
rect 28960 16668 28966 16680
rect 37550 16668 37556 16720
rect 37608 16668 37614 16720
rect 38470 16668 38476 16720
rect 38528 16668 38534 16720
rect 44821 16711 44879 16717
rect 44821 16677 44833 16711
rect 44867 16708 44879 16711
rect 44867 16680 45324 16708
rect 44867 16677 44879 16680
rect 44821 16671 44879 16677
rect 25869 16643 25927 16649
rect 25869 16640 25881 16643
rect 24820 16612 25881 16640
rect 24820 16600 24826 16612
rect 25869 16609 25881 16612
rect 25915 16609 25927 16643
rect 28261 16643 28319 16649
rect 25869 16603 25927 16609
rect 26344 16612 28120 16640
rect 23937 16575 23995 16581
rect 23937 16541 23949 16575
rect 23983 16541 23995 16575
rect 23937 16535 23995 16541
rect 24026 16532 24032 16584
rect 24084 16572 24090 16584
rect 24121 16575 24179 16581
rect 24121 16572 24133 16575
rect 24084 16544 24133 16572
rect 24084 16532 24090 16544
rect 24121 16541 24133 16544
rect 24167 16541 24179 16575
rect 24121 16535 24179 16541
rect 26145 16575 26203 16581
rect 26145 16541 26157 16575
rect 26191 16572 26203 16575
rect 26234 16572 26240 16584
rect 26191 16544 26240 16572
rect 26191 16541 26203 16544
rect 26145 16535 26203 16541
rect 26234 16532 26240 16544
rect 26292 16532 26298 16584
rect 26344 16572 26372 16612
rect 26421 16575 26479 16581
rect 26421 16572 26433 16575
rect 26344 16544 26433 16572
rect 26421 16541 26433 16544
rect 26467 16541 26479 16575
rect 26421 16535 26479 16541
rect 26786 16532 26792 16584
rect 26844 16532 26850 16584
rect 26878 16532 26884 16584
rect 26936 16572 26942 16584
rect 27617 16575 27675 16581
rect 27617 16572 27629 16575
rect 26936 16544 27629 16572
rect 26936 16532 26942 16544
rect 27617 16541 27629 16544
rect 27663 16541 27675 16575
rect 28092 16572 28120 16612
rect 28261 16609 28273 16643
rect 28307 16609 28319 16643
rect 28261 16603 28319 16609
rect 36446 16600 36452 16652
rect 36504 16600 36510 16652
rect 37568 16640 37596 16668
rect 38488 16640 38516 16668
rect 37568 16612 38424 16640
rect 38488 16612 38700 16640
rect 28353 16575 28411 16581
rect 28353 16572 28365 16575
rect 28092 16544 28365 16572
rect 27617 16535 27675 16541
rect 28353 16541 28365 16544
rect 28399 16572 28411 16575
rect 28534 16572 28540 16584
rect 28399 16544 28540 16572
rect 28399 16541 28411 16544
rect 28353 16535 28411 16541
rect 28534 16532 28540 16544
rect 28592 16532 28598 16584
rect 31202 16532 31208 16584
rect 31260 16572 31266 16584
rect 31570 16572 31576 16584
rect 31260 16544 31576 16572
rect 31260 16532 31266 16544
rect 31570 16532 31576 16544
rect 31628 16532 31634 16584
rect 33502 16572 33508 16584
rect 32982 16544 33508 16572
rect 33502 16532 33508 16544
rect 33560 16532 33566 16584
rect 33870 16532 33876 16584
rect 33928 16572 33934 16584
rect 36173 16575 36231 16581
rect 36173 16572 36185 16575
rect 33928 16544 36185 16572
rect 33928 16532 33934 16544
rect 36173 16541 36185 16544
rect 36219 16541 36231 16575
rect 38396 16572 38424 16612
rect 38519 16575 38577 16581
rect 38519 16572 38531 16575
rect 38396 16544 38531 16572
rect 36173 16535 36231 16541
rect 38519 16541 38531 16544
rect 38565 16541 38577 16575
rect 38672 16572 38700 16612
rect 40862 16600 40868 16652
rect 40920 16640 40926 16652
rect 41049 16643 41107 16649
rect 41049 16640 41061 16643
rect 40920 16612 41061 16640
rect 40920 16600 40926 16612
rect 41049 16609 41061 16612
rect 41095 16609 41107 16643
rect 41049 16603 41107 16609
rect 41322 16600 41328 16652
rect 41380 16600 41386 16652
rect 42794 16600 42800 16652
rect 42852 16640 42858 16652
rect 43073 16643 43131 16649
rect 43073 16640 43085 16643
rect 42852 16612 43085 16640
rect 42852 16600 42858 16612
rect 43073 16609 43085 16612
rect 43119 16609 43131 16643
rect 43073 16603 43131 16609
rect 43349 16643 43407 16649
rect 43349 16609 43361 16643
rect 43395 16640 43407 16643
rect 45002 16640 45008 16652
rect 43395 16612 45008 16640
rect 43395 16609 43407 16612
rect 43349 16603 43407 16609
rect 45002 16600 45008 16612
rect 45060 16600 45066 16652
rect 45296 16649 45324 16680
rect 45462 16668 45468 16720
rect 45520 16708 45526 16720
rect 45520 16680 45968 16708
rect 45520 16668 45526 16680
rect 45281 16643 45339 16649
rect 45281 16609 45293 16643
rect 45327 16640 45339 16643
rect 45738 16640 45744 16652
rect 45327 16612 45744 16640
rect 45327 16609 45339 16612
rect 45281 16603 45339 16609
rect 45738 16600 45744 16612
rect 45796 16600 45802 16652
rect 38749 16575 38807 16581
rect 38749 16572 38761 16575
rect 38672 16544 38761 16572
rect 38519 16535 38577 16541
rect 38749 16541 38761 16544
rect 38795 16541 38807 16575
rect 38930 16572 38936 16584
rect 38891 16544 38936 16572
rect 38749 16535 38807 16541
rect 38930 16532 38936 16544
rect 38988 16532 38994 16584
rect 39022 16532 39028 16584
rect 39080 16572 39086 16584
rect 39482 16572 39488 16584
rect 39080 16544 39488 16572
rect 39080 16532 39086 16544
rect 39482 16532 39488 16544
rect 39540 16532 39546 16584
rect 44358 16532 44364 16584
rect 44416 16572 44422 16584
rect 45940 16572 45968 16680
rect 46032 16640 46060 16736
rect 46753 16711 46811 16717
rect 46753 16677 46765 16711
rect 46799 16708 46811 16711
rect 48148 16708 48176 16748
rect 49970 16736 49976 16788
rect 50028 16776 50034 16788
rect 50801 16779 50859 16785
rect 50801 16776 50813 16779
rect 50028 16748 50813 16776
rect 50028 16736 50034 16748
rect 50801 16745 50813 16748
rect 50847 16745 50859 16779
rect 55306 16776 55312 16788
rect 50801 16739 50859 16745
rect 51046 16748 55312 16776
rect 51046 16708 51074 16748
rect 55306 16736 55312 16748
rect 55364 16776 55370 16788
rect 55585 16779 55643 16785
rect 55585 16776 55597 16779
rect 55364 16748 55597 16776
rect 55364 16736 55370 16748
rect 55585 16745 55597 16748
rect 55631 16745 55643 16779
rect 55585 16739 55643 16745
rect 46799 16680 46980 16708
rect 48148 16680 51074 16708
rect 46799 16677 46811 16680
rect 46753 16671 46811 16677
rect 46032 16612 46612 16640
rect 46106 16572 46112 16584
rect 44416 16558 44482 16572
rect 44416 16544 44496 16558
rect 45940 16544 46112 16572
rect 44416 16532 44422 16544
rect 23860 16476 25636 16504
rect 20864 16464 20870 16476
rect 12526 16396 12532 16448
rect 12584 16436 12590 16448
rect 14918 16436 14924 16448
rect 12584 16408 14924 16436
rect 12584 16396 12590 16408
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 17678 16396 17684 16448
rect 17736 16396 17742 16448
rect 18506 16396 18512 16448
rect 18564 16396 18570 16448
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 20901 16439 20959 16445
rect 20901 16436 20913 16439
rect 20772 16408 20913 16436
rect 20772 16396 20778 16408
rect 20901 16405 20913 16408
rect 20947 16436 20959 16439
rect 22738 16436 22744 16448
rect 20947 16408 22744 16436
rect 20947 16405 20959 16408
rect 20901 16399 20959 16405
rect 22738 16396 22744 16408
rect 22796 16436 22802 16448
rect 23216 16436 23244 16476
rect 25608 16448 25636 16476
rect 26510 16464 26516 16516
rect 26568 16464 26574 16516
rect 26602 16464 26608 16516
rect 26660 16464 26666 16516
rect 27338 16464 27344 16516
rect 27396 16504 27402 16516
rect 27433 16507 27491 16513
rect 27433 16504 27445 16507
rect 27396 16476 27445 16504
rect 27396 16464 27402 16476
rect 27433 16473 27445 16476
rect 27479 16473 27491 16507
rect 27433 16467 27491 16473
rect 27798 16464 27804 16516
rect 27856 16504 27862 16516
rect 28077 16507 28135 16513
rect 28077 16504 28089 16507
rect 27856 16476 28089 16504
rect 27856 16464 27862 16476
rect 28077 16473 28089 16476
rect 28123 16473 28135 16507
rect 28077 16467 28135 16473
rect 31846 16464 31852 16516
rect 31904 16464 31910 16516
rect 35434 16504 35440 16516
rect 33336 16476 35440 16504
rect 22796 16408 23244 16436
rect 23293 16439 23351 16445
rect 22796 16396 22802 16408
rect 23293 16405 23305 16439
rect 23339 16436 23351 16439
rect 23566 16436 23572 16448
rect 23339 16408 23572 16436
rect 23339 16405 23351 16408
rect 23293 16399 23351 16405
rect 23566 16396 23572 16408
rect 23624 16396 23630 16448
rect 23750 16396 23756 16448
rect 23808 16396 23814 16448
rect 23842 16396 23848 16448
rect 23900 16436 23906 16448
rect 24029 16439 24087 16445
rect 24029 16436 24041 16439
rect 23900 16408 24041 16436
rect 23900 16396 23906 16408
rect 24029 16405 24041 16408
rect 24075 16405 24087 16439
rect 24029 16399 24087 16405
rect 25590 16396 25596 16448
rect 25648 16436 25654 16448
rect 26053 16439 26111 16445
rect 26053 16436 26065 16439
rect 25648 16408 26065 16436
rect 25648 16396 25654 16408
rect 26053 16405 26065 16408
rect 26099 16405 26111 16439
rect 26620 16436 26648 16464
rect 27522 16436 27528 16448
rect 26620 16408 27528 16436
rect 26053 16399 26111 16405
rect 27522 16396 27528 16408
rect 27580 16396 27586 16448
rect 27890 16396 27896 16448
rect 27948 16436 27954 16448
rect 28537 16439 28595 16445
rect 28537 16436 28549 16439
rect 27948 16408 28549 16436
rect 27948 16396 27954 16408
rect 28537 16405 28549 16408
rect 28583 16405 28595 16439
rect 28537 16399 28595 16405
rect 32674 16396 32680 16448
rect 32732 16436 32738 16448
rect 33336 16445 33364 16476
rect 35434 16464 35440 16476
rect 35492 16464 35498 16516
rect 36078 16464 36084 16516
rect 36136 16504 36142 16516
rect 36538 16504 36544 16516
rect 36136 16476 36544 16504
rect 36136 16464 36142 16476
rect 36538 16464 36544 16476
rect 36596 16504 36602 16516
rect 38657 16507 38715 16513
rect 38657 16504 38669 16507
rect 36596 16476 36938 16504
rect 37936 16476 38669 16504
rect 36596 16464 36602 16476
rect 33321 16439 33379 16445
rect 33321 16436 33333 16439
rect 32732 16408 33333 16436
rect 32732 16396 32738 16408
rect 33321 16405 33333 16408
rect 33367 16405 33379 16439
rect 33321 16399 33379 16405
rect 33502 16396 33508 16448
rect 33560 16436 33566 16448
rect 35250 16436 35256 16448
rect 33560 16408 35256 16436
rect 33560 16396 33566 16408
rect 35250 16396 35256 16408
rect 35308 16396 35314 16448
rect 37090 16396 37096 16448
rect 37148 16436 37154 16448
rect 37936 16445 37964 16476
rect 38657 16473 38669 16476
rect 38703 16473 38715 16507
rect 39206 16504 39212 16516
rect 38657 16467 38715 16473
rect 39040 16476 39212 16504
rect 37921 16439 37979 16445
rect 37921 16436 37933 16439
rect 37148 16408 37933 16436
rect 37148 16396 37154 16408
rect 37921 16405 37933 16408
rect 37967 16405 37979 16439
rect 38672 16436 38700 16467
rect 39040 16436 39068 16476
rect 39206 16464 39212 16476
rect 39264 16464 39270 16516
rect 42550 16476 42653 16504
rect 42625 16448 42653 16476
rect 38672 16408 39068 16436
rect 37921 16399 37979 16405
rect 42610 16396 42616 16448
rect 42668 16436 42674 16448
rect 44266 16436 44272 16448
rect 42668 16408 44272 16436
rect 42668 16396 42674 16408
rect 44266 16396 44272 16408
rect 44324 16436 44330 16448
rect 44468 16436 44496 16544
rect 46106 16532 46112 16544
rect 46164 16532 46170 16584
rect 46201 16575 46259 16581
rect 46201 16541 46213 16575
rect 46247 16541 46259 16575
rect 46201 16535 46259 16541
rect 46216 16504 46244 16535
rect 46474 16532 46480 16584
rect 46532 16532 46538 16584
rect 46584 16581 46612 16612
rect 46842 16600 46848 16652
rect 46900 16600 46906 16652
rect 46952 16640 46980 16680
rect 47121 16643 47179 16649
rect 47121 16640 47133 16643
rect 46952 16612 47133 16640
rect 47121 16609 47133 16612
rect 47167 16609 47179 16643
rect 47121 16603 47179 16609
rect 47854 16600 47860 16652
rect 47912 16640 47918 16652
rect 50798 16640 50804 16652
rect 47912 16612 49004 16640
rect 47912 16600 47918 16612
rect 46569 16575 46627 16581
rect 46569 16541 46581 16575
rect 46615 16541 46627 16575
rect 46569 16535 46627 16541
rect 48222 16532 48228 16584
rect 48280 16532 48286 16584
rect 48866 16532 48872 16584
rect 48924 16532 48930 16584
rect 48976 16572 49004 16612
rect 49804 16612 50016 16640
rect 49237 16575 49295 16581
rect 49237 16572 49249 16575
rect 48976 16544 49249 16572
rect 49237 16541 49249 16544
rect 49283 16541 49295 16575
rect 49237 16535 49295 16541
rect 49326 16532 49332 16584
rect 49384 16572 49390 16584
rect 49513 16575 49571 16581
rect 49513 16572 49525 16575
rect 49384 16544 49525 16572
rect 49384 16532 49390 16544
rect 49513 16541 49525 16544
rect 49559 16541 49571 16575
rect 49513 16535 49571 16541
rect 47394 16504 47400 16516
rect 46216 16476 47400 16504
rect 47394 16464 47400 16476
rect 47452 16464 47458 16516
rect 44324 16408 44496 16436
rect 44324 16396 44330 16408
rect 47302 16396 47308 16448
rect 47360 16436 47366 16448
rect 48240 16436 48268 16532
rect 48608 16476 48820 16504
rect 47360 16408 48268 16436
rect 47360 16396 47366 16408
rect 48406 16396 48412 16448
rect 48464 16436 48470 16448
rect 48608 16445 48636 16476
rect 48593 16439 48651 16445
rect 48593 16436 48605 16439
rect 48464 16408 48605 16436
rect 48464 16396 48470 16408
rect 48593 16405 48605 16408
rect 48639 16405 48651 16439
rect 48593 16399 48651 16405
rect 48682 16396 48688 16448
rect 48740 16396 48746 16448
rect 48792 16436 48820 16476
rect 48958 16464 48964 16516
rect 49016 16464 49022 16516
rect 49050 16464 49056 16516
rect 49108 16464 49114 16516
rect 49605 16507 49663 16513
rect 49605 16504 49617 16507
rect 49160 16476 49617 16504
rect 49160 16436 49188 16476
rect 49605 16473 49617 16476
rect 49651 16473 49663 16507
rect 49605 16467 49663 16473
rect 49694 16464 49700 16516
rect 49752 16464 49758 16516
rect 48792 16408 49188 16436
rect 49329 16439 49387 16445
rect 49329 16405 49341 16439
rect 49375 16436 49387 16439
rect 49804 16436 49832 16612
rect 49881 16575 49939 16581
rect 49881 16541 49893 16575
rect 49927 16541 49939 16575
rect 49988 16572 50016 16612
rect 50540 16612 50804 16640
rect 50338 16581 50344 16584
rect 50157 16575 50215 16581
rect 50157 16572 50169 16575
rect 49988 16544 50169 16572
rect 49881 16535 49939 16541
rect 50157 16541 50169 16544
rect 50203 16541 50215 16575
rect 50157 16535 50215 16541
rect 50305 16575 50344 16581
rect 50305 16541 50317 16575
rect 50305 16535 50344 16541
rect 49375 16408 49832 16436
rect 49896 16436 49924 16535
rect 50338 16532 50344 16535
rect 50396 16532 50402 16584
rect 50540 16581 50568 16612
rect 50798 16600 50804 16612
rect 50856 16600 50862 16652
rect 51166 16600 51172 16652
rect 51224 16600 51230 16652
rect 51350 16600 51356 16652
rect 51408 16640 51414 16652
rect 51718 16640 51724 16652
rect 51408 16612 51724 16640
rect 51408 16600 51414 16612
rect 51718 16600 51724 16612
rect 51776 16640 51782 16652
rect 51997 16643 52055 16649
rect 51997 16640 52009 16643
rect 51776 16612 52009 16640
rect 51776 16600 51782 16612
rect 51997 16609 52009 16612
rect 52043 16609 52055 16643
rect 51997 16603 52055 16609
rect 52273 16643 52331 16649
rect 52273 16609 52285 16643
rect 52319 16640 52331 16643
rect 52638 16640 52644 16652
rect 52319 16612 52644 16640
rect 52319 16609 52331 16612
rect 52273 16603 52331 16609
rect 52638 16600 52644 16612
rect 52696 16600 52702 16652
rect 55600 16640 55628 16739
rect 55600 16612 56088 16640
rect 50706 16581 50712 16584
rect 50525 16575 50583 16581
rect 50525 16541 50537 16575
rect 50571 16541 50583 16575
rect 50525 16535 50583 16541
rect 50663 16575 50712 16581
rect 50663 16541 50675 16575
rect 50709 16541 50712 16575
rect 50663 16535 50712 16541
rect 50706 16532 50712 16535
rect 50764 16532 50770 16584
rect 51077 16575 51135 16581
rect 51077 16541 51089 16575
rect 51123 16572 51135 16575
rect 51184 16572 51212 16600
rect 51123 16544 51396 16572
rect 51123 16541 51135 16544
rect 51077 16535 51135 16541
rect 50062 16464 50068 16516
rect 50120 16504 50126 16516
rect 50433 16507 50491 16513
rect 50433 16504 50445 16507
rect 50120 16476 50445 16504
rect 50120 16464 50126 16476
rect 50433 16473 50445 16476
rect 50479 16473 50491 16507
rect 50982 16504 50988 16516
rect 50433 16467 50491 16473
rect 50724 16476 50988 16504
rect 50724 16436 50752 16476
rect 50982 16464 50988 16476
rect 51040 16464 51046 16516
rect 51169 16507 51227 16513
rect 51169 16473 51181 16507
rect 51215 16473 51227 16507
rect 51169 16467 51227 16473
rect 49896 16408 50752 16436
rect 49375 16405 49387 16408
rect 49329 16399 49387 16405
rect 50890 16396 50896 16448
rect 50948 16396 50954 16448
rect 51074 16396 51080 16448
rect 51132 16436 51138 16448
rect 51184 16436 51212 16467
rect 51258 16464 51264 16516
rect 51316 16464 51322 16516
rect 51132 16408 51212 16436
rect 51368 16436 51396 16544
rect 51442 16532 51448 16584
rect 51500 16532 51506 16584
rect 54202 16572 54208 16584
rect 53760 16544 54208 16572
rect 52546 16464 52552 16516
rect 52604 16504 52610 16516
rect 52604 16476 52762 16504
rect 52604 16464 52610 16476
rect 53760 16448 53788 16544
rect 54202 16532 54208 16544
rect 54260 16572 54266 16584
rect 54389 16575 54447 16581
rect 54389 16572 54401 16575
rect 54260 16544 54401 16572
rect 54260 16532 54266 16544
rect 54389 16541 54401 16544
rect 54435 16541 54447 16575
rect 54389 16535 54447 16541
rect 54754 16532 54760 16584
rect 54812 16532 54818 16584
rect 54938 16532 54944 16584
rect 54996 16532 55002 16584
rect 55030 16532 55036 16584
rect 55088 16532 55094 16584
rect 55766 16532 55772 16584
rect 55824 16532 55830 16584
rect 56060 16581 56088 16612
rect 56410 16600 56416 16652
rect 56468 16640 56474 16652
rect 56505 16643 56563 16649
rect 56505 16640 56517 16643
rect 56468 16612 56517 16640
rect 56468 16600 56474 16612
rect 56505 16609 56517 16612
rect 56551 16609 56563 16643
rect 56505 16603 56563 16609
rect 55953 16575 56011 16581
rect 55953 16541 55965 16575
rect 55999 16541 56011 16575
rect 55953 16535 56011 16541
rect 56045 16575 56103 16581
rect 56045 16541 56057 16575
rect 56091 16541 56103 16575
rect 56045 16535 56103 16541
rect 55674 16464 55680 16516
rect 55732 16504 55738 16516
rect 55968 16504 55996 16535
rect 56134 16532 56140 16584
rect 56192 16532 56198 16584
rect 77846 16572 77852 16584
rect 64846 16544 77852 16572
rect 55732 16476 55996 16504
rect 56413 16507 56471 16513
rect 55732 16464 55738 16476
rect 56413 16473 56425 16507
rect 56459 16504 56471 16507
rect 56750 16507 56808 16513
rect 56750 16504 56762 16507
rect 56459 16476 56762 16504
rect 56459 16473 56471 16476
rect 56413 16467 56471 16473
rect 56750 16473 56762 16476
rect 56796 16473 56808 16507
rect 56750 16467 56808 16473
rect 51442 16436 51448 16448
rect 51368 16408 51448 16436
rect 51132 16396 51138 16408
rect 51442 16396 51448 16408
rect 51500 16436 51506 16448
rect 51537 16439 51595 16445
rect 51537 16436 51549 16439
rect 51500 16408 51549 16436
rect 51500 16396 51506 16408
rect 51537 16405 51549 16408
rect 51583 16405 51595 16439
rect 51537 16399 51595 16405
rect 53742 16396 53748 16448
rect 53800 16396 53806 16448
rect 53834 16396 53840 16448
rect 53892 16396 53898 16448
rect 54570 16396 54576 16448
rect 54628 16396 54634 16448
rect 57885 16439 57943 16445
rect 57885 16405 57897 16439
rect 57931 16436 57943 16439
rect 57974 16436 57980 16448
rect 57931 16408 57980 16436
rect 57931 16405 57943 16408
rect 57885 16399 57943 16405
rect 57974 16396 57980 16408
rect 58032 16436 58038 16448
rect 64846 16436 64874 16544
rect 77846 16532 77852 16544
rect 77904 16532 77910 16584
rect 58032 16408 64874 16436
rect 58032 16396 58038 16408
rect 1104 16346 78844 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 66314 16346
rect 66366 16294 66378 16346
rect 66430 16294 66442 16346
rect 66494 16294 66506 16346
rect 66558 16294 66570 16346
rect 66622 16294 78844 16346
rect 1104 16272 78844 16294
rect 9490 16232 9496 16244
rect 8588 16204 9496 16232
rect 1302 16056 1308 16108
rect 1360 16096 1366 16108
rect 8588 16105 8616 16204
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 11440 16204 11744 16232
rect 11440 16164 11468 16204
rect 10074 16136 11468 16164
rect 11716 16164 11744 16204
rect 12618 16192 12624 16244
rect 12676 16232 12682 16244
rect 13265 16235 13323 16241
rect 13265 16232 13277 16235
rect 12676 16204 13277 16232
rect 12676 16192 12682 16204
rect 13265 16201 13277 16204
rect 13311 16232 13323 16235
rect 13354 16232 13360 16244
rect 13311 16204 13360 16232
rect 13311 16201 13323 16204
rect 13265 16195 13323 16201
rect 13354 16192 13360 16204
rect 13412 16192 13418 16244
rect 17034 16192 17040 16244
rect 17092 16192 17098 16244
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 17368 16204 17509 16232
rect 17368 16192 17374 16204
rect 17497 16201 17509 16204
rect 17543 16201 17555 16235
rect 17497 16195 17555 16201
rect 20806 16192 20812 16244
rect 20864 16192 20870 16244
rect 23198 16192 23204 16244
rect 23256 16232 23262 16244
rect 23256 16204 23704 16232
rect 23256 16192 23262 16204
rect 12250 16164 12256 16176
rect 11716 16136 12256 16164
rect 12250 16124 12256 16136
rect 12308 16124 12314 16176
rect 14918 16124 14924 16176
rect 14976 16124 14982 16176
rect 17221 16167 17279 16173
rect 17221 16133 17233 16167
rect 17267 16164 17279 16167
rect 18506 16164 18512 16176
rect 17267 16136 18512 16164
rect 17267 16133 17279 16136
rect 17221 16127 17279 16133
rect 18506 16124 18512 16136
rect 18564 16124 18570 16176
rect 23290 16164 23296 16176
rect 20364 16136 23296 16164
rect 20364 16108 20392 16136
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 1360 16068 1409 16096
rect 1360 16056 1366 16068
rect 1397 16065 1409 16068
rect 1443 16096 1455 16099
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1443 16068 1685 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16065 8631 16099
rect 8573 16059 8631 16065
rect 11514 16056 11520 16108
rect 11572 16056 11578 16108
rect 17126 16056 17132 16108
rect 17184 16056 17190 16108
rect 17678 16056 17684 16108
rect 17736 16096 17742 16108
rect 18049 16099 18107 16105
rect 18049 16096 18061 16099
rect 17736 16068 18061 16096
rect 17736 16056 17742 16068
rect 18049 16065 18061 16068
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 20346 16056 20352 16108
rect 20404 16056 20410 16108
rect 20533 16099 20591 16105
rect 20533 16065 20545 16099
rect 20579 16096 20591 16099
rect 20622 16096 20628 16108
rect 20579 16068 20628 16096
rect 20579 16065 20591 16068
rect 20533 16059 20591 16065
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 20714 16056 20720 16108
rect 20772 16056 20778 16108
rect 20806 16056 20812 16108
rect 20864 16096 20870 16108
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 20864 16068 21097 16096
rect 20864 16056 20870 16068
rect 21085 16065 21097 16068
rect 21131 16096 21143 16099
rect 21450 16096 21456 16108
rect 21131 16068 21456 16096
rect 21131 16065 21143 16068
rect 21085 16059 21143 16065
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 23216 16105 23244 16136
rect 23290 16124 23296 16136
rect 23348 16124 23354 16176
rect 23676 16105 23704 16204
rect 24578 16192 24584 16244
rect 24636 16192 24642 16244
rect 24762 16192 24768 16244
rect 24820 16192 24826 16244
rect 26053 16235 26111 16241
rect 26053 16201 26065 16235
rect 26099 16232 26111 16235
rect 26326 16232 26332 16244
rect 26099 16204 26332 16232
rect 26099 16201 26111 16204
rect 26053 16195 26111 16201
rect 26326 16192 26332 16204
rect 26384 16192 26390 16244
rect 27246 16192 27252 16244
rect 27304 16232 27310 16244
rect 27304 16204 27476 16232
rect 27304 16192 27310 16204
rect 23842 16124 23848 16176
rect 23900 16164 23906 16176
rect 26786 16164 26792 16176
rect 23900 16136 26792 16164
rect 23900 16124 23906 16136
rect 23201 16099 23259 16105
rect 23201 16065 23213 16099
rect 23247 16065 23259 16099
rect 23201 16059 23259 16065
rect 23385 16099 23443 16105
rect 23385 16065 23397 16099
rect 23431 16096 23443 16099
rect 23477 16099 23535 16105
rect 23477 16096 23489 16099
rect 23431 16068 23489 16096
rect 23431 16065 23443 16068
rect 23385 16059 23443 16065
rect 23477 16065 23489 16068
rect 23523 16065 23535 16099
rect 23477 16059 23535 16065
rect 23661 16099 23719 16105
rect 23661 16065 23673 16099
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 24029 16099 24087 16105
rect 24029 16065 24041 16099
rect 24075 16096 24087 16099
rect 24075 16068 24256 16096
rect 24075 16065 24087 16068
rect 24029 16059 24087 16065
rect 8294 15988 8300 16040
rect 8352 16028 8358 16040
rect 8849 16031 8907 16037
rect 8849 16028 8861 16031
rect 8352 16000 8861 16028
rect 8352 15988 8358 16000
rect 8849 15997 8861 16000
rect 8895 15997 8907 16031
rect 8849 15991 8907 15997
rect 11790 15988 11796 16040
rect 11848 15988 11854 16040
rect 12250 15988 12256 16040
rect 12308 16028 12314 16040
rect 12526 16028 12532 16040
rect 12308 16000 12532 16028
rect 12308 15988 12314 16000
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 13630 15988 13636 16040
rect 13688 15988 13694 16040
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 16028 13967 16031
rect 14274 16028 14280 16040
rect 13955 16000 14280 16028
rect 13955 15997 13967 16000
rect 13909 15991 13967 15997
rect 14274 15988 14280 16000
rect 14332 15988 14338 16040
rect 15381 16031 15439 16037
rect 15381 15997 15393 16031
rect 15427 16028 15439 16031
rect 15746 16028 15752 16040
rect 15427 16000 15752 16028
rect 15427 15997 15439 16000
rect 15381 15991 15439 15997
rect 15746 15988 15752 16000
rect 15804 16028 15810 16040
rect 16025 16031 16083 16037
rect 16025 16028 16037 16031
rect 15804 16000 16037 16028
rect 15804 15988 15810 16000
rect 16025 15997 16037 16000
rect 16071 15997 16083 16031
rect 16025 15991 16083 15997
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 16028 20959 16031
rect 20990 16028 20996 16040
rect 20947 16000 20996 16028
rect 20947 15997 20959 16000
rect 20901 15991 20959 15997
rect 20990 15988 20996 16000
rect 21048 15988 21054 16040
rect 22922 15988 22928 16040
rect 22980 16028 22986 16040
rect 23400 16028 23428 16059
rect 22980 16000 23428 16028
rect 22980 15988 22986 16000
rect 24118 15988 24124 16040
rect 24176 15988 24182 16040
rect 24228 16037 24256 16068
rect 24394 16056 24400 16108
rect 24452 16096 24458 16108
rect 24640 16099 24698 16105
rect 24640 16096 24652 16099
rect 24452 16068 24652 16096
rect 24452 16056 24458 16068
rect 24640 16065 24652 16068
rect 24686 16096 24698 16099
rect 24762 16096 24768 16108
rect 24686 16068 24768 16096
rect 24686 16065 24698 16068
rect 24640 16059 24698 16065
rect 24762 16056 24768 16068
rect 24820 16056 24826 16108
rect 25590 16056 25596 16108
rect 25648 16056 25654 16108
rect 25792 16105 25820 16136
rect 26786 16124 26792 16136
rect 26844 16124 26850 16176
rect 27338 16164 27344 16176
rect 26896 16136 27344 16164
rect 25777 16099 25835 16105
rect 25777 16065 25789 16099
rect 25823 16065 25835 16099
rect 25777 16059 25835 16065
rect 25869 16099 25927 16105
rect 25869 16065 25881 16099
rect 25915 16096 25927 16099
rect 25958 16096 25964 16108
rect 25915 16068 25964 16096
rect 25915 16065 25927 16068
rect 25869 16059 25927 16065
rect 25958 16056 25964 16068
rect 26016 16056 26022 16108
rect 26896 16096 26924 16136
rect 27338 16124 27344 16136
rect 27396 16124 27402 16176
rect 27448 16173 27476 16204
rect 27522 16192 27528 16244
rect 27580 16232 27586 16244
rect 27985 16235 28043 16241
rect 27985 16232 27997 16235
rect 27580 16204 27997 16232
rect 27580 16192 27586 16204
rect 27985 16201 27997 16204
rect 28031 16201 28043 16235
rect 27985 16195 28043 16201
rect 31846 16192 31852 16244
rect 31904 16232 31910 16244
rect 32125 16235 32183 16241
rect 32125 16232 32137 16235
rect 31904 16204 32137 16232
rect 31904 16192 31910 16204
rect 32125 16201 32137 16204
rect 32171 16201 32183 16235
rect 32125 16195 32183 16201
rect 34790 16192 34796 16244
rect 34848 16232 34854 16244
rect 35621 16235 35679 16241
rect 35621 16232 35633 16235
rect 34848 16204 35633 16232
rect 34848 16192 34854 16204
rect 35621 16201 35633 16204
rect 35667 16201 35679 16235
rect 35621 16195 35679 16201
rect 38194 16192 38200 16244
rect 38252 16232 38258 16244
rect 41506 16232 41512 16244
rect 38252 16204 41512 16232
rect 38252 16192 38258 16204
rect 41506 16192 41512 16204
rect 41564 16232 41570 16244
rect 42518 16232 42524 16244
rect 41564 16204 42524 16232
rect 41564 16192 41570 16204
rect 42518 16192 42524 16204
rect 42576 16192 42582 16244
rect 44450 16192 44456 16244
rect 44508 16232 44514 16244
rect 44729 16235 44787 16241
rect 44729 16232 44741 16235
rect 44508 16204 44741 16232
rect 44508 16192 44514 16204
rect 44729 16201 44741 16204
rect 44775 16201 44787 16235
rect 44729 16195 44787 16201
rect 27433 16167 27491 16173
rect 27433 16133 27445 16167
rect 27479 16164 27491 16167
rect 29178 16164 29184 16176
rect 27479 16136 29184 16164
rect 27479 16133 27491 16136
rect 27433 16127 27491 16133
rect 26252 16068 26924 16096
rect 24213 16031 24271 16037
rect 24213 15997 24225 16031
rect 24259 16028 24271 16031
rect 26252 16028 26280 16068
rect 27154 16056 27160 16108
rect 27212 16096 27218 16108
rect 27249 16099 27307 16105
rect 27249 16096 27261 16099
rect 27212 16068 27261 16096
rect 27212 16056 27218 16068
rect 27249 16065 27261 16068
rect 27295 16065 27307 16099
rect 27249 16059 27307 16065
rect 27982 16056 27988 16108
rect 28040 16056 28046 16108
rect 28184 16105 28212 16136
rect 29178 16124 29184 16136
rect 29236 16124 29242 16176
rect 34149 16167 34207 16173
rect 34149 16133 34161 16167
rect 34195 16164 34207 16167
rect 34238 16164 34244 16176
rect 34195 16136 34244 16164
rect 34195 16133 34207 16136
rect 34149 16127 34207 16133
rect 34238 16124 34244 16136
rect 34296 16124 34302 16176
rect 28169 16099 28227 16105
rect 28169 16065 28181 16099
rect 28215 16065 28227 16099
rect 28169 16059 28227 16065
rect 28445 16099 28503 16105
rect 28445 16065 28457 16099
rect 28491 16096 28503 16099
rect 28994 16096 29000 16108
rect 28491 16068 29000 16096
rect 28491 16065 28503 16068
rect 28445 16059 28503 16065
rect 28994 16056 29000 16068
rect 29052 16096 29058 16108
rect 29546 16096 29552 16108
rect 29052 16068 29552 16096
rect 29052 16056 29058 16068
rect 29546 16056 29552 16068
rect 29604 16056 29610 16108
rect 32030 16056 32036 16108
rect 32088 16096 32094 16108
rect 32309 16099 32367 16105
rect 32309 16096 32321 16099
rect 32088 16068 32321 16096
rect 32088 16056 32094 16068
rect 32309 16065 32321 16068
rect 32355 16065 32367 16099
rect 32309 16059 32367 16065
rect 32398 16056 32404 16108
rect 32456 16056 32462 16108
rect 32674 16056 32680 16108
rect 32732 16056 32738 16108
rect 33226 16056 33232 16108
rect 33284 16096 33290 16108
rect 33870 16096 33876 16108
rect 33284 16068 33876 16096
rect 33284 16056 33290 16068
rect 33870 16056 33876 16068
rect 33928 16056 33934 16108
rect 35250 16056 35256 16108
rect 35308 16056 35314 16108
rect 44744 16096 44772 16195
rect 44910 16192 44916 16244
rect 44968 16232 44974 16244
rect 45646 16232 45652 16244
rect 44968 16204 45652 16232
rect 44968 16192 44974 16204
rect 45388 16173 45416 16204
rect 45646 16192 45652 16204
rect 45704 16192 45710 16244
rect 46014 16232 46020 16244
rect 45756 16204 46020 16232
rect 45373 16167 45431 16173
rect 45373 16133 45385 16167
rect 45419 16133 45431 16167
rect 45756 16164 45784 16204
rect 46014 16192 46020 16204
rect 46072 16192 46078 16244
rect 46201 16235 46259 16241
rect 46201 16201 46213 16235
rect 46247 16232 46259 16235
rect 46474 16232 46480 16244
rect 46247 16204 46480 16232
rect 46247 16201 46259 16204
rect 46201 16195 46259 16201
rect 46474 16192 46480 16204
rect 46532 16192 46538 16244
rect 47305 16235 47363 16241
rect 47305 16232 47317 16235
rect 46676 16204 47317 16232
rect 45373 16127 45431 16133
rect 45664 16136 45784 16164
rect 45097 16099 45155 16105
rect 45097 16096 45109 16099
rect 44744 16068 45109 16096
rect 45097 16065 45109 16068
rect 45143 16065 45155 16099
rect 45097 16059 45155 16065
rect 45245 16099 45303 16105
rect 45245 16065 45257 16099
rect 45291 16096 45303 16099
rect 45291 16065 45324 16096
rect 45245 16059 45324 16065
rect 24259 16000 26280 16028
rect 24259 15997 24271 16000
rect 24213 15991 24271 15997
rect 26510 15988 26516 16040
rect 26568 16028 26574 16040
rect 32585 16031 32643 16037
rect 26568 16000 31754 16028
rect 26568 15988 26574 16000
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 8110 15960 8116 15972
rect 1627 15932 8116 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 8110 15920 8116 15932
rect 8168 15920 8174 15972
rect 16114 15920 16120 15972
rect 16172 15960 16178 15972
rect 16853 15963 16911 15969
rect 16853 15960 16865 15963
rect 16172 15932 16865 15960
rect 16172 15920 16178 15932
rect 16853 15929 16865 15932
rect 16899 15929 16911 15963
rect 16853 15923 16911 15929
rect 23937 15963 23995 15969
rect 23937 15929 23949 15963
rect 23983 15960 23995 15963
rect 27246 15960 27252 15972
rect 23983 15932 27252 15960
rect 23983 15929 23995 15932
rect 23937 15923 23995 15929
rect 27246 15920 27252 15932
rect 27304 15920 27310 15972
rect 27706 15920 27712 15972
rect 27764 15960 27770 15972
rect 30006 15960 30012 15972
rect 27764 15932 30012 15960
rect 27764 15920 27770 15932
rect 30006 15920 30012 15932
rect 30064 15920 30070 15972
rect 31726 15960 31754 16000
rect 32585 15997 32597 16031
rect 32631 16028 32643 16031
rect 33410 16028 33416 16040
rect 32631 16000 33416 16028
rect 32631 15997 32643 16000
rect 32585 15991 32643 15997
rect 33410 15988 33416 16000
rect 33468 15988 33474 16040
rect 36998 16028 37004 16040
rect 33980 16000 37004 16028
rect 33980 15960 34008 16000
rect 36998 15988 37004 16000
rect 37056 15988 37062 16040
rect 45296 16028 45324 16059
rect 45462 16056 45468 16108
rect 45520 16056 45526 16108
rect 45562 16099 45620 16105
rect 45562 16065 45574 16099
rect 45608 16096 45620 16099
rect 45664 16096 45692 16136
rect 45608 16068 45692 16096
rect 45608 16065 45620 16068
rect 45562 16059 45620 16065
rect 45738 16056 45744 16108
rect 45796 16096 45802 16108
rect 45833 16099 45891 16105
rect 45833 16096 45845 16099
rect 45796 16068 45845 16096
rect 45796 16056 45802 16068
rect 45833 16065 45845 16068
rect 45879 16065 45891 16099
rect 45833 16059 45891 16065
rect 46017 16099 46075 16105
rect 46017 16065 46029 16099
rect 46063 16096 46075 16099
rect 46198 16096 46204 16108
rect 46063 16068 46204 16096
rect 46063 16065 46075 16068
rect 46017 16059 46075 16065
rect 46198 16056 46204 16068
rect 46256 16096 46262 16108
rect 46676 16105 46704 16204
rect 47305 16201 47317 16204
rect 47351 16201 47363 16235
rect 47305 16195 47363 16201
rect 47394 16192 47400 16244
rect 47452 16232 47458 16244
rect 47581 16235 47639 16241
rect 47581 16232 47593 16235
rect 47452 16204 47593 16232
rect 47452 16192 47458 16204
rect 47581 16201 47593 16204
rect 47627 16201 47639 16235
rect 47581 16195 47639 16201
rect 48777 16235 48835 16241
rect 48777 16201 48789 16235
rect 48823 16232 48835 16235
rect 50154 16232 50160 16244
rect 48823 16204 49924 16232
rect 48823 16201 48835 16204
rect 48777 16195 48835 16201
rect 46753 16167 46811 16173
rect 46753 16133 46765 16167
rect 46799 16164 46811 16167
rect 47854 16164 47860 16176
rect 46799 16136 47860 16164
rect 46799 16133 46811 16136
rect 46753 16127 46811 16133
rect 47854 16124 47860 16136
rect 47912 16124 47918 16176
rect 48406 16164 48412 16176
rect 48240 16136 48412 16164
rect 48240 16105 48268 16136
rect 48406 16124 48412 16136
rect 48464 16124 48470 16176
rect 49053 16167 49111 16173
rect 49053 16133 49065 16167
rect 49099 16164 49111 16167
rect 49694 16164 49700 16176
rect 49099 16136 49700 16164
rect 49099 16133 49111 16136
rect 49053 16127 49111 16133
rect 49694 16124 49700 16136
rect 49752 16124 49758 16176
rect 49896 16173 49924 16204
rect 49988 16204 50160 16232
rect 49881 16167 49939 16173
rect 49881 16133 49893 16167
rect 49927 16133 49939 16167
rect 49881 16127 49939 16133
rect 49988 16164 50016 16204
rect 50154 16192 50160 16204
rect 50212 16192 50218 16244
rect 50614 16192 50620 16244
rect 50672 16232 50678 16244
rect 50672 16204 50752 16232
rect 50672 16192 50678 16204
rect 50724 16173 50752 16204
rect 50798 16192 50804 16244
rect 50856 16232 50862 16244
rect 50856 16204 52041 16232
rect 50856 16192 50862 16204
rect 50709 16167 50767 16173
rect 49988 16136 50385 16164
rect 46293 16099 46351 16105
rect 46293 16096 46305 16099
rect 46256 16068 46305 16096
rect 46256 16056 46262 16068
rect 46293 16065 46305 16068
rect 46339 16096 46351 16099
rect 46661 16099 46719 16105
rect 46661 16096 46673 16099
rect 46339 16068 46673 16096
rect 46339 16065 46351 16068
rect 46293 16059 46351 16065
rect 46661 16065 46673 16068
rect 46707 16065 46719 16099
rect 46661 16059 46719 16065
rect 46845 16099 46903 16105
rect 46845 16065 46857 16099
rect 46891 16065 46903 16099
rect 46845 16059 46903 16065
rect 47029 16099 47087 16105
rect 47029 16065 47041 16099
rect 47075 16096 47087 16099
rect 48225 16099 48283 16105
rect 48225 16096 48237 16099
rect 47075 16068 48237 16096
rect 47075 16065 47087 16068
rect 47029 16059 47087 16065
rect 48225 16065 48237 16068
rect 48271 16065 48283 16099
rect 48225 16059 48283 16065
rect 48317 16099 48375 16105
rect 48317 16065 48329 16099
rect 48363 16096 48375 16099
rect 48498 16096 48504 16108
rect 48363 16068 48504 16096
rect 48363 16065 48375 16068
rect 48317 16059 48375 16065
rect 45756 16028 45784 16056
rect 45296 16000 45784 16028
rect 45922 15988 45928 16040
rect 45980 16028 45986 16040
rect 46860 16028 46888 16059
rect 48498 16056 48504 16068
rect 48556 16056 48562 16108
rect 48590 16056 48596 16108
rect 48648 16056 48654 16108
rect 49510 16056 49516 16108
rect 49568 16056 49574 16108
rect 49789 16099 49847 16105
rect 49789 16065 49801 16099
rect 49835 16096 49847 16099
rect 49988 16096 50016 16136
rect 49835 16068 50016 16096
rect 50157 16099 50215 16105
rect 49835 16065 49847 16068
rect 49789 16059 49847 16065
rect 50157 16065 50169 16099
rect 50203 16096 50215 16099
rect 50246 16096 50252 16108
rect 50203 16068 50252 16096
rect 50203 16065 50215 16068
rect 50157 16059 50215 16065
rect 50246 16056 50252 16068
rect 50304 16056 50310 16108
rect 45980 16000 46888 16028
rect 48409 16031 48467 16037
rect 45980 15988 45986 16000
rect 48409 15997 48421 16031
rect 48455 15997 48467 16031
rect 48409 15991 48467 15997
rect 31726 15932 34008 15960
rect 35250 15920 35256 15972
rect 35308 15960 35314 15972
rect 35805 15963 35863 15969
rect 35805 15960 35817 15963
rect 35308 15932 35817 15960
rect 35308 15920 35314 15932
rect 35805 15929 35817 15932
rect 35851 15960 35863 15963
rect 36078 15960 36084 15972
rect 35851 15932 36084 15960
rect 35851 15929 35863 15932
rect 35805 15923 35863 15929
rect 36078 15920 36084 15932
rect 36136 15920 36142 15972
rect 45741 15963 45799 15969
rect 45741 15929 45753 15963
rect 45787 15960 45799 15963
rect 48424 15960 48452 15991
rect 49050 15988 49056 16040
rect 49108 16028 49114 16040
rect 49418 16028 49424 16040
rect 49108 16000 49424 16028
rect 49108 15988 49114 16000
rect 49418 15988 49424 16000
rect 49476 15988 49482 16040
rect 50065 16031 50123 16037
rect 50065 15997 50077 16031
rect 50111 15997 50123 16031
rect 50357 16028 50385 16136
rect 50709 16133 50721 16167
rect 50755 16133 50767 16167
rect 50709 16127 50767 16133
rect 50430 16056 50436 16108
rect 50488 16105 50494 16108
rect 50890 16105 50896 16108
rect 50488 16099 50511 16105
rect 50499 16065 50511 16099
rect 50488 16059 50511 16065
rect 50617 16099 50675 16105
rect 50617 16065 50629 16099
rect 50663 16065 50675 16099
rect 50617 16059 50675 16065
rect 50847 16099 50896 16105
rect 50847 16065 50859 16099
rect 50893 16065 50896 16099
rect 50847 16059 50896 16065
rect 50488 16056 50494 16059
rect 50632 16028 50660 16059
rect 50890 16056 50896 16059
rect 50948 16056 50954 16108
rect 51067 16099 51125 16105
rect 51067 16065 51079 16099
rect 51113 16065 51125 16099
rect 51067 16059 51125 16065
rect 50706 16028 50712 16040
rect 50357 16000 50712 16028
rect 50065 15991 50123 15997
rect 45787 15932 48452 15960
rect 45787 15929 45799 15932
rect 45741 15923 45799 15929
rect 10321 15895 10379 15901
rect 10321 15861 10333 15895
rect 10367 15892 10379 15895
rect 14642 15892 14648 15904
rect 10367 15864 14648 15892
rect 10367 15861 10379 15864
rect 10321 15855 10379 15861
rect 14642 15852 14648 15864
rect 14700 15852 14706 15904
rect 15470 15852 15476 15904
rect 15528 15852 15534 15904
rect 17402 15852 17408 15904
rect 17460 15852 17466 15904
rect 20530 15852 20536 15904
rect 20588 15852 20594 15904
rect 21082 15852 21088 15904
rect 21140 15852 21146 15904
rect 23382 15852 23388 15904
rect 23440 15852 23446 15904
rect 25866 15852 25872 15904
rect 25924 15852 25930 15904
rect 26326 15852 26332 15904
rect 26384 15892 26390 15904
rect 27065 15895 27123 15901
rect 27065 15892 27077 15895
rect 26384 15864 27077 15892
rect 26384 15852 26390 15864
rect 27065 15861 27077 15864
rect 27111 15861 27123 15895
rect 27065 15855 27123 15861
rect 28629 15895 28687 15901
rect 28629 15861 28641 15895
rect 28675 15892 28687 15895
rect 29546 15892 29552 15904
rect 28675 15864 29552 15892
rect 28675 15861 28687 15864
rect 28629 15855 28687 15861
rect 29546 15852 29552 15864
rect 29604 15852 29610 15904
rect 35986 15852 35992 15904
rect 36044 15852 36050 15904
rect 39666 15852 39672 15904
rect 39724 15892 39730 15904
rect 43346 15892 43352 15904
rect 39724 15864 43352 15892
rect 39724 15852 39730 15864
rect 43346 15852 43352 15864
rect 43404 15852 43410 15904
rect 46106 15852 46112 15904
rect 46164 15892 46170 15904
rect 46477 15895 46535 15901
rect 46477 15892 46489 15895
rect 46164 15864 46489 15892
rect 46164 15852 46170 15864
rect 46477 15861 46489 15864
rect 46523 15861 46535 15895
rect 46477 15855 46535 15861
rect 46750 15852 46756 15904
rect 46808 15892 46814 15904
rect 47121 15895 47179 15901
rect 47121 15892 47133 15895
rect 46808 15864 47133 15892
rect 46808 15852 46814 15864
rect 47121 15861 47133 15864
rect 47167 15861 47179 15895
rect 47121 15855 47179 15861
rect 48593 15895 48651 15901
rect 48593 15861 48605 15895
rect 48639 15892 48651 15895
rect 48682 15892 48688 15904
rect 48639 15864 48688 15892
rect 48639 15861 48651 15864
rect 48593 15855 48651 15861
rect 48682 15852 48688 15864
rect 48740 15852 48746 15904
rect 49237 15895 49295 15901
rect 49237 15861 49249 15895
rect 49283 15892 49295 15895
rect 49326 15892 49332 15904
rect 49283 15864 49332 15892
rect 49283 15861 49295 15864
rect 49237 15855 49295 15861
rect 49326 15852 49332 15864
rect 49384 15852 49390 15904
rect 49970 15852 49976 15904
rect 50028 15852 50034 15904
rect 50080 15892 50108 15991
rect 50706 15988 50712 16000
rect 50764 15988 50770 16040
rect 51092 16028 51120 16059
rect 51166 16056 51172 16108
rect 51224 16056 51230 16108
rect 51350 16056 51356 16108
rect 51408 16056 51414 16108
rect 51445 16099 51503 16105
rect 51445 16065 51457 16099
rect 51491 16096 51503 16099
rect 51534 16096 51540 16108
rect 51491 16068 51540 16096
rect 51491 16065 51503 16068
rect 51445 16059 51503 16065
rect 51534 16056 51540 16068
rect 51592 16096 51598 16108
rect 51721 16099 51779 16105
rect 51721 16096 51733 16099
rect 51592 16068 51733 16096
rect 51592 16056 51598 16068
rect 51721 16065 51733 16068
rect 51767 16065 51779 16099
rect 51721 16059 51779 16065
rect 51902 16056 51908 16108
rect 51960 16056 51966 16108
rect 52013 16105 52041 16204
rect 52362 16192 52368 16244
rect 52420 16192 52426 16244
rect 52549 16235 52607 16241
rect 52549 16201 52561 16235
rect 52595 16201 52607 16235
rect 52549 16195 52607 16201
rect 52181 16167 52239 16173
rect 52181 16133 52193 16167
rect 52227 16164 52239 16167
rect 52380 16164 52408 16192
rect 52227 16136 52408 16164
rect 52227 16133 52239 16136
rect 52181 16127 52239 16133
rect 51998 16099 52056 16105
rect 51998 16065 52010 16099
rect 52044 16065 52056 16099
rect 51998 16059 52056 16065
rect 51000 16000 51120 16028
rect 50341 15963 50399 15969
rect 50341 15929 50353 15963
rect 50387 15960 50399 15963
rect 50430 15960 50436 15972
rect 50387 15932 50436 15960
rect 50387 15929 50399 15932
rect 50341 15923 50399 15929
rect 50430 15920 50436 15932
rect 50488 15920 50494 15972
rect 51000 15969 51028 16000
rect 50985 15963 51043 15969
rect 50985 15929 50997 15963
rect 51031 15929 51043 15963
rect 52013 15960 52041 16059
rect 52270 16056 52276 16108
rect 52328 16056 52334 16108
rect 52454 16105 52460 16108
rect 52411 16099 52460 16105
rect 52411 16065 52423 16099
rect 52457 16065 52460 16099
rect 52411 16059 52460 16065
rect 52454 16056 52460 16059
rect 52512 16056 52518 16108
rect 52564 16096 52592 16195
rect 52638 16192 52644 16244
rect 52696 16232 52702 16244
rect 52733 16235 52791 16241
rect 52733 16232 52745 16235
rect 52696 16204 52745 16232
rect 52696 16192 52702 16204
rect 52733 16201 52745 16204
rect 52779 16201 52791 16235
rect 54938 16232 54944 16244
rect 52733 16195 52791 16201
rect 53208 16204 54944 16232
rect 53208 16164 53236 16204
rect 54938 16192 54944 16204
rect 54996 16192 55002 16244
rect 56134 16192 56140 16244
rect 56192 16232 56198 16244
rect 57057 16235 57115 16241
rect 57057 16232 57069 16235
rect 56192 16204 57069 16232
rect 56192 16192 56198 16204
rect 57057 16201 57069 16204
rect 57103 16201 57115 16235
rect 57057 16195 57115 16201
rect 57974 16192 57980 16244
rect 58032 16192 58038 16244
rect 53116 16136 53236 16164
rect 53116 16105 53144 16136
rect 53374 16124 53380 16176
rect 53432 16124 53438 16176
rect 54570 16124 54576 16176
rect 54628 16164 54634 16176
rect 54665 16167 54723 16173
rect 54665 16164 54677 16167
rect 54628 16136 54677 16164
rect 54628 16124 54634 16136
rect 54665 16133 54677 16136
rect 54711 16133 54723 16167
rect 54665 16127 54723 16133
rect 55674 16124 55680 16176
rect 55732 16124 55738 16176
rect 52917 16099 52975 16105
rect 52917 16096 52929 16099
rect 52564 16068 52929 16096
rect 52917 16065 52929 16068
rect 52963 16065 52975 16099
rect 52917 16059 52975 16065
rect 53101 16099 53159 16105
rect 53101 16065 53113 16099
rect 53147 16065 53159 16099
rect 53101 16059 53159 16065
rect 53193 16099 53251 16105
rect 53193 16065 53205 16099
rect 53239 16096 53251 16099
rect 53834 16096 53840 16108
rect 53239 16068 53840 16096
rect 53239 16065 53251 16068
rect 53193 16059 53251 16065
rect 53834 16056 53840 16068
rect 53892 16056 53898 16108
rect 57701 16099 57759 16105
rect 57701 16065 57713 16099
rect 57747 16096 57759 16099
rect 57992 16096 58020 16192
rect 57747 16068 58020 16096
rect 57747 16065 57759 16068
rect 57701 16059 57759 16065
rect 54018 15988 54024 16040
rect 54076 16028 54082 16040
rect 54113 16031 54171 16037
rect 54113 16028 54125 16031
rect 54076 16000 54125 16028
rect 54076 15988 54082 16000
rect 54113 15997 54125 16000
rect 54159 16028 54171 16031
rect 54389 16031 54447 16037
rect 54389 16028 54401 16031
rect 54159 16000 54401 16028
rect 54159 15997 54171 16000
rect 54113 15991 54171 15997
rect 54389 15997 54401 16000
rect 54435 15997 54447 16031
rect 55030 16028 55036 16040
rect 54389 15991 54447 15997
rect 54496 16000 55036 16028
rect 54496 15960 54524 16000
rect 55030 15988 55036 16000
rect 55088 16028 55094 16040
rect 56137 16031 56195 16037
rect 56137 16028 56149 16031
rect 55088 16000 56149 16028
rect 55088 15988 55094 16000
rect 56137 15997 56149 16000
rect 56183 15997 56195 16031
rect 56137 15991 56195 15997
rect 52013 15932 54524 15960
rect 50985 15923 51043 15929
rect 51629 15895 51687 15901
rect 51629 15892 51641 15895
rect 50080 15864 51641 15892
rect 51629 15861 51641 15864
rect 51675 15861 51687 15895
rect 51629 15855 51687 15861
rect 1104 15802 78844 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 78844 15802
rect 1104 15728 78844 15750
rect 8294 15648 8300 15700
rect 8352 15648 8358 15700
rect 11790 15648 11796 15700
rect 11848 15648 11854 15700
rect 14274 15648 14280 15700
rect 14332 15648 14338 15700
rect 16114 15648 16120 15700
rect 16172 15648 16178 15700
rect 19702 15688 19708 15700
rect 19306 15660 19708 15688
rect 15470 15620 15476 15632
rect 14752 15592 15476 15620
rect 12434 15512 12440 15564
rect 12492 15512 12498 15564
rect 13354 15512 13360 15564
rect 13412 15512 13418 15564
rect 14752 15561 14780 15592
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 14737 15555 14795 15561
rect 14737 15521 14749 15555
rect 14783 15521 14795 15555
rect 14737 15515 14795 15521
rect 14921 15555 14979 15561
rect 14921 15521 14933 15555
rect 14967 15552 14979 15555
rect 15010 15552 15016 15564
rect 14967 15524 15016 15552
rect 14967 15521 14979 15524
rect 14921 15515 14979 15521
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 15746 15512 15752 15564
rect 15804 15512 15810 15564
rect 19306 15552 19334 15660
rect 19702 15648 19708 15660
rect 19760 15648 19766 15700
rect 20533 15691 20591 15697
rect 20533 15657 20545 15691
rect 20579 15688 20591 15691
rect 24118 15688 24124 15700
rect 20579 15660 24124 15688
rect 20579 15657 20591 15660
rect 20533 15651 20591 15657
rect 24118 15648 24124 15660
rect 24176 15648 24182 15700
rect 25130 15648 25136 15700
rect 25188 15688 25194 15700
rect 25225 15691 25283 15697
rect 25225 15688 25237 15691
rect 25188 15660 25237 15688
rect 25188 15648 25194 15660
rect 25225 15657 25237 15660
rect 25271 15657 25283 15691
rect 25225 15651 25283 15657
rect 25685 15691 25743 15697
rect 25685 15657 25697 15691
rect 25731 15688 25743 15691
rect 27798 15688 27804 15700
rect 25731 15660 27804 15688
rect 25731 15657 25743 15660
rect 25685 15651 25743 15657
rect 27798 15648 27804 15660
rect 27856 15648 27862 15700
rect 27893 15691 27951 15697
rect 27893 15657 27905 15691
rect 27939 15688 27951 15691
rect 28994 15688 29000 15700
rect 27939 15660 29000 15688
rect 27939 15657 27951 15660
rect 27893 15651 27951 15657
rect 28994 15648 29000 15660
rect 29052 15648 29058 15700
rect 29641 15691 29699 15697
rect 29641 15657 29653 15691
rect 29687 15688 29699 15691
rect 31481 15691 31539 15697
rect 31481 15688 31493 15691
rect 29687 15660 31493 15688
rect 29687 15657 29699 15660
rect 29641 15651 29699 15657
rect 31481 15657 31493 15660
rect 31527 15688 31539 15691
rect 34333 15691 34391 15697
rect 34333 15688 34345 15691
rect 31527 15660 33456 15688
rect 31527 15657 31539 15660
rect 31481 15651 31539 15657
rect 19518 15580 19524 15632
rect 19576 15620 19582 15632
rect 19613 15623 19671 15629
rect 19613 15620 19625 15623
rect 19576 15592 19625 15620
rect 19576 15580 19582 15592
rect 19613 15589 19625 15592
rect 19659 15589 19671 15623
rect 19613 15583 19671 15589
rect 20073 15623 20131 15629
rect 20073 15589 20085 15623
rect 20119 15620 20131 15623
rect 22094 15620 22100 15632
rect 20119 15592 22100 15620
rect 20119 15589 20131 15592
rect 20073 15583 20131 15589
rect 22094 15580 22100 15592
rect 22152 15580 22158 15632
rect 24026 15620 24032 15632
rect 22664 15592 24032 15620
rect 18616 15524 19334 15552
rect 19797 15555 19855 15561
rect 18616 15496 18644 15524
rect 19797 15521 19809 15555
rect 19843 15521 19855 15555
rect 20441 15555 20499 15561
rect 20441 15552 20453 15555
rect 19797 15515 19855 15521
rect 20272 15524 20453 15552
rect 1394 15444 1400 15496
rect 1452 15484 1458 15496
rect 1673 15487 1731 15493
rect 1673 15484 1685 15487
rect 1452 15456 1685 15484
rect 1452 15444 1458 15456
rect 1673 15453 1685 15456
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 8110 15444 8116 15496
rect 8168 15444 8174 15496
rect 12158 15444 12164 15496
rect 12216 15444 12222 15496
rect 14642 15444 14648 15496
rect 14700 15484 14706 15496
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 14700 15456 15853 15484
rect 14700 15444 14706 15456
rect 15841 15453 15853 15456
rect 15887 15484 15899 15487
rect 18598 15484 18604 15496
rect 15887 15456 18604 15484
rect 15887 15453 15899 15456
rect 15841 15447 15899 15453
rect 18598 15444 18604 15456
rect 18656 15444 18662 15496
rect 18966 15444 18972 15496
rect 19024 15484 19030 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 19024 15456 19257 15484
rect 19024 15444 19030 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 19610 15444 19616 15496
rect 19668 15484 19674 15496
rect 19812 15484 19840 15515
rect 19668 15456 19840 15484
rect 19668 15444 19674 15456
rect 7926 15416 7932 15428
rect 1596 15388 7932 15416
rect 1596 15357 1624 15388
rect 7926 15376 7932 15388
rect 7984 15376 7990 15428
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15317 1639 15351
rect 1581 15311 1639 15317
rect 12253 15351 12311 15357
rect 12253 15317 12265 15351
rect 12299 15348 12311 15351
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 12299 15320 12817 15348
rect 12299 15317 12311 15320
rect 12253 15311 12311 15317
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 20272 15348 20300 15524
rect 20441 15521 20453 15524
rect 20487 15521 20499 15555
rect 20441 15515 20499 15521
rect 20533 15555 20591 15561
rect 20533 15521 20545 15555
rect 20579 15552 20591 15555
rect 20622 15552 20628 15564
rect 20579 15524 20628 15552
rect 20579 15521 20591 15524
rect 20533 15515 20591 15521
rect 20622 15512 20628 15524
rect 20680 15552 20686 15564
rect 20680 15524 20944 15552
rect 20680 15512 20686 15524
rect 20346 15444 20352 15496
rect 20404 15484 20410 15496
rect 20916 15493 20944 15524
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 22664 15552 22692 15592
rect 21508 15524 22692 15552
rect 21508 15512 21514 15524
rect 20901 15487 20959 15493
rect 20404 15456 20852 15484
rect 20404 15444 20410 15456
rect 20714 15376 20720 15428
rect 20772 15376 20778 15428
rect 20824 15416 20852 15456
rect 20901 15453 20913 15487
rect 20947 15453 20959 15487
rect 20901 15447 20959 15453
rect 21082 15444 21088 15496
rect 21140 15444 21146 15496
rect 21361 15487 21419 15493
rect 21361 15453 21373 15487
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15484 21695 15487
rect 22738 15484 22744 15496
rect 21683 15456 22744 15484
rect 21683 15453 21695 15456
rect 21637 15447 21695 15453
rect 21376 15416 21404 15447
rect 22738 15444 22744 15456
rect 22796 15444 22802 15496
rect 22848 15493 22876 15592
rect 24026 15580 24032 15592
rect 24084 15580 24090 15632
rect 24136 15552 24164 15648
rect 24762 15580 24768 15632
rect 24820 15620 24826 15632
rect 27982 15620 27988 15632
rect 24820 15592 27988 15620
rect 24820 15580 24826 15592
rect 27982 15580 27988 15592
rect 28040 15580 28046 15632
rect 28629 15623 28687 15629
rect 28629 15589 28641 15623
rect 28675 15589 28687 15623
rect 28629 15583 28687 15589
rect 25314 15552 25320 15564
rect 24136 15524 25320 15552
rect 25314 15512 25320 15524
rect 25372 15512 25378 15564
rect 25866 15512 25872 15564
rect 25924 15552 25930 15564
rect 26142 15552 26148 15564
rect 25924 15524 26148 15552
rect 25924 15512 25930 15524
rect 26142 15512 26148 15524
rect 26200 15552 26206 15564
rect 26200 15524 26832 15552
rect 26200 15512 26206 15524
rect 22833 15487 22891 15493
rect 22833 15453 22845 15487
rect 22879 15453 22891 15487
rect 22833 15447 22891 15453
rect 23014 15444 23020 15496
rect 23072 15444 23078 15496
rect 23198 15444 23204 15496
rect 23256 15444 23262 15496
rect 25222 15444 25228 15496
rect 25280 15444 25286 15496
rect 25498 15444 25504 15496
rect 25556 15444 25562 15496
rect 25958 15444 25964 15496
rect 26016 15484 26022 15496
rect 26053 15487 26111 15493
rect 26053 15484 26065 15487
rect 26016 15456 26065 15484
rect 26016 15444 26022 15456
rect 26053 15453 26065 15456
rect 26099 15453 26111 15487
rect 26053 15447 26111 15453
rect 26418 15444 26424 15496
rect 26476 15444 26482 15496
rect 26804 15493 26832 15524
rect 27430 15512 27436 15564
rect 27488 15552 27494 15564
rect 28644 15552 28672 15583
rect 29656 15552 29684 15651
rect 27488 15524 28396 15552
rect 28644 15524 29040 15552
rect 27488 15512 27494 15524
rect 26789 15487 26847 15493
rect 26789 15453 26801 15487
rect 26835 15453 26847 15487
rect 26789 15447 26847 15453
rect 27246 15444 27252 15496
rect 27304 15444 27310 15496
rect 27706 15444 27712 15496
rect 27764 15444 27770 15496
rect 28368 15493 28396 15524
rect 28353 15487 28411 15493
rect 28353 15453 28365 15487
rect 28399 15453 28411 15487
rect 28353 15447 28411 15453
rect 28810 15444 28816 15496
rect 28868 15444 28874 15496
rect 29012 15493 29040 15524
rect 29104 15524 29684 15552
rect 29104 15493 29132 15524
rect 28997 15487 29055 15493
rect 28997 15453 29009 15487
rect 29043 15453 29055 15487
rect 28997 15447 29055 15453
rect 29089 15487 29147 15493
rect 29089 15453 29101 15487
rect 29135 15453 29147 15487
rect 29089 15447 29147 15453
rect 29181 15487 29239 15493
rect 29181 15453 29193 15487
rect 29227 15484 29239 15487
rect 29546 15484 29552 15496
rect 29227 15456 29552 15484
rect 29227 15453 29239 15456
rect 29181 15447 29239 15453
rect 22922 15416 22928 15428
rect 20824 15388 21404 15416
rect 21082 15348 21088 15360
rect 20272 15320 21088 15348
rect 12805 15311 12863 15317
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 21376 15348 21404 15388
rect 22066 15388 22928 15416
rect 22066 15348 22094 15388
rect 22922 15376 22928 15388
rect 22980 15376 22986 15428
rect 25240 15416 25268 15444
rect 27062 15416 27068 15428
rect 25240 15388 27068 15416
rect 27062 15376 27068 15388
rect 27120 15376 27126 15428
rect 27522 15376 27528 15428
rect 27580 15416 27586 15428
rect 28445 15419 28503 15425
rect 28445 15416 28457 15419
rect 27580 15388 28457 15416
rect 27580 15376 27586 15388
rect 28445 15385 28457 15388
rect 28491 15385 28503 15419
rect 28445 15379 28503 15385
rect 28629 15419 28687 15425
rect 28629 15385 28641 15419
rect 28675 15416 28687 15419
rect 29196 15416 29224 15447
rect 29546 15444 29552 15456
rect 29604 15444 29610 15496
rect 29730 15444 29736 15496
rect 29788 15444 29794 15496
rect 31110 15444 31116 15496
rect 31168 15444 31174 15496
rect 30009 15419 30067 15425
rect 30009 15416 30021 15419
rect 28675 15388 29224 15416
rect 29380 15388 30021 15416
rect 28675 15385 28687 15388
rect 28629 15379 28687 15385
rect 21376 15320 22094 15348
rect 22462 15308 22468 15360
rect 22520 15348 22526 15360
rect 22649 15351 22707 15357
rect 22649 15348 22661 15351
rect 22520 15320 22661 15348
rect 22520 15308 22526 15320
rect 22649 15317 22661 15320
rect 22695 15317 22707 15351
rect 22649 15311 22707 15317
rect 23109 15351 23167 15357
rect 23109 15317 23121 15351
rect 23155 15348 23167 15351
rect 23934 15348 23940 15360
rect 23155 15320 23940 15348
rect 23155 15317 23167 15320
rect 23109 15311 23167 15317
rect 23934 15308 23940 15320
rect 23992 15348 23998 15360
rect 25498 15348 25504 15360
rect 23992 15320 25504 15348
rect 23992 15308 23998 15320
rect 25498 15308 25504 15320
rect 25556 15308 25562 15360
rect 26970 15308 26976 15360
rect 27028 15348 27034 15360
rect 28644 15348 28672 15379
rect 29380 15357 29408 15388
rect 30009 15385 30021 15388
rect 30055 15385 30067 15419
rect 30009 15379 30067 15385
rect 31570 15376 31576 15428
rect 31628 15416 31634 15428
rect 32677 15419 32735 15425
rect 32677 15416 32689 15419
rect 31628 15388 32689 15416
rect 31628 15376 31634 15388
rect 32677 15385 32689 15388
rect 32723 15416 32735 15419
rect 33226 15416 33232 15428
rect 32723 15388 33232 15416
rect 32723 15385 32735 15388
rect 32677 15379 32735 15385
rect 33226 15376 33232 15388
rect 33284 15376 33290 15428
rect 33428 15416 33456 15660
rect 33520 15660 34345 15688
rect 33520 15493 33548 15660
rect 34333 15657 34345 15660
rect 34379 15688 34391 15691
rect 38746 15688 38752 15700
rect 34379 15660 38752 15688
rect 34379 15657 34391 15660
rect 34333 15651 34391 15657
rect 38746 15648 38752 15660
rect 38804 15688 38810 15700
rect 40586 15688 40592 15700
rect 38804 15660 40592 15688
rect 38804 15648 38810 15660
rect 40586 15648 40592 15660
rect 40644 15648 40650 15700
rect 41414 15648 41420 15700
rect 41472 15688 41478 15700
rect 42610 15688 42616 15700
rect 41472 15660 42616 15688
rect 41472 15648 41478 15660
rect 42610 15648 42616 15660
rect 42668 15648 42674 15700
rect 45922 15648 45928 15700
rect 45980 15688 45986 15700
rect 46750 15688 46756 15700
rect 45980 15660 46756 15688
rect 45980 15648 45986 15660
rect 46750 15648 46756 15660
rect 46808 15648 46814 15700
rect 49878 15648 49884 15700
rect 49936 15648 49942 15700
rect 50709 15691 50767 15697
rect 50709 15657 50721 15691
rect 50755 15688 50767 15691
rect 51166 15688 51172 15700
rect 50755 15660 51172 15688
rect 50755 15657 50767 15660
rect 50709 15651 50767 15657
rect 51166 15648 51172 15660
rect 51224 15648 51230 15700
rect 53285 15691 53343 15697
rect 53285 15657 53297 15691
rect 53331 15688 53343 15691
rect 53374 15688 53380 15700
rect 53331 15660 53380 15688
rect 53331 15657 53343 15660
rect 53285 15651 53343 15657
rect 53374 15648 53380 15660
rect 53432 15648 53438 15700
rect 34422 15580 34428 15632
rect 34480 15620 34486 15632
rect 35986 15620 35992 15632
rect 34480 15592 35992 15620
rect 34480 15580 34486 15592
rect 35986 15580 35992 15592
rect 36044 15620 36050 15632
rect 37366 15620 37372 15632
rect 36044 15592 37372 15620
rect 36044 15580 36050 15592
rect 35434 15512 35440 15564
rect 35492 15512 35498 15564
rect 33505 15487 33563 15493
rect 33505 15453 33517 15487
rect 33551 15453 33563 15487
rect 33505 15447 33563 15453
rect 33686 15444 33692 15496
rect 33744 15484 33750 15496
rect 33873 15487 33931 15493
rect 33873 15484 33885 15487
rect 33744 15456 33885 15484
rect 33744 15444 33750 15456
rect 33873 15453 33885 15456
rect 33919 15453 33931 15487
rect 33873 15447 33931 15453
rect 34057 15487 34115 15493
rect 34057 15453 34069 15487
rect 34103 15453 34115 15487
rect 34057 15447 34115 15453
rect 34149 15487 34207 15493
rect 34149 15453 34161 15487
rect 34195 15484 34207 15487
rect 34701 15487 34759 15493
rect 34701 15484 34713 15487
rect 34195 15456 34713 15484
rect 34195 15453 34207 15456
rect 34149 15447 34207 15453
rect 34701 15453 34713 15456
rect 34747 15453 34759 15487
rect 34701 15447 34759 15453
rect 34072 15416 34100 15447
rect 34790 15444 34796 15496
rect 34848 15484 34854 15496
rect 35253 15487 35311 15493
rect 35253 15484 35265 15487
rect 34848 15456 35265 15484
rect 34848 15444 34854 15456
rect 35253 15453 35265 15456
rect 35299 15453 35311 15487
rect 35253 15447 35311 15453
rect 35342 15444 35348 15496
rect 35400 15484 35406 15496
rect 35621 15487 35679 15493
rect 35621 15484 35633 15487
rect 35400 15456 35633 15484
rect 35400 15444 35406 15456
rect 35621 15453 35633 15456
rect 35667 15453 35679 15487
rect 35621 15447 35679 15453
rect 35805 15487 35863 15493
rect 35805 15453 35817 15487
rect 35851 15453 35863 15487
rect 35805 15447 35863 15453
rect 35897 15487 35955 15493
rect 35897 15453 35909 15487
rect 35943 15484 35955 15487
rect 36541 15487 36599 15493
rect 36541 15484 36553 15487
rect 35943 15456 36553 15484
rect 35943 15453 35955 15456
rect 35897 15447 35955 15453
rect 36541 15453 36553 15456
rect 36587 15453 36599 15487
rect 36541 15447 36599 15453
rect 34238 15416 34244 15428
rect 33428 15388 33824 15416
rect 34072 15388 34244 15416
rect 27028 15320 28672 15348
rect 29365 15351 29423 15357
rect 27028 15308 27034 15320
rect 29365 15317 29377 15351
rect 29411 15317 29423 15351
rect 29365 15311 29423 15317
rect 33502 15308 33508 15360
rect 33560 15348 33566 15360
rect 33689 15351 33747 15357
rect 33689 15348 33701 15351
rect 33560 15320 33701 15348
rect 33560 15308 33566 15320
rect 33689 15317 33701 15320
rect 33735 15317 33747 15351
rect 33796 15348 33824 15388
rect 34238 15376 34244 15388
rect 34296 15376 34302 15428
rect 34330 15376 34336 15428
rect 34388 15416 34394 15428
rect 35820 15416 35848 15447
rect 35989 15419 36047 15425
rect 35989 15416 36001 15419
rect 34388 15388 36001 15416
rect 34388 15376 34394 15388
rect 35989 15385 36001 15388
rect 36035 15385 36047 15419
rect 35989 15379 36047 15385
rect 36357 15419 36415 15425
rect 36357 15385 36369 15419
rect 36403 15416 36415 15419
rect 36648 15416 36676 15592
rect 37366 15580 37372 15592
rect 37424 15620 37430 15632
rect 37424 15592 38056 15620
rect 37424 15580 37430 15592
rect 36998 15444 37004 15496
rect 37056 15484 37062 15496
rect 37093 15487 37151 15493
rect 37093 15484 37105 15487
rect 37056 15456 37105 15484
rect 37056 15444 37062 15456
rect 37093 15453 37105 15456
rect 37139 15453 37151 15487
rect 37093 15447 37151 15453
rect 37200 15456 37872 15484
rect 36403 15388 36676 15416
rect 36403 15385 36415 15388
rect 36357 15379 36415 15385
rect 37200 15348 37228 15456
rect 37274 15376 37280 15428
rect 37332 15416 37338 15428
rect 37369 15419 37427 15425
rect 37369 15416 37381 15419
rect 37332 15388 37381 15416
rect 37332 15376 37338 15388
rect 37369 15385 37381 15388
rect 37415 15385 37427 15419
rect 37369 15379 37427 15385
rect 37553 15419 37611 15425
rect 37553 15385 37565 15419
rect 37599 15416 37611 15419
rect 37642 15416 37648 15428
rect 37599 15388 37648 15416
rect 37599 15385 37611 15388
rect 37553 15379 37611 15385
rect 37642 15376 37648 15388
rect 37700 15376 37706 15428
rect 33796 15320 37228 15348
rect 33689 15311 33747 15317
rect 37734 15308 37740 15360
rect 37792 15308 37798 15360
rect 37844 15348 37872 15456
rect 37918 15444 37924 15496
rect 37976 15444 37982 15496
rect 38028 15416 38056 15592
rect 49602 15580 49608 15632
rect 49660 15620 49666 15632
rect 50890 15620 50896 15632
rect 49660 15592 50896 15620
rect 49660 15580 49666 15592
rect 50890 15580 50896 15592
rect 50948 15580 50954 15632
rect 56137 15623 56195 15629
rect 56137 15589 56149 15623
rect 56183 15589 56195 15623
rect 56137 15583 56195 15589
rect 38105 15555 38163 15561
rect 38105 15521 38117 15555
rect 38151 15552 38163 15555
rect 38562 15552 38568 15564
rect 38151 15524 38568 15552
rect 38151 15521 38163 15524
rect 38105 15515 38163 15521
rect 38562 15512 38568 15524
rect 38620 15512 38626 15564
rect 39853 15555 39911 15561
rect 39853 15521 39865 15555
rect 39899 15552 39911 15555
rect 40862 15552 40868 15564
rect 39899 15524 40868 15552
rect 39899 15521 39911 15524
rect 39853 15515 39911 15521
rect 40862 15512 40868 15524
rect 40920 15552 40926 15564
rect 40920 15524 41414 15552
rect 40920 15512 40926 15524
rect 38197 15487 38255 15493
rect 38197 15453 38209 15487
rect 38243 15484 38255 15487
rect 38841 15487 38899 15493
rect 38841 15484 38853 15487
rect 38243 15456 38853 15484
rect 38243 15453 38255 15456
rect 38197 15447 38255 15453
rect 38841 15453 38853 15456
rect 38887 15453 38899 15487
rect 38841 15447 38899 15453
rect 39298 15444 39304 15496
rect 39356 15484 39362 15496
rect 39393 15487 39451 15493
rect 39393 15484 39405 15487
rect 39356 15456 39405 15484
rect 39356 15444 39362 15456
rect 39393 15453 39405 15456
rect 39439 15453 39451 15487
rect 41386 15484 41414 15524
rect 45738 15512 45744 15564
rect 45796 15552 45802 15564
rect 46569 15555 46627 15561
rect 46569 15552 46581 15555
rect 45796 15524 46581 15552
rect 45796 15512 45802 15524
rect 46569 15521 46581 15524
rect 46615 15552 46627 15555
rect 46842 15552 46848 15564
rect 46615 15524 46848 15552
rect 46615 15521 46627 15524
rect 46569 15515 46627 15521
rect 46842 15512 46848 15524
rect 46900 15512 46906 15564
rect 49878 15512 49884 15564
rect 49936 15552 49942 15564
rect 52270 15552 52276 15564
rect 49936 15524 50384 15552
rect 49936 15512 49942 15524
rect 41877 15487 41935 15493
rect 41877 15484 41889 15487
rect 41386 15456 41889 15484
rect 39393 15447 39451 15453
rect 41877 15453 41889 15456
rect 41923 15453 41935 15487
rect 41877 15447 41935 15453
rect 43530 15444 43536 15496
rect 43588 15484 43594 15496
rect 44269 15487 44327 15493
rect 44269 15484 44281 15487
rect 43588 15456 44281 15484
rect 43588 15444 43594 15456
rect 44269 15453 44281 15456
rect 44315 15453 44327 15487
rect 44269 15447 44327 15453
rect 48130 15444 48136 15496
rect 48188 15484 48194 15496
rect 50356 15493 50384 15524
rect 50448 15524 52276 15552
rect 50448 15493 50476 15524
rect 52270 15512 52276 15524
rect 52328 15552 52334 15564
rect 54938 15552 54944 15564
rect 52328 15524 54944 15552
rect 52328 15512 52334 15524
rect 54938 15512 54944 15524
rect 54996 15552 55002 15564
rect 54996 15524 55720 15552
rect 54996 15512 55002 15524
rect 49697 15487 49755 15493
rect 49697 15484 49709 15487
rect 48188 15456 49709 15484
rect 48188 15444 48194 15456
rect 49697 15453 49709 15456
rect 49743 15484 49755 15487
rect 50157 15487 50215 15493
rect 50157 15484 50169 15487
rect 49743 15456 50169 15484
rect 49743 15453 49755 15456
rect 49697 15447 49755 15453
rect 50157 15453 50169 15456
rect 50203 15453 50215 15487
rect 50157 15447 50215 15453
rect 50341 15487 50399 15493
rect 50341 15453 50353 15487
rect 50387 15453 50399 15487
rect 50341 15447 50399 15453
rect 50433 15487 50491 15493
rect 50433 15453 50445 15487
rect 50479 15453 50491 15487
rect 50433 15447 50491 15453
rect 50525 15487 50583 15493
rect 50525 15453 50537 15487
rect 50571 15484 50583 15487
rect 50890 15484 50896 15496
rect 50571 15456 50896 15484
rect 50571 15453 50583 15456
rect 50525 15447 50583 15453
rect 50890 15444 50896 15456
rect 50948 15444 50954 15496
rect 54202 15444 54208 15496
rect 54260 15484 54266 15496
rect 54297 15487 54355 15493
rect 54297 15484 54309 15487
rect 54260 15456 54309 15484
rect 54260 15444 54266 15456
rect 54297 15453 54309 15456
rect 54343 15453 54355 15487
rect 54573 15487 54631 15493
rect 54573 15484 54585 15487
rect 54297 15447 54355 15453
rect 54404 15456 54585 15484
rect 38381 15419 38439 15425
rect 38381 15416 38393 15419
rect 38028 15388 38393 15416
rect 38381 15385 38393 15388
rect 38427 15416 38439 15419
rect 38749 15419 38807 15425
rect 38749 15416 38761 15419
rect 38427 15388 38761 15416
rect 38427 15385 38439 15388
rect 38381 15379 38439 15385
rect 38749 15385 38761 15388
rect 38795 15416 38807 15419
rect 40034 15416 40040 15428
rect 38795 15388 40040 15416
rect 38795 15385 38807 15388
rect 38749 15379 38807 15385
rect 40034 15376 40040 15388
rect 40092 15376 40098 15428
rect 40126 15376 40132 15428
rect 40184 15376 40190 15428
rect 41414 15416 41420 15428
rect 41354 15388 41420 15416
rect 41414 15376 41420 15388
rect 41472 15376 41478 15428
rect 41525 15388 42104 15416
rect 41525 15348 41553 15388
rect 37844 15320 41553 15348
rect 41598 15308 41604 15360
rect 41656 15308 41662 15360
rect 42076 15348 42104 15388
rect 42150 15376 42156 15428
rect 42208 15376 42214 15428
rect 42610 15376 42616 15428
rect 42668 15376 42674 15428
rect 45649 15419 45707 15425
rect 45649 15385 45661 15419
rect 45695 15416 45707 15419
rect 45741 15419 45799 15425
rect 45741 15416 45753 15419
rect 45695 15388 45753 15416
rect 45695 15385 45707 15388
rect 45649 15379 45707 15385
rect 45741 15385 45753 15388
rect 45787 15416 45799 15419
rect 45830 15416 45836 15428
rect 45787 15388 45836 15416
rect 45787 15385 45799 15388
rect 45741 15379 45799 15385
rect 45830 15376 45836 15388
rect 45888 15376 45894 15428
rect 48958 15376 48964 15428
rect 49016 15416 49022 15428
rect 50982 15416 50988 15428
rect 49016 15388 50988 15416
rect 49016 15376 49022 15388
rect 50982 15376 50988 15388
rect 51040 15416 51046 15428
rect 53834 15416 53840 15428
rect 51040 15388 53840 15416
rect 51040 15376 51046 15388
rect 53834 15376 53840 15388
rect 53892 15416 53898 15428
rect 54404 15416 54432 15456
rect 54573 15453 54585 15456
rect 54619 15453 54631 15487
rect 54573 15447 54631 15453
rect 54662 15444 54668 15496
rect 54720 15444 54726 15496
rect 55490 15444 55496 15496
rect 55548 15444 55554 15496
rect 55585 15487 55643 15493
rect 55585 15453 55597 15487
rect 55631 15453 55643 15487
rect 55692 15484 55720 15524
rect 55766 15512 55772 15564
rect 55824 15552 55830 15564
rect 56152 15552 56180 15583
rect 55824 15524 56180 15552
rect 55824 15512 55830 15524
rect 55861 15487 55919 15493
rect 55861 15484 55873 15487
rect 55692 15456 55873 15484
rect 55585 15447 55643 15453
rect 55861 15453 55873 15456
rect 55907 15453 55919 15487
rect 55861 15447 55919 15453
rect 53892 15388 54432 15416
rect 53892 15376 53898 15388
rect 54478 15376 54484 15428
rect 54536 15376 54542 15428
rect 55600 15416 55628 15447
rect 54864 15388 55628 15416
rect 55876 15416 55904 15447
rect 55950 15444 55956 15496
rect 56008 15444 56014 15496
rect 56502 15416 56508 15428
rect 55876 15388 56508 15416
rect 43438 15348 43444 15360
rect 42076 15320 43444 15348
rect 43438 15308 43444 15320
rect 43496 15308 43502 15360
rect 43530 15308 43536 15360
rect 43588 15348 43594 15360
rect 43625 15351 43683 15357
rect 43625 15348 43637 15351
rect 43588 15320 43637 15348
rect 43588 15308 43594 15320
rect 43625 15317 43637 15320
rect 43671 15317 43683 15351
rect 43625 15311 43683 15317
rect 43714 15308 43720 15360
rect 43772 15308 43778 15360
rect 45462 15308 45468 15360
rect 45520 15348 45526 15360
rect 46753 15351 46811 15357
rect 46753 15348 46765 15351
rect 45520 15320 46765 15348
rect 45520 15308 45526 15320
rect 46753 15317 46765 15320
rect 46799 15348 46811 15351
rect 47486 15348 47492 15360
rect 46799 15320 47492 15348
rect 46799 15317 46811 15320
rect 46753 15311 46811 15317
rect 47486 15308 47492 15320
rect 47544 15308 47550 15360
rect 48590 15308 48596 15360
rect 48648 15348 48654 15360
rect 49970 15348 49976 15360
rect 48648 15320 49976 15348
rect 48648 15308 48654 15320
rect 49970 15308 49976 15320
rect 50028 15308 50034 15360
rect 50890 15308 50896 15360
rect 50948 15308 50954 15360
rect 54864 15357 54892 15388
rect 56502 15376 56508 15388
rect 56560 15376 56566 15428
rect 54849 15351 54907 15357
rect 54849 15317 54861 15351
rect 54895 15317 54907 15351
rect 54849 15311 54907 15317
rect 55214 15308 55220 15360
rect 55272 15348 55278 15360
rect 55309 15351 55367 15357
rect 55309 15348 55321 15351
rect 55272 15320 55321 15348
rect 55272 15308 55278 15320
rect 55309 15317 55321 15320
rect 55355 15317 55367 15351
rect 55309 15311 55367 15317
rect 1104 15258 78844 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 66314 15258
rect 66366 15206 66378 15258
rect 66430 15206 66442 15258
rect 66494 15206 66506 15258
rect 66558 15206 66570 15258
rect 66622 15206 78844 15258
rect 1104 15184 78844 15206
rect 8110 15144 8116 15156
rect 7852 15116 8116 15144
rect 7561 15011 7619 15017
rect 7561 14977 7573 15011
rect 7607 15008 7619 15011
rect 7650 15008 7656 15020
rect 7607 14980 7656 15008
rect 7607 14977 7619 14980
rect 7561 14971 7619 14977
rect 7650 14968 7656 14980
rect 7708 14968 7714 15020
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 15008 7803 15011
rect 7852 15008 7880 15116
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 17126 15104 17132 15156
rect 17184 15144 17190 15156
rect 17221 15147 17279 15153
rect 17221 15144 17233 15147
rect 17184 15116 17233 15144
rect 17184 15104 17190 15116
rect 17221 15113 17233 15116
rect 17267 15113 17279 15147
rect 17221 15107 17279 15113
rect 25685 15147 25743 15153
rect 25685 15113 25697 15147
rect 25731 15113 25743 15147
rect 25685 15107 25743 15113
rect 26329 15147 26387 15153
rect 26329 15113 26341 15147
rect 26375 15144 26387 15147
rect 26418 15144 26424 15156
rect 26375 15116 26424 15144
rect 26375 15113 26387 15116
rect 26329 15107 26387 15113
rect 9766 15076 9772 15088
rect 7944 15048 8800 15076
rect 7944 15020 7972 15048
rect 7791 14980 7880 15008
rect 7791 14977 7803 14980
rect 7745 14971 7803 14977
rect 7926 14968 7932 15020
rect 7984 14968 7990 15020
rect 8205 15011 8263 15017
rect 8205 14977 8217 15011
rect 8251 15008 8263 15011
rect 8570 15008 8576 15020
rect 8251 14980 8576 15008
rect 8251 14977 8263 14980
rect 8205 14971 8263 14977
rect 8570 14968 8576 14980
rect 8628 14968 8634 15020
rect 8772 15017 8800 15048
rect 8864 15048 9772 15076
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 14977 8815 15011
rect 8757 14971 8815 14977
rect 8297 14943 8355 14949
rect 8297 14909 8309 14943
rect 8343 14940 8355 14943
rect 8864 14940 8892 15048
rect 9766 15036 9772 15048
rect 9824 15036 9830 15088
rect 19521 15079 19579 15085
rect 19521 15045 19533 15079
rect 19567 15076 19579 15079
rect 20346 15076 20352 15088
rect 19567 15048 20352 15076
rect 19567 15045 19579 15048
rect 19521 15039 19579 15045
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 20533 15079 20591 15085
rect 20533 15045 20545 15079
rect 20579 15076 20591 15079
rect 20622 15076 20628 15088
rect 20579 15048 20628 15076
rect 20579 15045 20591 15048
rect 20533 15039 20591 15045
rect 20622 15036 20628 15048
rect 20680 15076 20686 15088
rect 23014 15076 23020 15088
rect 20680 15048 22094 15076
rect 20680 15036 20686 15048
rect 9490 14968 9496 15020
rect 9548 14968 9554 15020
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 12250 15008 12256 15020
rect 10928 14980 12256 15008
rect 10928 14968 10934 14980
rect 12250 14968 12256 14980
rect 12308 14968 12314 15020
rect 12342 14968 12348 15020
rect 12400 15008 12406 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12400 14980 13001 15008
rect 12400 14968 12406 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 9769 14943 9827 14949
rect 9769 14940 9781 14943
rect 8343 14912 8892 14940
rect 8956 14912 9781 14940
rect 8343 14909 8355 14912
rect 8297 14903 8355 14909
rect 8956 14881 8984 14912
rect 9769 14909 9781 14912
rect 9815 14909 9827 14943
rect 9769 14903 9827 14909
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14940 11299 14943
rect 12360 14940 12388 14968
rect 11287 14912 12388 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 8941 14875 8999 14881
rect 8941 14841 8953 14875
rect 8987 14841 8999 14875
rect 13004 14872 13032 14971
rect 16850 14968 16856 15020
rect 16908 15008 16914 15020
rect 16908 14980 17724 15008
rect 16908 14968 16914 14980
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14940 13139 14943
rect 13446 14940 13452 14952
rect 13127 14912 13452 14940
rect 13127 14909 13139 14912
rect 13081 14903 13139 14909
rect 13446 14900 13452 14912
rect 13504 14900 13510 14952
rect 16942 14900 16948 14952
rect 17000 14900 17006 14952
rect 17696 14940 17724 14980
rect 18598 14968 18604 15020
rect 18656 14968 18662 15020
rect 22066 15008 22094 15048
rect 22480 15048 23020 15076
rect 22480 15017 22508 15048
rect 23014 15036 23020 15048
rect 23072 15076 23078 15088
rect 23072 15048 23244 15076
rect 23072 15036 23078 15048
rect 22465 15011 22523 15017
rect 22465 15008 22477 15011
rect 22066 14980 22477 15008
rect 22465 14977 22477 14980
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 22649 15011 22707 15017
rect 22649 14977 22661 15011
rect 22695 15008 22707 15011
rect 22738 15008 22744 15020
rect 22695 14980 22744 15008
rect 22695 14977 22707 14980
rect 22649 14971 22707 14977
rect 22738 14968 22744 14980
rect 22796 14968 22802 15020
rect 22922 14968 22928 15020
rect 22980 14968 22986 15020
rect 23216 15017 23244 15048
rect 24026 15036 24032 15088
rect 24084 15076 24090 15088
rect 24121 15079 24179 15085
rect 24121 15076 24133 15079
rect 24084 15048 24133 15076
rect 24084 15036 24090 15048
rect 24121 15045 24133 15048
rect 24167 15045 24179 15079
rect 25700 15076 25728 15107
rect 26418 15104 26424 15116
rect 26476 15104 26482 15156
rect 28902 15104 28908 15156
rect 28960 15144 28966 15156
rect 28997 15147 29055 15153
rect 28997 15144 29009 15147
rect 28960 15116 29009 15144
rect 28960 15104 28966 15116
rect 28997 15113 29009 15116
rect 29043 15113 29055 15147
rect 28997 15107 29055 15113
rect 33226 15104 33232 15156
rect 33284 15144 33290 15156
rect 33284 15116 37596 15144
rect 33284 15104 33290 15116
rect 27341 15079 27399 15085
rect 27341 15076 27353 15079
rect 25700 15048 27353 15076
rect 24121 15039 24179 15045
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 14977 23167 15011
rect 23109 14971 23167 14977
rect 23201 15011 23259 15017
rect 23201 14977 23213 15011
rect 23247 14977 23259 15011
rect 23201 14971 23259 14977
rect 23385 15011 23443 15017
rect 23385 14977 23397 15011
rect 23431 15008 23443 15011
rect 23937 15011 23995 15017
rect 23937 15008 23949 15011
rect 23431 14980 23949 15008
rect 23431 14977 23443 14980
rect 23385 14971 23443 14977
rect 23937 14977 23949 14980
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 19153 14943 19211 14949
rect 19153 14940 19165 14943
rect 17696 14912 19165 14940
rect 19153 14909 19165 14912
rect 19199 14940 19211 14943
rect 19610 14940 19616 14952
rect 19199 14912 19616 14940
rect 19199 14909 19211 14912
rect 19153 14903 19211 14909
rect 19610 14900 19616 14912
rect 19668 14900 19674 14952
rect 19702 14900 19708 14952
rect 19760 14940 19766 14952
rect 20165 14943 20223 14949
rect 20165 14940 20177 14943
rect 19760 14912 20177 14940
rect 19760 14900 19766 14912
rect 20165 14909 20177 14912
rect 20211 14909 20223 14943
rect 23124 14940 23152 14971
rect 23400 14940 23428 14971
rect 25314 14968 25320 15020
rect 25372 14968 25378 15020
rect 25498 14968 25504 15020
rect 25556 14968 25562 15020
rect 26252 15017 26280 15048
rect 27341 15045 27353 15048
rect 27387 15045 27399 15079
rect 27341 15039 27399 15045
rect 27433 15079 27491 15085
rect 27433 15045 27445 15079
rect 27479 15076 27491 15079
rect 31478 15076 31484 15088
rect 27479 15048 31484 15076
rect 27479 15045 27491 15048
rect 27433 15039 27491 15045
rect 31478 15036 31484 15048
rect 31536 15036 31542 15088
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 14977 26295 15011
rect 26415 15011 26473 15017
rect 26415 15008 26427 15011
rect 26237 14971 26295 14977
rect 26344 14980 26427 15008
rect 26344 14940 26372 14980
rect 26415 14977 26427 14980
rect 26461 15008 26473 15011
rect 26970 15008 26976 15020
rect 26461 14980 26976 15008
rect 26461 14977 26473 14980
rect 26415 14971 26473 14977
rect 26970 14968 26976 14980
rect 27028 14968 27034 15020
rect 27062 14968 27068 15020
rect 27120 14968 27126 15020
rect 27154 14968 27160 15020
rect 27212 14968 27218 15020
rect 27571 15011 27629 15017
rect 27571 14977 27583 15011
rect 27617 15008 27629 15011
rect 27706 15008 27712 15020
rect 27617 14980 27712 15008
rect 27617 14977 27629 14980
rect 27571 14971 27629 14977
rect 27706 14968 27712 14980
rect 27764 15008 27770 15020
rect 28350 15008 28356 15020
rect 27764 14980 28356 15008
rect 27764 14968 27770 14980
rect 28350 14968 28356 14980
rect 28408 14968 28414 15020
rect 28626 14968 28632 15020
rect 28684 14968 28690 15020
rect 28718 14968 28724 15020
rect 28776 15008 28782 15020
rect 28905 15011 28963 15017
rect 28905 15008 28917 15011
rect 28776 14980 28917 15008
rect 28776 14968 28782 14980
rect 28905 14977 28917 14980
rect 28951 14977 28963 15011
rect 28905 14971 28963 14977
rect 29089 15011 29147 15017
rect 29089 14977 29101 15011
rect 29135 15008 29147 15011
rect 29178 15008 29184 15020
rect 29135 14980 29184 15008
rect 29135 14977 29147 14980
rect 29089 14971 29147 14977
rect 29178 14968 29184 14980
rect 29236 14968 29242 15020
rect 32214 14968 32220 15020
rect 32272 15008 32278 15020
rect 33134 15008 33140 15020
rect 32272 14980 33140 15008
rect 32272 14968 32278 14980
rect 33134 14968 33140 14980
rect 33192 14968 33198 15020
rect 33226 14968 33232 15020
rect 33284 14968 33290 15020
rect 35268 15017 35296 15116
rect 35434 15036 35440 15088
rect 35492 15076 35498 15088
rect 35529 15079 35587 15085
rect 35529 15076 35541 15079
rect 35492 15048 35541 15076
rect 35492 15036 35498 15048
rect 35529 15045 35541 15048
rect 35575 15045 35587 15079
rect 35529 15039 35587 15045
rect 37568 15017 37596 15116
rect 37642 15104 37648 15156
rect 37700 15144 37706 15156
rect 37700 15116 39993 15144
rect 37700 15104 37706 15116
rect 37734 15036 37740 15088
rect 37792 15076 37798 15088
rect 37829 15079 37887 15085
rect 37829 15076 37841 15079
rect 37792 15048 37841 15076
rect 37792 15036 37798 15048
rect 37829 15045 37841 15048
rect 37875 15045 37887 15079
rect 39114 15076 39120 15088
rect 39054 15048 39120 15076
rect 37829 15039 37887 15045
rect 39114 15036 39120 15048
rect 39172 15076 39178 15088
rect 39390 15076 39396 15088
rect 39172 15048 39396 15076
rect 39172 15036 39178 15048
rect 39390 15036 39396 15048
rect 39448 15036 39454 15088
rect 35253 15011 35311 15017
rect 34638 14980 34744 15008
rect 20165 14903 20223 14909
rect 22066 14912 23428 14940
rect 24228 14912 26372 14940
rect 13004 14844 17264 14872
rect 8941 14835 8999 14841
rect 13265 14807 13323 14813
rect 13265 14773 13277 14807
rect 13311 14804 13323 14807
rect 14274 14804 14280 14816
rect 13311 14776 14280 14804
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 17236 14804 17264 14844
rect 18984 14844 19196 14872
rect 18984 14816 19012 14844
rect 18966 14804 18972 14816
rect 17236 14776 18972 14804
rect 18966 14764 18972 14776
rect 19024 14764 19030 14816
rect 19058 14764 19064 14816
rect 19116 14764 19122 14816
rect 19168 14804 19196 14844
rect 19242 14832 19248 14884
rect 19300 14872 19306 14884
rect 19518 14872 19524 14884
rect 19300 14844 19524 14872
rect 19300 14832 19306 14844
rect 19518 14832 19524 14844
rect 19576 14872 19582 14884
rect 20073 14875 20131 14881
rect 20073 14872 20085 14875
rect 19576 14844 20085 14872
rect 19576 14832 19582 14844
rect 20073 14841 20085 14844
rect 20119 14841 20131 14875
rect 20073 14835 20131 14841
rect 21082 14832 21088 14884
rect 21140 14872 21146 14884
rect 22066 14872 22094 14912
rect 21140 14844 22094 14872
rect 21140 14832 21146 14844
rect 22462 14832 22468 14884
rect 22520 14872 22526 14884
rect 24228 14872 24256 14912
rect 22520 14844 24256 14872
rect 24305 14875 24363 14881
rect 22520 14832 22526 14844
rect 24305 14841 24317 14875
rect 24351 14872 24363 14875
rect 25590 14872 25596 14884
rect 24351 14844 25596 14872
rect 24351 14841 24363 14844
rect 24305 14835 24363 14841
rect 25590 14832 25596 14844
rect 25648 14832 25654 14884
rect 25958 14832 25964 14884
rect 26016 14872 26022 14884
rect 27172 14872 27200 14968
rect 26016 14844 27200 14872
rect 28537 14875 28595 14881
rect 26016 14832 26022 14844
rect 28537 14841 28549 14875
rect 28583 14872 28595 14875
rect 28644 14872 28672 14968
rect 32309 14943 32367 14949
rect 32309 14909 32321 14943
rect 32355 14909 32367 14943
rect 32309 14903 32367 14909
rect 32585 14943 32643 14949
rect 32585 14909 32597 14943
rect 32631 14940 32643 14943
rect 32631 14912 33364 14940
rect 32631 14909 32643 14912
rect 32585 14903 32643 14909
rect 30006 14872 30012 14884
rect 28583 14844 30012 14872
rect 28583 14841 28595 14844
rect 28537 14835 28595 14841
rect 30006 14832 30012 14844
rect 30064 14832 30070 14884
rect 32324 14872 32352 14903
rect 33226 14872 33232 14884
rect 32324 14844 33232 14872
rect 33226 14832 33232 14844
rect 33284 14832 33290 14884
rect 19981 14807 20039 14813
rect 19981 14804 19993 14807
rect 19168 14776 19993 14804
rect 19981 14773 19993 14776
rect 20027 14773 20039 14807
rect 19981 14767 20039 14773
rect 22646 14764 22652 14816
rect 22704 14764 22710 14816
rect 22738 14764 22744 14816
rect 22796 14804 22802 14816
rect 23109 14807 23167 14813
rect 23109 14804 23121 14807
rect 22796 14776 23121 14804
rect 22796 14764 22802 14776
rect 23109 14773 23121 14776
rect 23155 14773 23167 14807
rect 23109 14767 23167 14773
rect 23290 14764 23296 14816
rect 23348 14804 23354 14816
rect 23385 14807 23443 14813
rect 23385 14804 23397 14807
rect 23348 14776 23397 14804
rect 23348 14764 23354 14776
rect 23385 14773 23397 14776
rect 23431 14773 23443 14807
rect 23385 14767 23443 14773
rect 25130 14764 25136 14816
rect 25188 14804 25194 14816
rect 25317 14807 25375 14813
rect 25317 14804 25329 14807
rect 25188 14776 25329 14804
rect 25188 14764 25194 14776
rect 25317 14773 25329 14776
rect 25363 14773 25375 14807
rect 25317 14767 25375 14773
rect 27709 14807 27767 14813
rect 27709 14773 27721 14807
rect 27755 14804 27767 14807
rect 27798 14804 27804 14816
rect 27755 14776 27804 14804
rect 27755 14773 27767 14776
rect 27709 14767 27767 14773
rect 27798 14764 27804 14776
rect 27856 14764 27862 14816
rect 28718 14764 28724 14816
rect 28776 14764 28782 14816
rect 33336 14804 33364 14912
rect 33502 14900 33508 14952
rect 33560 14900 33566 14952
rect 34716 14884 34744 14980
rect 35253 14977 35265 15011
rect 35299 14977 35311 15011
rect 37277 15011 37335 15017
rect 37277 15008 37289 15011
rect 36662 14994 37289 15008
rect 35253 14971 35311 14977
rect 36648 14980 37289 14994
rect 36078 14940 36084 14952
rect 35084 14912 36084 14940
rect 34698 14832 34704 14884
rect 34756 14872 34762 14884
rect 35084 14881 35112 14912
rect 36078 14900 36084 14912
rect 36136 14940 36142 14952
rect 36648 14940 36676 14980
rect 37277 14977 37289 14980
rect 37323 14977 37335 15011
rect 37277 14971 37335 14977
rect 37553 15011 37611 15017
rect 37553 14977 37565 15011
rect 37599 14977 37611 15011
rect 37553 14971 37611 14977
rect 39482 14968 39488 15020
rect 39540 14968 39546 15020
rect 39666 15017 39672 15020
rect 39633 15011 39672 15017
rect 39633 14977 39645 15011
rect 39633 14971 39672 14977
rect 39666 14968 39672 14971
rect 39724 14968 39730 15020
rect 39758 14968 39764 15020
rect 39816 14968 39822 15020
rect 39965 15017 39993 15116
rect 40126 15104 40132 15156
rect 40184 15144 40190 15156
rect 40221 15147 40279 15153
rect 40221 15144 40233 15147
rect 40184 15116 40233 15144
rect 40184 15104 40190 15116
rect 40221 15113 40233 15116
rect 40267 15113 40279 15147
rect 40221 15107 40279 15113
rect 42150 15104 42156 15156
rect 42208 15144 42214 15156
rect 42429 15147 42487 15153
rect 42429 15144 42441 15147
rect 42208 15116 42441 15144
rect 42208 15104 42214 15116
rect 42429 15113 42441 15116
rect 42475 15113 42487 15147
rect 42429 15107 42487 15113
rect 43346 15104 43352 15156
rect 43404 15104 43410 15156
rect 43438 15104 43444 15156
rect 43496 15144 43502 15156
rect 47673 15147 47731 15153
rect 47673 15144 47685 15147
rect 43496 15116 47685 15144
rect 43496 15104 43502 15116
rect 47673 15113 47685 15116
rect 47719 15144 47731 15147
rect 48130 15144 48136 15156
rect 47719 15116 48136 15144
rect 47719 15113 47731 15116
rect 47673 15107 47731 15113
rect 48130 15104 48136 15116
rect 48188 15104 48194 15156
rect 48222 15104 48228 15156
rect 48280 15144 48286 15156
rect 55950 15144 55956 15156
rect 48280 15104 48314 15144
rect 43364 15076 43392 15104
rect 43625 15079 43683 15085
rect 43625 15076 43637 15079
rect 43364 15048 43637 15076
rect 43625 15045 43637 15048
rect 43671 15045 43683 15079
rect 48286 15076 48314 15104
rect 51046 15116 55956 15144
rect 51046 15076 51074 15116
rect 55950 15104 55956 15116
rect 56008 15104 56014 15156
rect 56502 15104 56508 15156
rect 56560 15144 56566 15156
rect 56597 15147 56655 15153
rect 56597 15144 56609 15147
rect 56560 15116 56609 15144
rect 56560 15104 56566 15116
rect 56597 15113 56609 15116
rect 56643 15113 56655 15147
rect 56597 15107 56655 15113
rect 48286 15048 51074 15076
rect 55125 15079 55183 15085
rect 43625 15039 43683 15045
rect 39853 15011 39911 15017
rect 39853 14977 39865 15011
rect 39899 14977 39911 15011
rect 39853 14971 39911 14977
rect 39950 15011 40008 15017
rect 39950 14977 39962 15011
rect 39996 14977 40008 15011
rect 40405 15011 40463 15017
rect 40405 15008 40417 15011
rect 39950 14971 40008 14977
rect 40144 14980 40417 15008
rect 39868 14940 39896 14971
rect 36136 14912 36676 14940
rect 39316 14912 39896 14940
rect 36136 14900 36142 14912
rect 35069 14875 35127 14881
rect 35069 14872 35081 14875
rect 34756 14844 35081 14872
rect 34756 14832 34762 14844
rect 35069 14841 35081 14844
rect 35115 14841 35127 14875
rect 35069 14835 35127 14841
rect 39316 14816 39344 14912
rect 40144 14881 40172 14980
rect 40405 14977 40417 14980
rect 40451 14977 40463 15011
rect 40405 14971 40463 14977
rect 41046 14968 41052 15020
rect 41104 15008 41110 15020
rect 41104 14980 41414 15008
rect 41104 14968 41110 14980
rect 40681 14943 40739 14949
rect 40681 14909 40693 14943
rect 40727 14940 40739 14943
rect 41233 14943 41291 14949
rect 41233 14940 41245 14943
rect 40727 14912 41245 14940
rect 40727 14909 40739 14912
rect 40681 14903 40739 14909
rect 41233 14909 41245 14912
rect 41279 14909 41291 14943
rect 41386 14940 41414 14980
rect 41598 14968 41604 15020
rect 41656 15008 41662 15020
rect 41782 15008 41788 15020
rect 41656 14980 41788 15008
rect 41656 14968 41662 14980
rect 41782 14968 41788 14980
rect 41840 14968 41846 15020
rect 41969 15011 42027 15017
rect 41969 14977 41981 15011
rect 42015 14977 42027 15011
rect 41969 14971 42027 14977
rect 41984 14940 42012 14971
rect 42058 14968 42064 15020
rect 42116 15008 42122 15020
rect 42613 15011 42671 15017
rect 42613 15008 42625 15011
rect 42116 14980 42625 15008
rect 42116 14968 42122 14980
rect 42613 14977 42625 14980
rect 42659 14977 42671 15011
rect 42978 15008 42984 15020
rect 42613 14971 42671 14977
rect 42720 14980 42984 15008
rect 42720 14940 42748 14980
rect 42978 14968 42984 14980
rect 43036 14968 43042 15020
rect 43990 14968 43996 15020
rect 44048 15008 44054 15020
rect 44269 15011 44327 15017
rect 44269 15008 44281 15011
rect 44048 14980 44281 15008
rect 44048 14968 44054 14980
rect 44269 14977 44281 14980
rect 44315 14977 44327 15011
rect 44269 14971 44327 14977
rect 45554 14968 45560 15020
rect 45612 15008 45618 15020
rect 46477 15011 46535 15017
rect 46477 15008 46489 15011
rect 45612 14980 46489 15008
rect 45612 14968 45618 14980
rect 46477 14977 46489 14980
rect 46523 15008 46535 15011
rect 46658 15008 46664 15020
rect 46523 14980 46664 15008
rect 46523 14977 46535 14980
rect 46477 14971 46535 14977
rect 46658 14968 46664 14980
rect 46716 15008 46722 15020
rect 46845 15011 46903 15017
rect 46845 15008 46857 15011
rect 46716 14980 46857 15008
rect 46716 14968 46722 14980
rect 46845 14977 46857 14980
rect 46891 14977 46903 15011
rect 46845 14971 46903 14977
rect 48038 14968 48044 15020
rect 48096 14968 48102 15020
rect 48130 14968 48136 15020
rect 48188 14968 48194 15020
rect 49344 15017 49372 15048
rect 51000 15017 51028 15048
rect 55125 15045 55137 15079
rect 55171 15076 55183 15079
rect 55214 15076 55220 15088
rect 55171 15048 55220 15076
rect 55171 15045 55183 15048
rect 55125 15039 55183 15045
rect 55214 15036 55220 15048
rect 55272 15036 55278 15088
rect 55582 15036 55588 15088
rect 55640 15036 55646 15088
rect 48225 15011 48283 15017
rect 48225 14977 48237 15011
rect 48271 14977 48283 15011
rect 48225 14971 48283 14977
rect 48409 15011 48467 15017
rect 48409 14977 48421 15011
rect 48455 15008 48467 15011
rect 49329 15011 49387 15017
rect 48455 14980 49280 15008
rect 48455 14977 48467 14980
rect 48409 14971 48467 14977
rect 41386 14912 42748 14940
rect 42889 14943 42947 14949
rect 41233 14903 41291 14909
rect 42889 14909 42901 14943
rect 42935 14940 42947 14943
rect 43714 14940 43720 14952
rect 42935 14912 43720 14940
rect 42935 14909 42947 14912
rect 42889 14903 42947 14909
rect 43714 14900 43720 14912
rect 43772 14900 43778 14952
rect 44545 14943 44603 14949
rect 44545 14909 44557 14943
rect 44591 14940 44603 14943
rect 45097 14943 45155 14949
rect 45097 14940 45109 14943
rect 44591 14912 45109 14940
rect 44591 14909 44603 14912
rect 44545 14903 44603 14909
rect 45097 14909 45109 14912
rect 45143 14909 45155 14943
rect 45097 14903 45155 14909
rect 45370 14900 45376 14952
rect 45428 14940 45434 14952
rect 45649 14943 45707 14949
rect 45649 14940 45661 14943
rect 45428 14912 45661 14940
rect 45428 14900 45434 14912
rect 45649 14909 45661 14912
rect 45695 14909 45707 14943
rect 45649 14903 45707 14909
rect 47946 14900 47952 14952
rect 48004 14940 48010 14952
rect 48240 14940 48268 14971
rect 48004 14912 48268 14940
rect 49252 14940 49280 14980
rect 49329 14977 49341 15011
rect 49375 14977 49387 15011
rect 50525 15011 50583 15017
rect 50525 15008 50537 15011
rect 49329 14971 49387 14977
rect 50264 14980 50537 15008
rect 49694 14940 49700 14952
rect 49252 14912 49700 14940
rect 48004 14900 48010 14912
rect 49694 14900 49700 14912
rect 49752 14900 49758 14952
rect 40129 14875 40187 14881
rect 40129 14841 40141 14875
rect 40175 14841 40187 14875
rect 40129 14835 40187 14841
rect 40589 14875 40647 14881
rect 40589 14841 40601 14875
rect 40635 14872 40647 14875
rect 41414 14872 41420 14884
rect 40635 14844 41420 14872
rect 40635 14841 40647 14844
rect 40589 14835 40647 14841
rect 41414 14832 41420 14844
rect 41472 14872 41478 14884
rect 42797 14875 42855 14881
rect 42797 14872 42809 14875
rect 41472 14844 42809 14872
rect 41472 14832 41478 14844
rect 42797 14841 42809 14844
rect 42843 14841 42855 14875
rect 42797 14835 42855 14841
rect 43901 14875 43959 14881
rect 43901 14841 43913 14875
rect 43947 14872 43959 14875
rect 44358 14872 44364 14884
rect 43947 14844 44364 14872
rect 43947 14841 43959 14844
rect 43901 14835 43959 14841
rect 44358 14832 44364 14844
rect 44416 14832 44422 14884
rect 34238 14804 34244 14816
rect 33336 14776 34244 14804
rect 34238 14764 34244 14776
rect 34296 14764 34302 14816
rect 34790 14764 34796 14816
rect 34848 14804 34854 14816
rect 34977 14807 35035 14813
rect 34977 14804 34989 14807
rect 34848 14776 34989 14804
rect 34848 14764 34854 14776
rect 34977 14773 34989 14776
rect 35023 14773 35035 14807
rect 34977 14767 35035 14773
rect 36538 14764 36544 14816
rect 36596 14804 36602 14816
rect 36998 14804 37004 14816
rect 36596 14776 37004 14804
rect 36596 14764 36602 14776
rect 36998 14764 37004 14776
rect 37056 14764 37062 14816
rect 39298 14764 39304 14816
rect 39356 14764 39362 14816
rect 42150 14764 42156 14816
rect 42208 14804 42214 14816
rect 43622 14804 43628 14816
rect 42208 14776 43628 14804
rect 42208 14764 42214 14776
rect 43622 14764 43628 14776
rect 43680 14764 43686 14816
rect 44082 14764 44088 14816
rect 44140 14764 44146 14816
rect 44453 14807 44511 14813
rect 44453 14773 44465 14807
rect 44499 14804 44511 14807
rect 45002 14804 45008 14816
rect 44499 14776 45008 14804
rect 44499 14773 44511 14776
rect 44453 14767 44511 14773
rect 45002 14764 45008 14776
rect 45060 14764 45066 14816
rect 46661 14807 46719 14813
rect 46661 14773 46673 14807
rect 46707 14804 46719 14807
rect 47118 14804 47124 14816
rect 46707 14776 47124 14804
rect 46707 14773 46719 14776
rect 46661 14767 46719 14773
rect 47118 14764 47124 14776
rect 47176 14764 47182 14816
rect 47854 14764 47860 14816
rect 47912 14764 47918 14816
rect 48774 14764 48780 14816
rect 48832 14804 48838 14816
rect 49053 14807 49111 14813
rect 49053 14804 49065 14807
rect 48832 14776 49065 14804
rect 48832 14764 48838 14776
rect 49053 14773 49065 14776
rect 49099 14773 49111 14807
rect 49053 14767 49111 14773
rect 49510 14764 49516 14816
rect 49568 14804 49574 14816
rect 50264 14813 50292 14980
rect 50525 14977 50537 14980
rect 50571 14977 50583 15011
rect 50525 14971 50583 14977
rect 50985 15011 51043 15017
rect 50985 14977 50997 15011
rect 51031 14977 51043 15011
rect 50985 14971 51043 14977
rect 54018 14968 54024 15020
rect 54076 15008 54082 15020
rect 54849 15011 54907 15017
rect 54849 15008 54861 15011
rect 54076 14980 54861 15008
rect 54076 14968 54082 14980
rect 54849 14977 54861 14980
rect 54895 14977 54907 15011
rect 54849 14971 54907 14977
rect 51534 14872 51540 14884
rect 50632 14844 51540 14872
rect 50632 14816 50660 14844
rect 51534 14832 51540 14844
rect 51592 14832 51598 14884
rect 50249 14807 50307 14813
rect 50249 14804 50261 14807
rect 49568 14776 50261 14804
rect 49568 14764 49574 14776
rect 50249 14773 50261 14776
rect 50295 14773 50307 14807
rect 50249 14767 50307 14773
rect 50614 14764 50620 14816
rect 50672 14764 50678 14816
rect 50893 14807 50951 14813
rect 50893 14773 50905 14807
rect 50939 14804 50951 14807
rect 51810 14804 51816 14816
rect 50939 14776 51816 14804
rect 50939 14773 50951 14776
rect 50893 14767 50951 14773
rect 51810 14764 51816 14776
rect 51868 14764 51874 14816
rect 54202 14764 54208 14816
rect 54260 14764 54266 14816
rect 1104 14714 78844 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 78844 14714
rect 1104 14640 78844 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 8570 14600 8576 14612
rect 1627 14572 8576 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 14645 14603 14703 14609
rect 14645 14569 14657 14603
rect 14691 14600 14703 14603
rect 17954 14600 17960 14612
rect 14691 14572 17960 14600
rect 14691 14569 14703 14572
rect 14645 14563 14703 14569
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 18966 14560 18972 14612
rect 19024 14600 19030 14612
rect 19613 14603 19671 14609
rect 19613 14600 19625 14603
rect 19024 14572 19625 14600
rect 19024 14560 19030 14572
rect 19613 14569 19625 14572
rect 19659 14569 19671 14603
rect 19613 14563 19671 14569
rect 19702 14560 19708 14612
rect 19760 14560 19766 14612
rect 20073 14603 20131 14609
rect 20073 14569 20085 14603
rect 20119 14600 20131 14603
rect 20806 14600 20812 14612
rect 20119 14572 20812 14600
rect 20119 14569 20131 14572
rect 20073 14563 20131 14569
rect 20806 14560 20812 14572
rect 20864 14560 20870 14612
rect 22646 14560 22652 14612
rect 22704 14600 22710 14612
rect 22925 14603 22983 14609
rect 22925 14600 22937 14603
rect 22704 14572 22937 14600
rect 22704 14560 22710 14572
rect 22925 14569 22937 14572
rect 22971 14569 22983 14603
rect 22925 14563 22983 14569
rect 23198 14560 23204 14612
rect 23256 14560 23262 14612
rect 28166 14560 28172 14612
rect 28224 14560 28230 14612
rect 30650 14560 30656 14612
rect 30708 14600 30714 14612
rect 32030 14600 32036 14612
rect 30708 14572 32036 14600
rect 30708 14560 30714 14572
rect 32030 14560 32036 14572
rect 32088 14600 32094 14612
rect 33042 14600 33048 14612
rect 32088 14572 33048 14600
rect 32088 14560 32094 14572
rect 33042 14560 33048 14572
rect 33100 14560 33106 14612
rect 33226 14560 33232 14612
rect 33284 14600 33290 14612
rect 34149 14603 34207 14609
rect 34149 14600 34161 14603
rect 33284 14572 34161 14600
rect 33284 14560 33290 14572
rect 34149 14569 34161 14572
rect 34195 14600 34207 14603
rect 34422 14600 34428 14612
rect 34195 14572 34428 14600
rect 34195 14569 34207 14572
rect 34149 14563 34207 14569
rect 34422 14560 34428 14572
rect 34480 14560 34486 14612
rect 35342 14560 35348 14612
rect 35400 14600 35406 14612
rect 35529 14603 35587 14609
rect 35529 14600 35541 14603
rect 35400 14572 35541 14600
rect 35400 14560 35406 14572
rect 35529 14569 35541 14572
rect 35575 14569 35587 14603
rect 35529 14563 35587 14569
rect 37277 14603 37335 14609
rect 37277 14569 37289 14603
rect 37323 14600 37335 14603
rect 37918 14600 37924 14612
rect 37323 14572 37924 14600
rect 37323 14569 37335 14572
rect 37277 14563 37335 14569
rect 37918 14560 37924 14572
rect 37976 14560 37982 14612
rect 42058 14560 42064 14612
rect 42116 14560 42122 14612
rect 42334 14560 42340 14612
rect 42392 14600 42398 14612
rect 42981 14603 43039 14609
rect 42981 14600 42993 14603
rect 42392 14572 42993 14600
rect 42392 14560 42398 14572
rect 42981 14569 42993 14572
rect 43027 14600 43039 14603
rect 43070 14600 43076 14612
rect 43027 14572 43076 14600
rect 43027 14569 43039 14572
rect 42981 14563 43039 14569
rect 43070 14560 43076 14572
rect 43128 14600 43134 14612
rect 43898 14600 43904 14612
rect 43128 14572 43904 14600
rect 43128 14560 43134 14572
rect 43898 14560 43904 14572
rect 43956 14560 43962 14612
rect 43990 14560 43996 14612
rect 44048 14560 44054 14612
rect 45848 14572 47072 14600
rect 14090 14492 14096 14544
rect 14148 14492 14154 14544
rect 24762 14532 24768 14544
rect 22756 14504 24768 14532
rect 12434 14424 12440 14476
rect 12492 14464 12498 14476
rect 12621 14467 12679 14473
rect 12621 14464 12633 14467
rect 12492 14436 12633 14464
rect 12492 14424 12498 14436
rect 12621 14433 12633 14436
rect 12667 14433 12679 14467
rect 12621 14427 12679 14433
rect 1210 14356 1216 14408
rect 1268 14396 1274 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 1268 14368 1409 14396
rect 1268 14356 1274 14368
rect 1397 14365 1409 14368
rect 1443 14396 1455 14399
rect 1673 14399 1731 14405
rect 1673 14396 1685 14399
rect 1443 14368 1685 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 1673 14365 1685 14368
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 7650 14356 7656 14408
rect 7708 14356 7714 14408
rect 12342 14356 12348 14408
rect 12400 14356 12406 14408
rect 12636 14328 12664 14427
rect 13446 14424 13452 14476
rect 13504 14424 13510 14476
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 16482 14464 16488 14476
rect 14967 14436 16488 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 16669 14467 16727 14473
rect 16669 14433 16681 14467
rect 16715 14464 16727 14467
rect 16942 14464 16948 14476
rect 16715 14436 16948 14464
rect 16715 14433 16727 14436
rect 16669 14427 16727 14433
rect 16942 14424 16948 14436
rect 17000 14464 17006 14476
rect 17313 14467 17371 14473
rect 17313 14464 17325 14467
rect 17000 14436 17325 14464
rect 17000 14424 17006 14436
rect 17313 14433 17325 14436
rect 17359 14433 17371 14467
rect 17313 14427 17371 14433
rect 19610 14424 19616 14476
rect 19668 14464 19674 14476
rect 19797 14467 19855 14473
rect 19797 14464 19809 14467
rect 19668 14436 19809 14464
rect 19668 14424 19674 14436
rect 19797 14433 19809 14436
rect 19843 14433 19855 14467
rect 19797 14427 19855 14433
rect 20530 14424 20536 14476
rect 20588 14424 20594 14476
rect 14274 14356 14280 14408
rect 14332 14356 14338 14408
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14396 14427 14399
rect 14458 14396 14464 14408
rect 14415 14368 14464 14396
rect 14415 14365 14427 14368
rect 14369 14359 14427 14365
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 18506 14356 18512 14408
rect 18564 14396 18570 14408
rect 19058 14396 19064 14408
rect 18564 14368 19064 14396
rect 18564 14356 18570 14368
rect 19058 14356 19064 14368
rect 19116 14396 19122 14408
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 19116 14368 19257 14396
rect 19116 14356 19122 14368
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14396 20499 14399
rect 21450 14396 21456 14408
rect 20487 14368 21456 14396
rect 20487 14365 20499 14368
rect 20441 14359 20499 14365
rect 21450 14356 21456 14368
rect 21508 14356 21514 14408
rect 22370 14356 22376 14408
rect 22428 14396 22434 14408
rect 22756 14405 22784 14504
rect 24762 14492 24768 14504
rect 24820 14492 24826 14544
rect 27706 14532 27712 14544
rect 26160 14504 27712 14532
rect 23017 14467 23075 14473
rect 23017 14433 23029 14467
rect 23063 14464 23075 14467
rect 23290 14464 23296 14476
rect 23063 14436 23296 14464
rect 23063 14433 23075 14436
rect 23017 14427 23075 14433
rect 23290 14424 23296 14436
rect 23348 14424 23354 14476
rect 23566 14424 23572 14476
rect 23624 14464 23630 14476
rect 24854 14464 24860 14476
rect 23624 14436 24860 14464
rect 23624 14424 23630 14436
rect 24854 14424 24860 14436
rect 24912 14424 24918 14476
rect 22741 14399 22799 14405
rect 22741 14396 22753 14399
rect 22428 14368 22753 14396
rect 22428 14356 22434 14368
rect 22741 14365 22753 14368
rect 22787 14365 22799 14399
rect 22741 14359 22799 14365
rect 23106 14356 23112 14408
rect 23164 14396 23170 14408
rect 23201 14399 23259 14405
rect 23201 14396 23213 14399
rect 23164 14368 23213 14396
rect 23164 14356 23170 14368
rect 23201 14365 23213 14368
rect 23247 14365 23259 14399
rect 23201 14359 23259 14365
rect 23382 14356 23388 14408
rect 23440 14396 23446 14408
rect 23661 14399 23719 14405
rect 23661 14396 23673 14399
rect 23440 14368 23673 14396
rect 23440 14356 23446 14368
rect 23661 14365 23673 14368
rect 23707 14396 23719 14399
rect 26160 14396 26188 14504
rect 27706 14492 27712 14504
rect 27764 14492 27770 14544
rect 27985 14535 28043 14541
rect 27985 14501 27997 14535
rect 28031 14532 28043 14535
rect 28031 14504 28212 14532
rect 28031 14501 28043 14504
rect 27985 14495 28043 14501
rect 27154 14424 27160 14476
rect 27212 14464 27218 14476
rect 28074 14464 28080 14476
rect 27212 14436 27477 14464
rect 27212 14424 27218 14436
rect 23707 14368 26188 14396
rect 23707 14365 23719 14368
rect 23661 14359 23719 14365
rect 26878 14356 26884 14408
rect 26936 14396 26942 14408
rect 27338 14396 27344 14408
rect 26936 14368 27344 14396
rect 26936 14356 26942 14368
rect 27338 14356 27344 14368
rect 27396 14356 27402 14408
rect 27449 14405 27477 14436
rect 27908 14436 28080 14464
rect 27434 14399 27492 14405
rect 27434 14365 27446 14399
rect 27480 14365 27492 14399
rect 27434 14359 27492 14365
rect 27522 14356 27528 14408
rect 27580 14396 27586 14408
rect 27632 14405 27849 14406
rect 27632 14399 27864 14405
rect 27632 14396 27818 14399
rect 27580 14378 27818 14396
rect 27580 14368 27660 14378
rect 27580 14356 27586 14368
rect 27806 14365 27818 14378
rect 27852 14365 27864 14399
rect 27806 14359 27864 14365
rect 15102 14328 15108 14340
rect 12636 14300 15108 14328
rect 15102 14288 15108 14300
rect 15160 14288 15166 14340
rect 15194 14288 15200 14340
rect 15252 14288 15258 14340
rect 17589 14331 17647 14337
rect 15580 14300 15686 14328
rect 16500 14300 16896 14328
rect 7834 14220 7840 14272
rect 7892 14220 7898 14272
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 11977 14263 12035 14269
rect 11977 14260 11989 14263
rect 11848 14232 11989 14260
rect 11848 14220 11854 14232
rect 11977 14229 11989 14232
rect 12023 14229 12035 14263
rect 11977 14223 12035 14229
rect 12437 14263 12495 14269
rect 12437 14229 12449 14263
rect 12483 14260 12495 14263
rect 12897 14263 12955 14269
rect 12897 14260 12909 14263
rect 12483 14232 12909 14260
rect 12483 14229 12495 14232
rect 12437 14223 12495 14229
rect 12897 14229 12909 14232
rect 12943 14229 12955 14263
rect 12897 14223 12955 14229
rect 14458 14220 14464 14272
rect 14516 14220 14522 14272
rect 14918 14220 14924 14272
rect 14976 14260 14982 14272
rect 15580 14260 15608 14300
rect 16500 14260 16528 14300
rect 14976 14232 16528 14260
rect 14976 14220 14982 14232
rect 16758 14220 16764 14272
rect 16816 14220 16822 14272
rect 16868 14260 16896 14300
rect 17589 14297 17601 14331
rect 17635 14328 17647 14331
rect 17635 14300 18184 14328
rect 17635 14297 17647 14300
rect 17589 14291 17647 14297
rect 18156 14269 18184 14300
rect 23290 14288 23296 14340
rect 23348 14328 23354 14340
rect 24762 14328 24768 14340
rect 23348 14300 24768 14328
rect 23348 14288 23354 14300
rect 17681 14263 17739 14269
rect 17681 14260 17693 14263
rect 16868 14232 17693 14260
rect 17681 14229 17693 14232
rect 17727 14229 17739 14263
rect 17681 14223 17739 14229
rect 18141 14263 18199 14269
rect 18141 14229 18153 14263
rect 18187 14260 18199 14263
rect 18322 14260 18328 14272
rect 18187 14232 18328 14260
rect 18187 14229 18199 14232
rect 18141 14223 18199 14229
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 20809 14263 20867 14269
rect 20809 14229 20821 14263
rect 20855 14260 20867 14263
rect 20898 14260 20904 14272
rect 20855 14232 20904 14260
rect 20855 14229 20867 14232
rect 20809 14223 20867 14229
rect 20898 14220 20904 14232
rect 20956 14220 20962 14272
rect 22554 14220 22560 14272
rect 22612 14220 22618 14272
rect 22646 14220 22652 14272
rect 22704 14260 22710 14272
rect 23382 14260 23388 14272
rect 22704 14232 23388 14260
rect 22704 14220 22710 14232
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 23569 14263 23627 14269
rect 23569 14229 23581 14263
rect 23615 14260 23627 14263
rect 23658 14260 23664 14272
rect 23615 14232 23664 14260
rect 23615 14229 23627 14232
rect 23569 14223 23627 14229
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 23860 14269 23888 14300
rect 24762 14288 24768 14300
rect 24820 14288 24826 14340
rect 26970 14288 26976 14340
rect 27028 14328 27034 14340
rect 27617 14331 27675 14337
rect 27617 14328 27629 14331
rect 27028 14300 27629 14328
rect 27028 14288 27034 14300
rect 27617 14297 27629 14300
rect 27663 14297 27675 14331
rect 27617 14291 27675 14297
rect 27709 14331 27767 14337
rect 27709 14297 27721 14331
rect 27755 14328 27767 14331
rect 27908 14328 27936 14436
rect 28074 14424 28080 14436
rect 28132 14424 28138 14476
rect 28184 14464 28212 14504
rect 33870 14492 33876 14544
rect 33928 14532 33934 14544
rect 34793 14535 34851 14541
rect 34793 14532 34805 14535
rect 33928 14504 34805 14532
rect 33928 14492 33934 14504
rect 34793 14501 34805 14504
rect 34839 14501 34851 14535
rect 34793 14495 34851 14501
rect 35084 14504 37320 14532
rect 28184 14436 28396 14464
rect 27755 14300 27936 14328
rect 27755 14297 27767 14300
rect 27709 14291 27767 14297
rect 23845 14263 23903 14269
rect 23845 14229 23857 14263
rect 23891 14229 23903 14263
rect 23845 14223 23903 14229
rect 24302 14220 24308 14272
rect 24360 14260 24366 14272
rect 26234 14260 26240 14272
rect 24360 14232 26240 14260
rect 24360 14220 24366 14232
rect 26234 14220 26240 14232
rect 26292 14220 26298 14272
rect 28074 14220 28080 14272
rect 28132 14260 28138 14272
rect 28368 14260 28396 14436
rect 29454 14424 29460 14476
rect 29512 14464 29518 14476
rect 29730 14464 29736 14476
rect 29512 14436 29736 14464
rect 29512 14424 29518 14436
rect 29730 14424 29736 14436
rect 29788 14464 29794 14476
rect 31297 14467 31355 14473
rect 31297 14464 31309 14467
rect 29788 14436 31309 14464
rect 29788 14424 29794 14436
rect 31297 14433 31309 14436
rect 31343 14464 31355 14467
rect 31570 14464 31576 14476
rect 31343 14436 31576 14464
rect 31343 14433 31355 14436
rect 31297 14427 31355 14433
rect 31570 14424 31576 14436
rect 31628 14424 31634 14476
rect 29546 14356 29552 14408
rect 29604 14396 29610 14408
rect 30285 14399 30343 14405
rect 30285 14396 30297 14399
rect 29604 14368 30297 14396
rect 29604 14356 29610 14368
rect 30285 14365 30297 14368
rect 30331 14365 30343 14399
rect 30285 14359 30343 14365
rect 30469 14399 30527 14405
rect 30469 14365 30481 14399
rect 30515 14396 30527 14399
rect 30926 14396 30932 14408
rect 30515 14368 30932 14396
rect 30515 14365 30527 14368
rect 30469 14359 30527 14365
rect 30926 14356 30932 14368
rect 30984 14356 30990 14408
rect 33134 14356 33140 14408
rect 33192 14356 33198 14408
rect 33410 14356 33416 14408
rect 33468 14396 33474 14408
rect 34977 14399 35035 14405
rect 34977 14396 34989 14399
rect 33468 14368 34989 14396
rect 33468 14356 33474 14368
rect 34977 14365 34989 14368
rect 35023 14396 35035 14399
rect 35084 14396 35112 14504
rect 37292 14476 37320 14504
rect 39666 14492 39672 14544
rect 39724 14532 39730 14544
rect 43346 14532 43352 14544
rect 39724 14504 42564 14532
rect 39724 14492 39730 14504
rect 35802 14424 35808 14476
rect 35860 14464 35866 14476
rect 36814 14464 36820 14476
rect 35860 14436 36308 14464
rect 35860 14424 35866 14436
rect 35023 14368 35112 14396
rect 35708 14399 35766 14405
rect 35023 14365 35035 14368
rect 34977 14359 35035 14365
rect 35708 14365 35720 14399
rect 35754 14396 35766 14399
rect 36080 14399 36138 14405
rect 35754 14368 36032 14396
rect 35754 14365 35766 14368
rect 35708 14359 35766 14365
rect 31570 14288 31576 14340
rect 31628 14288 31634 14340
rect 32858 14328 32864 14340
rect 32798 14300 32864 14328
rect 32858 14288 32864 14300
rect 32916 14288 32922 14340
rect 33502 14288 33508 14340
rect 33560 14328 33566 14340
rect 34790 14328 34796 14340
rect 33560 14300 34796 14328
rect 33560 14288 33566 14300
rect 34790 14288 34796 14300
rect 34848 14328 34854 14340
rect 35802 14328 35808 14340
rect 34848 14300 35808 14328
rect 34848 14288 34854 14300
rect 35802 14288 35808 14300
rect 35860 14288 35866 14340
rect 35897 14331 35955 14337
rect 35897 14297 35909 14331
rect 35943 14297 35955 14331
rect 35897 14291 35955 14297
rect 28132 14232 28396 14260
rect 30101 14263 30159 14269
rect 28132 14220 28138 14232
rect 30101 14229 30113 14263
rect 30147 14260 30159 14263
rect 30374 14260 30380 14272
rect 30147 14232 30380 14260
rect 30147 14229 30159 14232
rect 30101 14223 30159 14229
rect 30374 14220 30380 14232
rect 30432 14220 30438 14272
rect 31938 14220 31944 14272
rect 31996 14260 32002 14272
rect 33045 14263 33103 14269
rect 33045 14260 33057 14263
rect 31996 14232 33057 14260
rect 31996 14220 32002 14232
rect 33045 14229 33057 14232
rect 33091 14260 33103 14263
rect 33962 14260 33968 14272
rect 33091 14232 33968 14260
rect 33091 14229 33103 14232
rect 33045 14223 33103 14229
rect 33962 14220 33968 14232
rect 34020 14220 34026 14272
rect 34146 14220 34152 14272
rect 34204 14260 34210 14272
rect 35342 14260 35348 14272
rect 34204 14232 35348 14260
rect 34204 14220 34210 14232
rect 35342 14220 35348 14232
rect 35400 14260 35406 14272
rect 35912 14260 35940 14291
rect 35400 14232 35940 14260
rect 36004 14260 36032 14368
rect 36080 14365 36092 14399
rect 36126 14365 36138 14399
rect 36080 14359 36138 14365
rect 36096 14328 36124 14359
rect 36170 14356 36176 14408
rect 36228 14356 36234 14408
rect 36280 14405 36308 14436
rect 36464 14436 36820 14464
rect 36464 14405 36492 14436
rect 36814 14424 36820 14436
rect 36872 14464 36878 14476
rect 37093 14467 37151 14473
rect 37093 14464 37105 14467
rect 36872 14436 37105 14464
rect 36872 14424 36878 14436
rect 37093 14433 37105 14436
rect 37139 14464 37151 14467
rect 37182 14464 37188 14476
rect 37139 14436 37188 14464
rect 37139 14433 37151 14436
rect 37093 14427 37151 14433
rect 37182 14424 37188 14436
rect 37240 14424 37246 14476
rect 37274 14424 37280 14476
rect 37332 14424 37338 14476
rect 37550 14424 37556 14476
rect 37608 14424 37614 14476
rect 39758 14464 39764 14476
rect 37660 14436 39764 14464
rect 36265 14399 36323 14405
rect 36265 14365 36277 14399
rect 36311 14365 36323 14399
rect 36265 14359 36323 14365
rect 36449 14399 36507 14405
rect 36449 14365 36461 14399
rect 36495 14365 36507 14399
rect 36449 14359 36507 14365
rect 36630 14356 36636 14408
rect 36688 14356 36694 14408
rect 37456 14399 37514 14405
rect 37456 14396 37468 14399
rect 36740 14368 37468 14396
rect 36354 14328 36360 14340
rect 36096 14300 36360 14328
rect 36354 14288 36360 14300
rect 36412 14288 36418 14340
rect 36538 14288 36544 14340
rect 36596 14288 36602 14340
rect 36740 14260 36768 14368
rect 37456 14365 37468 14368
rect 37502 14396 37514 14399
rect 37568 14396 37596 14424
rect 37660 14405 37688 14436
rect 39758 14424 39764 14436
rect 39816 14424 39822 14476
rect 39850 14424 39856 14476
rect 39908 14464 39914 14476
rect 39908 14436 41460 14464
rect 39908 14424 39914 14436
rect 37502 14368 37596 14396
rect 37645 14399 37703 14405
rect 37502 14365 37514 14368
rect 37456 14359 37514 14365
rect 37645 14365 37657 14399
rect 37691 14365 37703 14399
rect 37645 14359 37703 14365
rect 37828 14399 37886 14405
rect 37828 14365 37840 14399
rect 37874 14365 37886 14399
rect 37828 14359 37886 14365
rect 37921 14399 37979 14405
rect 37921 14365 37933 14399
rect 37967 14396 37979 14399
rect 39482 14396 39488 14408
rect 37967 14368 39488 14396
rect 37967 14365 37979 14368
rect 37921 14359 37979 14365
rect 36998 14288 37004 14340
rect 37056 14328 37062 14340
rect 37553 14331 37611 14337
rect 37553 14328 37565 14331
rect 37056 14300 37565 14328
rect 37056 14288 37062 14300
rect 37553 14297 37565 14300
rect 37599 14297 37611 14331
rect 37553 14291 37611 14297
rect 36004 14232 36768 14260
rect 35400 14220 35406 14232
rect 36814 14220 36820 14272
rect 36872 14220 36878 14272
rect 36906 14220 36912 14272
rect 36964 14220 36970 14272
rect 37734 14220 37740 14272
rect 37792 14260 37798 14272
rect 37845 14260 37873 14359
rect 39482 14356 39488 14368
rect 39540 14356 39546 14408
rect 39776 14328 39804 14424
rect 41432 14405 41460 14436
rect 42334 14424 42340 14476
rect 42392 14424 42398 14476
rect 41417 14399 41475 14405
rect 41417 14365 41429 14399
rect 41463 14365 41475 14399
rect 41417 14359 41475 14365
rect 41506 14356 41512 14408
rect 41564 14396 41570 14408
rect 41564 14368 41609 14396
rect 41564 14356 41570 14368
rect 41782 14356 41788 14408
rect 41840 14356 41846 14408
rect 41923 14399 41981 14405
rect 41923 14365 41935 14399
rect 41969 14396 41981 14399
rect 42150 14396 42156 14408
rect 41969 14368 42156 14396
rect 41969 14365 41981 14368
rect 41923 14359 41981 14365
rect 42150 14356 42156 14368
rect 42208 14356 42214 14408
rect 42352 14396 42380 14424
rect 42536 14405 42564 14504
rect 43272 14504 43352 14532
rect 43272 14464 43300 14504
rect 43346 14492 43352 14504
rect 43404 14492 43410 14544
rect 44453 14535 44511 14541
rect 44453 14532 44465 14535
rect 43456 14504 44465 14532
rect 43456 14464 43484 14504
rect 44453 14501 44465 14504
rect 44499 14532 44511 14535
rect 44910 14532 44916 14544
rect 44499 14504 44916 14532
rect 44499 14501 44511 14504
rect 44453 14495 44511 14501
rect 44910 14492 44916 14504
rect 44968 14532 44974 14544
rect 45848 14532 45876 14572
rect 44968 14504 45876 14532
rect 47044 14532 47072 14572
rect 47486 14560 47492 14612
rect 47544 14560 47550 14612
rect 50798 14600 50804 14612
rect 48056 14572 50804 14600
rect 47762 14532 47768 14544
rect 47044 14504 47768 14532
rect 44968 14492 44974 14504
rect 47762 14492 47768 14504
rect 47820 14492 47826 14544
rect 42725 14436 43300 14464
rect 43364 14436 43484 14464
rect 42429 14399 42487 14405
rect 42429 14396 42441 14399
rect 42352 14368 42441 14396
rect 42429 14365 42441 14368
rect 42475 14365 42487 14399
rect 42429 14359 42487 14365
rect 42521 14399 42579 14405
rect 42521 14365 42533 14399
rect 42567 14396 42579 14399
rect 42725 14396 42753 14436
rect 42567 14368 42753 14396
rect 42567 14365 42579 14368
rect 42521 14359 42579 14365
rect 42794 14356 42800 14408
rect 42852 14356 42858 14408
rect 43364 14405 43392 14436
rect 43622 14424 43628 14476
rect 43680 14464 43686 14476
rect 44634 14464 44640 14476
rect 43680 14436 44640 14464
rect 43680 14424 43686 14436
rect 43349 14399 43407 14405
rect 43349 14365 43361 14399
rect 43395 14365 43407 14399
rect 43349 14359 43407 14365
rect 43442 14399 43500 14405
rect 43442 14365 43454 14399
rect 43488 14365 43500 14399
rect 43442 14359 43500 14365
rect 41690 14328 41696 14340
rect 39776 14300 41696 14328
rect 41690 14288 41696 14300
rect 41748 14288 41754 14340
rect 41800 14260 41828 14356
rect 42613 14331 42671 14337
rect 42613 14328 42625 14331
rect 41892 14300 42625 14328
rect 41892 14272 41920 14300
rect 42613 14297 42625 14300
rect 42659 14297 42671 14331
rect 42812 14328 42840 14356
rect 43457 14328 43485 14359
rect 43530 14356 43536 14408
rect 43588 14396 43594 14408
rect 43870 14405 43898 14436
rect 44634 14424 44640 14436
rect 44692 14424 44698 14476
rect 45094 14424 45100 14476
rect 45152 14464 45158 14476
rect 45738 14464 45744 14476
rect 45152 14436 45744 14464
rect 45152 14424 45158 14436
rect 45738 14424 45744 14436
rect 45796 14424 45802 14476
rect 46750 14424 46756 14476
rect 46808 14464 46814 14476
rect 47780 14464 47808 14492
rect 46808 14436 47164 14464
rect 46808 14424 46814 14436
rect 43717 14399 43775 14405
rect 43717 14396 43729 14399
rect 43588 14368 43729 14396
rect 43588 14356 43594 14368
rect 43717 14365 43729 14368
rect 43763 14365 43775 14399
rect 43717 14359 43775 14365
rect 43855 14399 43913 14405
rect 43855 14365 43867 14399
rect 43901 14365 43913 14399
rect 47136 14396 47164 14436
rect 47688 14436 47808 14464
rect 47302 14396 47308 14408
rect 43855 14359 43913 14365
rect 44100 14368 45324 14396
rect 47136 14382 47308 14396
rect 47150 14368 47308 14382
rect 42812 14300 43485 14328
rect 43625 14331 43683 14337
rect 42613 14291 42671 14297
rect 43625 14297 43637 14331
rect 43671 14328 43683 14331
rect 44100 14328 44128 14368
rect 43671 14300 44128 14328
rect 44177 14331 44235 14337
rect 43671 14297 43683 14300
rect 43625 14291 43683 14297
rect 44177 14297 44189 14331
rect 44223 14328 44235 14331
rect 44358 14328 44364 14340
rect 44223 14300 44364 14328
rect 44223 14297 44235 14300
rect 44177 14291 44235 14297
rect 37792 14232 41828 14260
rect 37792 14220 37798 14232
rect 41874 14220 41880 14272
rect 41932 14220 41938 14272
rect 42242 14220 42248 14272
rect 42300 14220 42306 14272
rect 42628 14260 42656 14291
rect 44358 14288 44364 14300
rect 44416 14328 44422 14340
rect 44637 14331 44695 14337
rect 44637 14328 44649 14331
rect 44416 14300 44649 14328
rect 44416 14288 44422 14300
rect 44637 14297 44649 14300
rect 44683 14297 44695 14331
rect 44637 14291 44695 14297
rect 45002 14288 45008 14340
rect 45060 14288 45066 14340
rect 45186 14288 45192 14340
rect 45244 14288 45250 14340
rect 45296 14272 45324 14368
rect 47302 14356 47308 14368
rect 47360 14396 47366 14408
rect 47578 14396 47584 14408
rect 47360 14368 47584 14396
rect 47360 14356 47366 14368
rect 47578 14356 47584 14368
rect 47636 14356 47642 14408
rect 47688 14405 47716 14436
rect 47673 14399 47731 14405
rect 47673 14365 47685 14399
rect 47719 14365 47731 14399
rect 47673 14359 47731 14365
rect 47821 14399 47879 14405
rect 47821 14365 47833 14399
rect 47867 14396 47879 14399
rect 48056 14396 48084 14572
rect 50798 14560 50804 14572
rect 50856 14560 50862 14612
rect 51074 14600 51080 14612
rect 50908 14572 51080 14600
rect 48317 14535 48375 14541
rect 48317 14501 48329 14535
rect 48363 14501 48375 14535
rect 48317 14495 48375 14501
rect 47867 14368 48084 14396
rect 47867 14365 47879 14368
rect 47821 14359 47879 14365
rect 48130 14356 48136 14408
rect 48188 14405 48194 14408
rect 48188 14396 48196 14405
rect 48332 14396 48360 14495
rect 50430 14492 50436 14544
rect 50488 14532 50494 14544
rect 50488 14504 50568 14532
rect 50488 14492 50494 14504
rect 49694 14424 49700 14476
rect 49752 14464 49758 14476
rect 49878 14464 49884 14476
rect 49752 14436 49884 14464
rect 49752 14424 49758 14436
rect 49878 14424 49884 14436
rect 49936 14464 49942 14476
rect 49973 14467 50031 14473
rect 49973 14464 49985 14467
rect 49936 14436 49985 14464
rect 49936 14424 49942 14436
rect 49973 14433 49985 14436
rect 50019 14464 50031 14467
rect 50019 14436 50476 14464
rect 50019 14433 50031 14436
rect 49973 14427 50031 14433
rect 50448 14408 50476 14436
rect 48593 14399 48651 14405
rect 48593 14396 48605 14399
rect 48188 14368 48233 14396
rect 48332 14368 48605 14396
rect 48188 14359 48196 14368
rect 48593 14365 48605 14368
rect 48639 14365 48651 14399
rect 48593 14359 48651 14365
rect 48188 14356 48194 14359
rect 48774 14356 48780 14408
rect 48832 14356 48838 14408
rect 48869 14399 48927 14405
rect 48869 14365 48881 14399
rect 48915 14396 48927 14399
rect 49329 14399 49387 14405
rect 49329 14396 49341 14399
rect 48915 14368 49341 14396
rect 48915 14365 48927 14368
rect 48869 14359 48927 14365
rect 49329 14365 49341 14368
rect 49375 14365 49387 14399
rect 49329 14359 49387 14365
rect 50341 14399 50399 14405
rect 50341 14365 50353 14399
rect 50387 14365 50399 14399
rect 50341 14359 50399 14365
rect 46014 14288 46020 14340
rect 46072 14288 46078 14340
rect 47946 14328 47952 14340
rect 47320 14300 47952 14328
rect 43073 14263 43131 14269
rect 43073 14260 43085 14263
rect 42628 14232 43085 14260
rect 43073 14229 43085 14232
rect 43119 14229 43131 14263
rect 43073 14223 43131 14229
rect 45278 14220 45284 14272
rect 45336 14260 45342 14272
rect 47320 14260 47348 14300
rect 47946 14288 47952 14300
rect 48004 14288 48010 14340
rect 48041 14331 48099 14337
rect 48041 14297 48053 14331
rect 48087 14297 48099 14331
rect 50356 14328 50384 14359
rect 50430 14356 50436 14408
rect 50488 14356 50494 14408
rect 50540 14337 50568 14504
rect 50709 14399 50767 14405
rect 50709 14365 50721 14399
rect 50755 14396 50767 14399
rect 50908 14396 50936 14572
rect 51074 14560 51080 14572
rect 51132 14600 51138 14612
rect 53558 14600 53564 14612
rect 51132 14572 53564 14600
rect 51132 14560 51138 14572
rect 53558 14560 53564 14572
rect 53616 14560 53622 14612
rect 51350 14492 51356 14544
rect 51408 14532 51414 14544
rect 51408 14504 51488 14532
rect 51408 14492 51414 14504
rect 50982 14424 50988 14476
rect 51040 14464 51046 14476
rect 51040 14436 51212 14464
rect 51040 14424 51046 14436
rect 51184 14405 51212 14436
rect 51460 14405 51488 14504
rect 54202 14492 54208 14544
rect 54260 14532 54266 14544
rect 54260 14504 55076 14532
rect 54260 14492 54266 14504
rect 51084 14399 51142 14405
rect 51084 14396 51096 14399
rect 50755 14368 50936 14396
rect 51000 14368 51096 14396
rect 50755 14365 50767 14368
rect 50709 14359 50767 14365
rect 51000 14340 51028 14368
rect 51084 14365 51096 14368
rect 51130 14365 51142 14399
rect 51084 14359 51142 14365
rect 51170 14399 51228 14405
rect 51170 14365 51182 14399
rect 51216 14365 51228 14399
rect 51170 14359 51228 14365
rect 51445 14399 51503 14405
rect 51445 14365 51457 14399
rect 51491 14365 51503 14399
rect 51445 14359 51503 14365
rect 51534 14356 51540 14408
rect 51592 14405 51598 14408
rect 51592 14399 51619 14405
rect 51607 14365 51619 14399
rect 51592 14359 51619 14365
rect 51592 14356 51598 14359
rect 51718 14356 51724 14408
rect 51776 14396 51782 14408
rect 51813 14399 51871 14405
rect 51813 14396 51825 14399
rect 51776 14368 51825 14396
rect 51776 14356 51782 14368
rect 51813 14365 51825 14368
rect 51859 14365 51871 14399
rect 51813 14359 51871 14365
rect 53558 14356 53564 14408
rect 53616 14396 53622 14408
rect 54570 14405 54576 14408
rect 54205 14399 54263 14405
rect 54205 14396 54217 14399
rect 53616 14368 54217 14396
rect 53616 14356 53622 14368
rect 54205 14365 54217 14368
rect 54251 14365 54263 14399
rect 54568 14396 54576 14405
rect 54531 14368 54576 14396
rect 54205 14359 54263 14365
rect 54568 14359 54576 14368
rect 50525 14331 50583 14337
rect 50356 14300 50476 14328
rect 48041 14291 48099 14297
rect 45336 14232 47348 14260
rect 45336 14220 45342 14232
rect 47486 14220 47492 14272
rect 47544 14260 47550 14272
rect 48056 14260 48084 14291
rect 50448 14272 50476 14300
rect 50525 14297 50537 14331
rect 50571 14297 50583 14331
rect 50525 14291 50583 14297
rect 50982 14288 50988 14340
rect 51040 14288 51046 14340
rect 51353 14331 51411 14337
rect 51353 14328 51365 14331
rect 51276 14300 51365 14328
rect 51276 14272 51304 14300
rect 51353 14297 51365 14300
rect 51399 14297 51411 14331
rect 51353 14291 51411 14297
rect 52086 14288 52092 14340
rect 52144 14288 52150 14340
rect 52546 14288 52552 14340
rect 52604 14288 52610 14340
rect 53466 14288 53472 14340
rect 53524 14328 53530 14340
rect 53653 14331 53711 14337
rect 53653 14328 53665 14331
rect 53524 14300 53665 14328
rect 53524 14288 53530 14300
rect 53653 14297 53665 14300
rect 53699 14297 53711 14331
rect 54220 14328 54248 14359
rect 54570 14356 54576 14359
rect 54628 14356 54634 14408
rect 54754 14356 54760 14408
rect 54812 14356 54818 14408
rect 54938 14396 54944 14408
rect 54899 14368 54944 14396
rect 54938 14356 54944 14368
rect 54996 14356 55002 14408
rect 55048 14405 55076 14504
rect 55033 14399 55091 14405
rect 55033 14365 55045 14399
rect 55079 14365 55091 14399
rect 55033 14359 55091 14365
rect 54665 14331 54723 14337
rect 54665 14328 54677 14331
rect 54220 14300 54677 14328
rect 53653 14291 53711 14297
rect 54665 14297 54677 14300
rect 54711 14297 54723 14331
rect 54665 14291 54723 14297
rect 47544 14232 48084 14260
rect 47544 14220 47550 14232
rect 48406 14220 48412 14272
rect 48464 14220 48470 14272
rect 50157 14263 50215 14269
rect 50157 14229 50169 14263
rect 50203 14260 50215 14263
rect 50246 14260 50252 14272
rect 50203 14232 50252 14260
rect 50203 14229 50215 14232
rect 50157 14223 50215 14229
rect 50246 14220 50252 14232
rect 50304 14220 50310 14272
rect 50430 14220 50436 14272
rect 50488 14260 50494 14272
rect 50614 14260 50620 14272
rect 50488 14232 50620 14260
rect 50488 14220 50494 14232
rect 50614 14220 50620 14232
rect 50672 14220 50678 14272
rect 51258 14220 51264 14272
rect 51316 14220 51322 14272
rect 51721 14263 51779 14269
rect 51721 14229 51733 14263
rect 51767 14260 51779 14263
rect 52178 14260 52184 14272
rect 51767 14232 52184 14260
rect 51767 14229 51779 14232
rect 51721 14223 51779 14229
rect 52178 14220 52184 14232
rect 52236 14220 52242 14272
rect 54110 14220 54116 14272
rect 54168 14260 54174 14272
rect 54389 14263 54447 14269
rect 54389 14260 54401 14263
rect 54168 14232 54401 14260
rect 54168 14220 54174 14232
rect 54389 14229 54401 14232
rect 54435 14229 54447 14263
rect 54389 14223 54447 14229
rect 1104 14170 78844 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 66314 14170
rect 66366 14118 66378 14170
rect 66430 14118 66442 14170
rect 66494 14118 66506 14170
rect 66558 14118 66570 14170
rect 66622 14118 78844 14170
rect 1104 14096 78844 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 7650 14056 7656 14068
rect 1627 14028 7656 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 12710 14056 12716 14068
rect 11532 14028 12716 14056
rect 7834 13948 7840 14000
rect 7892 13988 7898 14000
rect 8205 13991 8263 13997
rect 8205 13988 8217 13991
rect 7892 13960 8217 13988
rect 7892 13948 7898 13960
rect 8205 13957 8217 13960
rect 8251 13957 8263 13991
rect 10870 13988 10876 14000
rect 9430 13960 10876 13988
rect 8205 13951 8263 13957
rect 10870 13948 10876 13960
rect 10928 13948 10934 14000
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 11532 13929 11560 14028
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 13265 14059 13323 14065
rect 13265 14025 13277 14059
rect 13311 14056 13323 14059
rect 13446 14056 13452 14068
rect 13311 14028 13452 14056
rect 13311 14025 13323 14028
rect 13265 14019 13323 14025
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 15749 14059 15807 14065
rect 15749 14056 15761 14059
rect 15252 14028 15761 14056
rect 15252 14016 15258 14028
rect 15749 14025 15761 14028
rect 15795 14025 15807 14059
rect 15749 14019 15807 14025
rect 16209 14059 16267 14065
rect 16209 14025 16221 14059
rect 16255 14056 16267 14059
rect 16758 14056 16764 14068
rect 16255 14028 16764 14056
rect 16255 14025 16267 14028
rect 16209 14019 16267 14025
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 21450 14016 21456 14068
rect 21508 14016 21514 14068
rect 22189 14059 22247 14065
rect 22189 14025 22201 14059
rect 22235 14056 22247 14059
rect 23106 14056 23112 14068
rect 22235 14028 23112 14056
rect 22235 14025 22247 14028
rect 22189 14019 22247 14025
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 25498 14056 25504 14068
rect 23216 14028 24716 14056
rect 11790 13948 11796 14000
rect 11848 13948 11854 14000
rect 12250 13948 12256 14000
rect 12308 13948 12314 14000
rect 18417 13991 18475 13997
rect 18417 13988 18429 13991
rect 17788 13960 18429 13988
rect 1673 13923 1731 13929
rect 1673 13920 1685 13923
rect 1452 13892 1685 13920
rect 1452 13880 1458 13892
rect 1673 13889 1685 13892
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16850 13920 16856 13932
rect 16163 13892 16856 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 7929 13855 7987 13861
rect 7929 13821 7941 13855
rect 7975 13852 7987 13855
rect 9398 13852 9404 13864
rect 7975 13824 9404 13852
rect 7975 13821 7987 13824
rect 7929 13815 7987 13821
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13852 9735 13855
rect 16132 13852 16160 13883
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17402 13880 17408 13932
rect 17460 13920 17466 13932
rect 17788 13929 17816 13960
rect 18417 13957 18429 13960
rect 18463 13957 18475 13991
rect 18417 13951 18475 13957
rect 17773 13923 17831 13929
rect 17773 13920 17785 13923
rect 17460 13892 17785 13920
rect 17460 13880 17466 13892
rect 17773 13889 17785 13892
rect 17819 13889 17831 13923
rect 17773 13883 17831 13889
rect 17954 13880 17960 13932
rect 18012 13920 18018 13932
rect 18233 13923 18291 13929
rect 18233 13920 18245 13923
rect 18012 13892 18245 13920
rect 18012 13880 18018 13892
rect 18233 13889 18245 13892
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13920 18567 13923
rect 19242 13920 19248 13932
rect 18555 13892 19248 13920
rect 18555 13889 18567 13892
rect 18509 13883 18567 13889
rect 19242 13880 19248 13892
rect 19300 13880 19306 13932
rect 21545 13923 21603 13929
rect 21545 13889 21557 13923
rect 21591 13920 21603 13923
rect 22370 13920 22376 13932
rect 21591 13892 22376 13920
rect 21591 13889 21603 13892
rect 21545 13883 21603 13889
rect 22370 13880 22376 13892
rect 22428 13880 22434 13932
rect 22462 13880 22468 13932
rect 22520 13920 22526 13932
rect 22557 13923 22615 13929
rect 22557 13920 22569 13923
rect 22520 13892 22569 13920
rect 22520 13880 22526 13892
rect 22557 13889 22569 13892
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 22738 13920 22744 13932
rect 22695 13892 22744 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 22738 13880 22744 13892
rect 22796 13880 22802 13932
rect 22925 13923 22983 13929
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 22925 13883 22983 13889
rect 9723 13824 16160 13852
rect 9723 13821 9735 13824
rect 9677 13815 9735 13821
rect 16390 13812 16396 13864
rect 16448 13812 16454 13864
rect 22940 13852 22968 13883
rect 23014 13880 23020 13932
rect 23072 13920 23078 13932
rect 23216 13929 23244 14028
rect 23382 13948 23388 14000
rect 23440 13988 23446 14000
rect 24688 13997 24716 14028
rect 25240 14028 25504 14056
rect 25240 13997 25268 14028
rect 25498 14016 25504 14028
rect 25556 14016 25562 14068
rect 25777 14059 25835 14065
rect 25777 14025 25789 14059
rect 25823 14056 25835 14059
rect 28353 14059 28411 14065
rect 25823 14028 27936 14056
rect 25823 14025 25835 14028
rect 25777 14019 25835 14025
rect 24029 13991 24087 13997
rect 24029 13988 24041 13991
rect 23440 13960 24041 13988
rect 23440 13948 23446 13960
rect 24029 13957 24041 13960
rect 24075 13988 24087 13991
rect 24673 13991 24731 13997
rect 24075 13960 24532 13988
rect 24075 13957 24087 13960
rect 24029 13951 24087 13957
rect 23201 13923 23259 13929
rect 23201 13920 23213 13923
rect 23072 13892 23213 13920
rect 23072 13880 23078 13892
rect 23201 13889 23213 13892
rect 23247 13889 23259 13923
rect 23474 13920 23480 13932
rect 23201 13883 23259 13889
rect 23308 13892 23480 13920
rect 23308 13852 23336 13892
rect 23474 13880 23480 13892
rect 23532 13880 23538 13932
rect 23658 13880 23664 13932
rect 23716 13880 23722 13932
rect 23842 13929 23848 13932
rect 23809 13923 23848 13929
rect 23809 13889 23821 13923
rect 23809 13883 23848 13889
rect 23842 13880 23848 13883
rect 23900 13880 23906 13932
rect 23934 13880 23940 13932
rect 23992 13880 23998 13932
rect 24118 13880 24124 13932
rect 24176 13929 24182 13932
rect 24504 13929 24532 13960
rect 24673 13957 24685 13991
rect 24719 13957 24731 13991
rect 24673 13951 24731 13957
rect 25225 13991 25283 13997
rect 25225 13957 25237 13991
rect 25271 13957 25283 13991
rect 26329 13991 26387 13997
rect 26329 13988 26341 13991
rect 25225 13951 25283 13957
rect 25332 13960 26341 13988
rect 25332 13932 25360 13960
rect 26329 13957 26341 13960
rect 26375 13957 26387 13991
rect 26329 13951 26387 13957
rect 27522 13948 27528 14000
rect 27580 13948 27586 14000
rect 27908 13997 27936 14028
rect 28353 14025 28365 14059
rect 28399 14056 28411 14059
rect 28810 14056 28816 14068
rect 28399 14028 28816 14056
rect 28399 14025 28411 14028
rect 28353 14019 28411 14025
rect 28810 14016 28816 14028
rect 28868 14016 28874 14068
rect 31481 14059 31539 14065
rect 31481 14025 31493 14059
rect 31527 14056 31539 14059
rect 31570 14056 31576 14068
rect 31527 14028 31576 14056
rect 31527 14025 31539 14028
rect 31481 14019 31539 14025
rect 31570 14016 31576 14028
rect 31628 14016 31634 14068
rect 32217 14059 32275 14065
rect 32217 14025 32229 14059
rect 32263 14025 32275 14059
rect 32217 14019 32275 14025
rect 27893 13991 27951 13997
rect 27893 13957 27905 13991
rect 27939 13957 27951 13991
rect 31202 13988 31208 14000
rect 31050 13960 31208 13988
rect 27893 13951 27951 13957
rect 31202 13948 31208 13960
rect 31260 13988 31266 14000
rect 32122 13988 32128 14000
rect 31260 13960 32128 13988
rect 31260 13948 31266 13960
rect 32122 13948 32128 13960
rect 32180 13948 32186 14000
rect 24176 13920 24184 13929
rect 24397 13923 24455 13929
rect 24176 13892 24221 13920
rect 24176 13883 24184 13892
rect 24397 13889 24409 13923
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 24490 13923 24548 13929
rect 24490 13889 24502 13923
rect 24536 13889 24548 13923
rect 24490 13883 24548 13889
rect 24765 13923 24823 13929
rect 24765 13889 24777 13923
rect 24811 13889 24823 13923
rect 24765 13883 24823 13889
rect 24176 13880 24182 13883
rect 22940 13824 23336 13852
rect 23385 13855 23443 13861
rect 23385 13821 23397 13855
rect 23431 13852 23443 13855
rect 24412 13852 24440 13883
rect 23431 13824 24440 13852
rect 24780 13852 24808 13883
rect 24854 13880 24860 13932
rect 24912 13929 24918 13932
rect 24912 13920 24920 13929
rect 25133 13923 25191 13929
rect 24912 13892 24957 13920
rect 24912 13883 24920 13892
rect 25133 13889 25145 13923
rect 25179 13920 25191 13923
rect 25314 13920 25320 13932
rect 25179 13892 25320 13920
rect 25179 13889 25191 13892
rect 25133 13883 25191 13889
rect 24912 13880 24918 13883
rect 25314 13880 25320 13892
rect 25372 13880 25378 13932
rect 25498 13880 25504 13932
rect 25556 13880 25562 13932
rect 25590 13880 25596 13932
rect 25648 13880 25654 13932
rect 26053 13923 26111 13929
rect 26053 13889 26065 13923
rect 26099 13889 26111 13923
rect 26053 13883 26111 13889
rect 24780 13824 24992 13852
rect 23431 13821 23443 13824
rect 23385 13815 23443 13821
rect 24302 13744 24308 13796
rect 24360 13744 24366 13796
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 18141 13719 18199 13725
rect 18141 13716 18153 13719
rect 18104 13688 18153 13716
rect 18104 13676 18110 13688
rect 18141 13685 18153 13688
rect 18187 13685 18199 13719
rect 18141 13679 18199 13685
rect 18509 13719 18567 13725
rect 18509 13685 18521 13719
rect 18555 13716 18567 13719
rect 18874 13716 18880 13728
rect 18555 13688 18880 13716
rect 18555 13685 18567 13688
rect 18509 13679 18567 13685
rect 18874 13676 18880 13688
rect 18932 13676 18938 13728
rect 24964 13716 24992 13824
rect 25958 13812 25964 13864
rect 26016 13812 26022 13864
rect 26068 13852 26096 13883
rect 26142 13880 26148 13932
rect 26200 13880 26206 13932
rect 27338 13880 27344 13932
rect 27396 13880 27402 13932
rect 27430 13880 27436 13932
rect 27488 13880 27494 13932
rect 27706 13880 27712 13932
rect 27764 13880 27770 13932
rect 27798 13880 27804 13932
rect 27856 13880 27862 13932
rect 28074 13880 28080 13932
rect 28132 13880 28138 13932
rect 28169 13923 28227 13929
rect 28169 13889 28181 13923
rect 28215 13889 28227 13923
rect 28169 13883 28227 13889
rect 31665 13923 31723 13929
rect 31665 13889 31677 13923
rect 31711 13920 31723 13923
rect 32232 13920 32260 14019
rect 32582 14016 32588 14068
rect 32640 14016 32646 14068
rect 32858 14016 32864 14068
rect 32916 14056 32922 14068
rect 33137 14059 33195 14065
rect 33137 14056 33149 14059
rect 32916 14028 33149 14056
rect 32916 14016 32922 14028
rect 33137 14025 33149 14028
rect 33183 14025 33195 14059
rect 33137 14019 33195 14025
rect 36170 14016 36176 14068
rect 36228 14056 36234 14068
rect 39850 14056 39856 14068
rect 36228 14028 39856 14056
rect 36228 14016 36234 14028
rect 39850 14016 39856 14028
rect 39908 14016 39914 14068
rect 45738 14056 45744 14068
rect 41386 14028 45744 14056
rect 32493 13991 32551 13997
rect 32493 13957 32505 13991
rect 32539 13988 32551 13991
rect 32600 13988 32628 14016
rect 33502 13988 33508 14000
rect 32539 13960 32628 13988
rect 32784 13960 33508 13988
rect 32539 13957 32551 13960
rect 32493 13951 32551 13957
rect 32398 13929 32404 13932
rect 32396 13920 32404 13929
rect 31711 13892 32260 13920
rect 32359 13892 32404 13920
rect 31711 13889 31723 13892
rect 31665 13883 31723 13889
rect 32396 13883 32404 13892
rect 26418 13852 26424 13864
rect 26068 13824 26424 13852
rect 26418 13812 26424 13824
rect 26476 13812 26482 13864
rect 27062 13812 27068 13864
rect 27120 13852 27126 13864
rect 28184 13852 28212 13883
rect 32398 13880 32404 13883
rect 32456 13880 32462 13932
rect 27120 13824 28212 13852
rect 27120 13812 27126 13824
rect 29454 13812 29460 13864
rect 29512 13852 29518 13864
rect 29549 13855 29607 13861
rect 29549 13852 29561 13855
rect 29512 13824 29561 13852
rect 29512 13812 29518 13824
rect 29549 13821 29561 13824
rect 29595 13821 29607 13855
rect 29549 13815 29607 13821
rect 29822 13812 29828 13864
rect 29880 13812 29886 13864
rect 31938 13812 31944 13864
rect 31996 13812 32002 13864
rect 32508 13852 32536 13951
rect 32784 13929 32812 13960
rect 33502 13948 33508 13960
rect 33560 13948 33566 14000
rect 36188 13988 36216 14016
rect 33704 13960 36216 13988
rect 32585 13923 32643 13929
rect 32585 13889 32597 13923
rect 32631 13889 32643 13923
rect 32585 13883 32643 13889
rect 32768 13923 32826 13929
rect 32768 13889 32780 13923
rect 32814 13889 32826 13923
rect 32768 13883 32826 13889
rect 32861 13923 32919 13929
rect 32861 13889 32873 13923
rect 32907 13920 32919 13923
rect 33042 13920 33048 13932
rect 32907 13892 33048 13920
rect 32907 13889 32919 13892
rect 32861 13883 32919 13889
rect 32048 13824 32536 13852
rect 32600 13852 32628 13883
rect 33042 13880 33048 13892
rect 33100 13920 33106 13932
rect 33704 13920 33732 13960
rect 33100 13892 33732 13920
rect 33100 13880 33106 13892
rect 33778 13880 33784 13932
rect 33836 13920 33842 13932
rect 33919 13923 33977 13929
rect 33919 13920 33931 13923
rect 33836 13892 33931 13920
rect 33836 13880 33842 13892
rect 33919 13889 33931 13892
rect 33965 13889 33977 13923
rect 33919 13883 33977 13889
rect 34054 13880 34060 13932
rect 34112 13880 34118 13932
rect 34146 13880 34152 13932
rect 34204 13880 34210 13932
rect 34440 13929 34468 13960
rect 36262 13948 36268 14000
rect 36320 13948 36326 14000
rect 36354 13948 36360 14000
rect 36412 13988 36418 14000
rect 39298 13988 39304 14000
rect 36412 13960 39304 13988
rect 36412 13948 36418 13960
rect 39298 13948 39304 13960
rect 39356 13948 39362 14000
rect 39574 13948 39580 14000
rect 39632 13988 39638 14000
rect 40865 13991 40923 13997
rect 40865 13988 40877 13991
rect 39632 13960 40877 13988
rect 39632 13948 39638 13960
rect 34332 13923 34390 13929
rect 34332 13889 34344 13923
rect 34378 13889 34390 13923
rect 34332 13883 34390 13889
rect 34425 13923 34483 13929
rect 34425 13889 34437 13923
rect 34471 13889 34483 13923
rect 34425 13883 34483 13889
rect 33594 13852 33600 13864
rect 32600 13824 33600 13852
rect 25038 13744 25044 13796
rect 25096 13744 25102 13796
rect 25682 13744 25688 13796
rect 25740 13784 25746 13796
rect 25869 13787 25927 13793
rect 25869 13784 25881 13787
rect 25740 13756 25881 13784
rect 25740 13744 25746 13756
rect 25869 13753 25881 13756
rect 25915 13753 25927 13787
rect 25869 13747 25927 13753
rect 30926 13744 30932 13796
rect 30984 13784 30990 13796
rect 31297 13787 31355 13793
rect 31297 13784 31309 13787
rect 30984 13756 31309 13784
rect 30984 13744 30990 13756
rect 31297 13753 31309 13756
rect 31343 13784 31355 13787
rect 32048 13784 32076 13824
rect 33594 13812 33600 13824
rect 33652 13852 33658 13864
rect 34164 13852 34192 13880
rect 33652 13824 34192 13852
rect 34348 13852 34376 13883
rect 35986 13880 35992 13932
rect 36044 13920 36050 13932
rect 36081 13923 36139 13929
rect 36081 13920 36093 13923
rect 36044 13892 36093 13920
rect 36044 13880 36050 13892
rect 36081 13889 36093 13892
rect 36127 13889 36139 13923
rect 36081 13883 36139 13889
rect 36446 13880 36452 13932
rect 36504 13920 36510 13932
rect 36817 13923 36875 13929
rect 36817 13920 36829 13923
rect 36504 13892 36829 13920
rect 36504 13880 36510 13892
rect 36817 13889 36829 13892
rect 36863 13920 36875 13923
rect 38838 13920 38844 13932
rect 36863 13892 38844 13920
rect 36863 13889 36875 13892
rect 36817 13883 36875 13889
rect 38838 13880 38844 13892
rect 38896 13880 38902 13932
rect 40586 13880 40592 13932
rect 40644 13880 40650 13932
rect 40788 13929 40816 13960
rect 40865 13957 40877 13960
rect 40911 13957 40923 13991
rect 40865 13951 40923 13957
rect 40773 13923 40831 13929
rect 40773 13889 40785 13923
rect 40819 13920 40831 13923
rect 41386 13920 41414 14028
rect 45738 14016 45744 14028
rect 45796 14016 45802 14068
rect 46014 14016 46020 14068
rect 46072 14056 46078 14068
rect 46385 14059 46443 14065
rect 46385 14056 46397 14059
rect 46072 14028 46397 14056
rect 46072 14016 46078 14028
rect 46385 14025 46397 14028
rect 46431 14025 46443 14059
rect 46750 14056 46756 14068
rect 46385 14019 46443 14025
rect 46584 14028 46756 14056
rect 44082 13948 44088 14000
rect 44140 13948 44146 14000
rect 46584 13988 46612 14028
rect 46750 14016 46756 14028
rect 46808 14016 46814 14068
rect 46934 14016 46940 14068
rect 46992 14056 46998 14068
rect 47121 14059 47179 14065
rect 47121 14056 47133 14059
rect 46992 14028 47133 14056
rect 46992 14016 46998 14028
rect 47121 14025 47133 14028
rect 47167 14056 47179 14059
rect 47486 14056 47492 14068
rect 47167 14028 47492 14056
rect 47167 14025 47179 14028
rect 47121 14019 47179 14025
rect 47486 14016 47492 14028
rect 47544 14056 47550 14068
rect 47581 14059 47639 14065
rect 47581 14056 47593 14059
rect 47544 14028 47593 14056
rect 47544 14016 47550 14028
rect 47581 14025 47593 14028
rect 47627 14025 47639 14059
rect 47581 14019 47639 14025
rect 47670 14016 47676 14068
rect 47728 14056 47734 14068
rect 51718 14056 51724 14068
rect 47728 14028 49280 14056
rect 47728 14016 47734 14028
rect 47854 13988 47860 14000
rect 45310 13960 46612 13988
rect 46676 13960 47860 13988
rect 46676 13929 46704 13960
rect 47854 13948 47860 13960
rect 47912 13948 47918 14000
rect 48133 13991 48191 13997
rect 48133 13957 48145 13991
rect 48179 13988 48191 13991
rect 48406 13988 48412 14000
rect 48179 13960 48412 13988
rect 48179 13957 48191 13960
rect 48133 13951 48191 13957
rect 48406 13948 48412 13960
rect 48464 13948 48470 14000
rect 49252 13932 49280 14028
rect 49896 14028 51724 14056
rect 40819 13892 41414 13920
rect 46569 13923 46627 13929
rect 40819 13889 40831 13892
rect 40773 13883 40831 13889
rect 46569 13889 46581 13923
rect 46615 13889 46627 13923
rect 46569 13883 46627 13889
rect 46661 13923 46719 13929
rect 46661 13889 46673 13923
rect 46707 13889 46719 13923
rect 46661 13883 46719 13889
rect 36538 13852 36544 13864
rect 34348 13824 36544 13852
rect 33652 13812 33658 13824
rect 36538 13812 36544 13824
rect 36596 13812 36602 13864
rect 36909 13855 36967 13861
rect 36909 13852 36921 13855
rect 36648 13824 36921 13852
rect 34238 13784 34244 13796
rect 31343 13756 32076 13784
rect 32140 13756 34244 13784
rect 31343 13753 31355 13756
rect 31297 13747 31355 13753
rect 26602 13716 26608 13728
rect 24964 13688 26608 13716
rect 26602 13676 26608 13688
rect 26660 13716 26666 13728
rect 26786 13716 26792 13728
rect 26660 13688 26792 13716
rect 26660 13676 26666 13688
rect 26786 13676 26792 13688
rect 26844 13676 26850 13728
rect 27154 13676 27160 13728
rect 27212 13676 27218 13728
rect 27614 13676 27620 13728
rect 27672 13716 27678 13728
rect 27893 13719 27951 13725
rect 27893 13716 27905 13719
rect 27672 13688 27905 13716
rect 27672 13676 27678 13688
rect 27893 13685 27905 13688
rect 27939 13685 27951 13719
rect 27893 13679 27951 13685
rect 31849 13719 31907 13725
rect 31849 13685 31861 13719
rect 31895 13716 31907 13719
rect 32140 13716 32168 13756
rect 34238 13744 34244 13756
rect 34296 13744 34302 13796
rect 36262 13744 36268 13796
rect 36320 13784 36326 13796
rect 36648 13784 36676 13824
rect 36909 13821 36921 13824
rect 36955 13821 36967 13855
rect 36909 13815 36967 13821
rect 40497 13855 40555 13861
rect 40497 13821 40509 13855
rect 40543 13852 40555 13855
rect 43809 13855 43867 13861
rect 40543 13824 40632 13852
rect 40543 13821 40555 13824
rect 40497 13815 40555 13821
rect 36320 13756 36676 13784
rect 40313 13787 40371 13793
rect 36320 13744 36326 13756
rect 40313 13753 40325 13787
rect 40359 13784 40371 13787
rect 40604 13784 40632 13824
rect 43809 13821 43821 13855
rect 43855 13852 43867 13855
rect 46584 13852 46612 13883
rect 46934 13880 46940 13932
rect 46992 13880 46998 13932
rect 49234 13880 49240 13932
rect 49292 13880 49298 13932
rect 49896 13929 49924 14028
rect 51718 14016 51724 14028
rect 51776 14016 51782 14068
rect 52270 14016 52276 14068
rect 52328 14056 52334 14068
rect 54202 14056 54208 14068
rect 52328 14028 54208 14056
rect 52328 14016 52334 14028
rect 54202 14016 54208 14028
rect 54260 14016 54266 14068
rect 51534 13988 51540 14000
rect 51382 13960 51540 13988
rect 51534 13948 51540 13960
rect 51592 13948 51598 14000
rect 51736 13988 51764 14016
rect 54018 13988 54024 14000
rect 51736 13960 54024 13988
rect 49881 13923 49939 13929
rect 49881 13889 49893 13923
rect 49927 13889 49939 13923
rect 49881 13883 49939 13889
rect 51997 13923 52055 13929
rect 51997 13889 52009 13923
rect 52043 13920 52055 13923
rect 52086 13920 52092 13932
rect 52043 13892 52092 13920
rect 52043 13889 52055 13892
rect 51997 13883 52055 13889
rect 52086 13880 52092 13892
rect 52144 13880 52150 13932
rect 52178 13880 52184 13932
rect 52236 13880 52242 13932
rect 52457 13923 52515 13929
rect 52457 13889 52469 13923
rect 52503 13920 52515 13923
rect 53466 13920 53472 13932
rect 52503 13892 53472 13920
rect 52503 13889 52515 13892
rect 52457 13883 52515 13889
rect 53466 13880 53472 13892
rect 53524 13880 53530 13932
rect 53668 13929 53696 13960
rect 54018 13948 54024 13960
rect 54076 13948 54082 14000
rect 53653 13923 53711 13929
rect 53653 13889 53665 13923
rect 53699 13889 53711 13923
rect 55582 13920 55588 13932
rect 55062 13906 55588 13920
rect 53653 13883 53711 13889
rect 55048 13892 55588 13906
rect 43855 13824 43944 13852
rect 46584 13824 46796 13852
rect 43855 13821 43867 13824
rect 43809 13815 43867 13821
rect 42242 13784 42248 13796
rect 40359 13756 40540 13784
rect 40604 13756 42248 13784
rect 40359 13753 40371 13756
rect 40313 13747 40371 13753
rect 31895 13688 32168 13716
rect 33045 13719 33103 13725
rect 31895 13685 31907 13688
rect 31849 13679 31907 13685
rect 33045 13685 33057 13719
rect 33091 13716 33103 13719
rect 33134 13716 33140 13728
rect 33091 13688 33140 13716
rect 33091 13685 33103 13688
rect 33045 13679 33103 13685
rect 33134 13676 33140 13688
rect 33192 13676 33198 13728
rect 33686 13676 33692 13728
rect 33744 13716 33750 13728
rect 33781 13719 33839 13725
rect 33781 13716 33793 13719
rect 33744 13688 33793 13716
rect 33744 13676 33750 13688
rect 33781 13685 33793 13688
rect 33827 13685 33839 13719
rect 33781 13679 33839 13685
rect 36630 13676 36636 13728
rect 36688 13676 36694 13728
rect 39390 13676 39396 13728
rect 39448 13716 39454 13728
rect 40037 13719 40095 13725
rect 40037 13716 40049 13719
rect 39448 13688 40049 13716
rect 39448 13676 39454 13688
rect 40037 13685 40049 13688
rect 40083 13685 40095 13719
rect 40037 13679 40095 13685
rect 40402 13676 40408 13728
rect 40460 13676 40466 13728
rect 40512 13716 40540 13756
rect 42242 13744 42248 13756
rect 42300 13744 42306 13796
rect 41966 13716 41972 13728
rect 40512 13688 41972 13716
rect 41966 13676 41972 13688
rect 42024 13676 42030 13728
rect 43916 13716 43944 13824
rect 46768 13784 46796 13824
rect 46842 13812 46848 13864
rect 46900 13852 46906 13864
rect 47857 13855 47915 13861
rect 47857 13852 47869 13855
rect 46900 13824 47869 13852
rect 46900 13812 46906 13824
rect 47857 13821 47869 13824
rect 47903 13821 47915 13855
rect 47857 13815 47915 13821
rect 49605 13855 49663 13861
rect 49605 13821 49617 13855
rect 49651 13852 49663 13855
rect 49651 13824 49924 13852
rect 49651 13821 49663 13824
rect 49605 13815 49663 13821
rect 49896 13796 49924 13824
rect 50154 13812 50160 13864
rect 50212 13812 50218 13864
rect 50614 13812 50620 13864
rect 50672 13852 50678 13864
rect 50798 13852 50804 13864
rect 50672 13824 50804 13852
rect 50672 13812 50678 13824
rect 50798 13812 50804 13824
rect 50856 13852 50862 13864
rect 51350 13852 51356 13864
rect 50856 13824 51356 13852
rect 50856 13812 50862 13824
rect 51350 13812 51356 13824
rect 51408 13852 51414 13864
rect 51629 13855 51687 13861
rect 51629 13852 51641 13855
rect 51408 13824 51641 13852
rect 51408 13812 51414 13824
rect 51629 13821 51641 13824
rect 51675 13821 51687 13855
rect 54938 13852 54944 13864
rect 51629 13815 51687 13821
rect 52564 13824 54944 13852
rect 52564 13796 52592 13824
rect 54938 13812 54944 13824
rect 54996 13852 55002 13864
rect 55048 13852 55076 13892
rect 55582 13880 55588 13892
rect 55640 13880 55646 13932
rect 54996 13824 55076 13852
rect 54996 13812 55002 13824
rect 47118 13784 47124 13796
rect 46768 13756 47124 13784
rect 47118 13744 47124 13756
rect 47176 13784 47182 13796
rect 47762 13784 47768 13796
rect 47176 13756 47768 13784
rect 47176 13744 47182 13756
rect 47762 13744 47768 13756
rect 47820 13744 47826 13796
rect 49878 13744 49884 13796
rect 49936 13744 49942 13796
rect 51534 13744 51540 13796
rect 51592 13784 51598 13796
rect 52546 13784 52552 13796
rect 51592 13756 52552 13784
rect 51592 13744 51598 13756
rect 52546 13744 52552 13756
rect 52604 13744 52610 13796
rect 45094 13716 45100 13728
rect 43916 13688 45100 13716
rect 45094 13676 45100 13688
rect 45152 13676 45158 13728
rect 45370 13676 45376 13728
rect 45428 13716 45434 13728
rect 45557 13719 45615 13725
rect 45557 13716 45569 13719
rect 45428 13688 45569 13716
rect 45428 13676 45434 13688
rect 45557 13685 45569 13688
rect 45603 13685 45615 13719
rect 45557 13679 45615 13685
rect 46845 13719 46903 13725
rect 46845 13685 46857 13719
rect 46891 13716 46903 13719
rect 46934 13716 46940 13728
rect 46891 13688 46940 13716
rect 46891 13685 46903 13688
rect 46845 13679 46903 13685
rect 46934 13676 46940 13688
rect 46992 13676 46998 13728
rect 51166 13676 51172 13728
rect 51224 13716 51230 13728
rect 51810 13716 51816 13728
rect 51224 13688 51816 13716
rect 51224 13676 51230 13688
rect 51810 13676 51816 13688
rect 51868 13716 51874 13728
rect 52362 13716 52368 13728
rect 51868 13688 52368 13716
rect 51868 13676 51874 13688
rect 52362 13676 52368 13688
rect 52420 13676 52426 13728
rect 53926 13725 53932 13728
rect 53916 13719 53932 13725
rect 53916 13685 53928 13719
rect 53916 13679 53932 13685
rect 53926 13676 53932 13679
rect 53984 13676 53990 13728
rect 55398 13676 55404 13728
rect 55456 13676 55462 13728
rect 1104 13626 78844 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 78844 13626
rect 1104 13552 78844 13574
rect 18601 13515 18659 13521
rect 18601 13512 18613 13515
rect 17696 13484 18613 13512
rect 9033 13379 9091 13385
rect 9033 13345 9045 13379
rect 9079 13376 9091 13379
rect 9398 13376 9404 13388
rect 9079 13348 9404 13376
rect 9079 13345 9091 13348
rect 9033 13339 9091 13345
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 8570 13268 8576 13320
rect 8628 13268 8634 13320
rect 16390 13268 16396 13320
rect 16448 13308 16454 13320
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 16448 13280 17233 13308
rect 16448 13268 16454 13280
rect 17221 13277 17233 13280
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 9309 13243 9367 13249
rect 9309 13209 9321 13243
rect 9355 13209 9367 13243
rect 10870 13240 10876 13252
rect 10534 13212 10876 13240
rect 9309 13203 9367 13209
rect 8757 13175 8815 13181
rect 8757 13141 8769 13175
rect 8803 13172 8815 13175
rect 9324 13172 9352 13203
rect 10870 13200 10876 13212
rect 10928 13200 10934 13252
rect 16942 13200 16948 13252
rect 17000 13200 17006 13252
rect 17236 13240 17264 13271
rect 17310 13268 17316 13320
rect 17368 13268 17374 13320
rect 17402 13268 17408 13320
rect 17460 13308 17466 13320
rect 17696 13317 17724 13484
rect 18601 13481 18613 13484
rect 18647 13481 18659 13515
rect 18601 13475 18659 13481
rect 21542 13472 21548 13524
rect 21600 13472 21606 13524
rect 21729 13515 21787 13521
rect 21729 13481 21741 13515
rect 21775 13512 21787 13515
rect 23014 13512 23020 13524
rect 21775 13484 23020 13512
rect 21775 13481 21787 13484
rect 21729 13475 21787 13481
rect 23014 13472 23020 13484
rect 23072 13472 23078 13524
rect 23198 13472 23204 13524
rect 23256 13472 23262 13524
rect 27430 13472 27436 13524
rect 27488 13472 27494 13524
rect 29178 13472 29184 13524
rect 29236 13472 29242 13524
rect 29822 13472 29828 13524
rect 29880 13512 29886 13524
rect 29917 13515 29975 13521
rect 29917 13512 29929 13515
rect 29880 13484 29929 13512
rect 29880 13472 29886 13484
rect 29917 13481 29929 13484
rect 29963 13481 29975 13515
rect 29917 13475 29975 13481
rect 32122 13472 32128 13524
rect 32180 13512 32186 13524
rect 32493 13515 32551 13521
rect 32493 13512 32505 13515
rect 32180 13484 32505 13512
rect 32180 13472 32186 13484
rect 32493 13481 32505 13484
rect 32539 13481 32551 13515
rect 32493 13475 32551 13481
rect 36630 13472 36636 13524
rect 36688 13512 36694 13524
rect 37093 13515 37151 13521
rect 37093 13512 37105 13515
rect 36688 13484 37105 13512
rect 36688 13472 36694 13484
rect 37093 13481 37105 13484
rect 37139 13481 37151 13515
rect 37093 13475 37151 13481
rect 37826 13472 37832 13524
rect 37884 13512 37890 13524
rect 38378 13512 38384 13524
rect 37884 13484 38384 13512
rect 37884 13472 37890 13484
rect 38378 13472 38384 13484
rect 38436 13512 38442 13524
rect 38933 13515 38991 13521
rect 38933 13512 38945 13515
rect 38436 13484 38945 13512
rect 38436 13472 38442 13484
rect 38933 13481 38945 13484
rect 38979 13481 38991 13515
rect 38933 13475 38991 13481
rect 39390 13472 39396 13524
rect 39448 13472 39454 13524
rect 40402 13472 40408 13524
rect 40460 13472 40466 13524
rect 40494 13472 40500 13524
rect 40552 13472 40558 13524
rect 41509 13515 41567 13521
rect 41509 13481 41521 13515
rect 41555 13512 41567 13515
rect 41690 13512 41696 13524
rect 41555 13484 41696 13512
rect 41555 13481 41567 13484
rect 41509 13475 41567 13481
rect 41690 13472 41696 13484
rect 41748 13512 41754 13524
rect 42334 13512 42340 13524
rect 41748 13484 42340 13512
rect 41748 13472 41754 13484
rect 42334 13472 42340 13484
rect 42392 13512 42398 13524
rect 42702 13512 42708 13524
rect 42392 13484 42708 13512
rect 42392 13472 42398 13484
rect 42702 13472 42708 13484
rect 42760 13472 42766 13524
rect 43165 13515 43223 13521
rect 43165 13481 43177 13515
rect 43211 13512 43223 13515
rect 44174 13512 44180 13524
rect 43211 13484 44180 13512
rect 43211 13481 43223 13484
rect 43165 13475 43223 13481
rect 44174 13472 44180 13484
rect 44232 13512 44238 13524
rect 45002 13512 45008 13524
rect 44232 13484 45008 13512
rect 44232 13472 44238 13484
rect 45002 13472 45008 13484
rect 45060 13472 45066 13524
rect 50154 13472 50160 13524
rect 50212 13472 50218 13524
rect 53837 13515 53895 13521
rect 53837 13481 53849 13515
rect 53883 13512 53895 13515
rect 53926 13512 53932 13524
rect 53883 13484 53932 13512
rect 53883 13481 53895 13484
rect 53837 13475 53895 13481
rect 53926 13472 53932 13484
rect 53984 13472 53990 13524
rect 18414 13444 18420 13456
rect 17788 13416 18420 13444
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 17460 13280 17693 13308
rect 17460 13268 17466 13280
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 17788 13240 17816 13416
rect 18414 13404 18420 13416
rect 18472 13444 18478 13456
rect 19426 13444 19432 13456
rect 18472 13416 19432 13444
rect 18472 13404 18478 13416
rect 19426 13404 19432 13416
rect 19484 13404 19490 13456
rect 21450 13404 21456 13456
rect 21508 13444 21514 13456
rect 25958 13444 25964 13456
rect 21508 13416 25964 13444
rect 21508 13404 21514 13416
rect 19242 13336 19248 13388
rect 19300 13376 19306 13388
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 19300 13348 19901 13376
rect 19300 13336 19306 13348
rect 19889 13345 19901 13348
rect 19935 13345 19947 13379
rect 19889 13339 19947 13345
rect 23474 13336 23480 13388
rect 23532 13376 23538 13388
rect 23532 13348 23612 13376
rect 23532 13336 23538 13348
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18049 13311 18107 13317
rect 18049 13308 18061 13311
rect 18012 13280 18061 13308
rect 18012 13268 18018 13280
rect 18049 13277 18061 13280
rect 18095 13308 18107 13311
rect 18095 13280 18552 13308
rect 18095 13277 18107 13280
rect 18049 13271 18107 13277
rect 17236 13212 17816 13240
rect 18414 13200 18420 13252
rect 18472 13200 18478 13252
rect 18524 13240 18552 13280
rect 18782 13268 18788 13320
rect 18840 13308 18846 13320
rect 19337 13311 19395 13317
rect 19337 13308 19349 13311
rect 18840 13280 19349 13308
rect 18840 13268 18846 13280
rect 19337 13277 19349 13280
rect 19383 13277 19395 13311
rect 19337 13271 19395 13277
rect 19702 13268 19708 13320
rect 19760 13268 19766 13320
rect 23290 13268 23296 13320
rect 23348 13308 23354 13320
rect 23584 13317 23612 13348
rect 23768 13317 23796 13416
rect 25958 13404 25964 13416
rect 26016 13404 26022 13456
rect 26142 13404 26148 13456
rect 26200 13444 26206 13456
rect 26200 13416 27384 13444
rect 26200 13404 26206 13416
rect 24118 13336 24124 13388
rect 24176 13376 24182 13388
rect 24302 13376 24308 13388
rect 24176 13348 24308 13376
rect 24176 13336 24182 13348
rect 24302 13336 24308 13348
rect 24360 13376 24366 13388
rect 26605 13379 26663 13385
rect 26605 13376 26617 13379
rect 24360 13348 26617 13376
rect 24360 13336 24366 13348
rect 26605 13345 26617 13348
rect 26651 13345 26663 13379
rect 26605 13339 26663 13345
rect 26694 13336 26700 13388
rect 26752 13336 26758 13388
rect 26786 13336 26792 13388
rect 26844 13336 26850 13388
rect 26881 13379 26939 13385
rect 26881 13345 26893 13379
rect 26927 13376 26939 13379
rect 27154 13376 27160 13388
rect 26927 13348 27160 13376
rect 26927 13345 26939 13348
rect 26881 13339 26939 13345
rect 27154 13336 27160 13348
rect 27212 13336 27218 13388
rect 27356 13317 27384 13416
rect 32582 13404 32588 13456
rect 32640 13444 32646 13456
rect 32640 13416 35940 13444
rect 32640 13404 32646 13416
rect 27522 13336 27528 13388
rect 27580 13376 27586 13388
rect 27580 13348 28304 13376
rect 27580 13336 27586 13348
rect 23385 13311 23443 13317
rect 23385 13308 23397 13311
rect 23348 13280 23397 13308
rect 23348 13268 23354 13280
rect 23385 13277 23397 13280
rect 23431 13277 23443 13311
rect 23385 13271 23443 13277
rect 23569 13311 23627 13317
rect 23569 13277 23581 13311
rect 23615 13277 23627 13311
rect 23569 13271 23627 13277
rect 23753 13311 23811 13317
rect 23753 13277 23765 13311
rect 23799 13277 23811 13311
rect 23753 13271 23811 13277
rect 27341 13311 27399 13317
rect 27341 13277 27353 13311
rect 27387 13277 27399 13311
rect 27341 13271 27399 13277
rect 27706 13268 27712 13320
rect 27764 13308 27770 13320
rect 28276 13317 28304 13348
rect 28350 13336 28356 13388
rect 28408 13376 28414 13388
rect 30193 13379 30251 13385
rect 30193 13376 30205 13379
rect 28408 13348 30205 13376
rect 28408 13336 28414 13348
rect 30193 13345 30205 13348
rect 30239 13345 30251 13379
rect 30193 13339 30251 13345
rect 30285 13379 30343 13385
rect 30285 13345 30297 13379
rect 30331 13376 30343 13379
rect 30331 13348 31754 13376
rect 30331 13345 30343 13348
rect 30285 13339 30343 13345
rect 28077 13311 28135 13317
rect 28077 13308 28089 13311
rect 27764 13280 28089 13308
rect 27764 13268 27770 13280
rect 28077 13277 28089 13280
rect 28123 13277 28135 13311
rect 28077 13271 28135 13277
rect 28261 13311 28319 13317
rect 28261 13277 28273 13311
rect 28307 13277 28319 13311
rect 28261 13271 28319 13277
rect 28445 13311 28503 13317
rect 28445 13277 28457 13311
rect 28491 13277 28503 13311
rect 28445 13271 28503 13277
rect 18617 13243 18675 13249
rect 18617 13240 18629 13243
rect 18524 13212 18629 13240
rect 18617 13209 18629 13212
rect 18663 13209 18675 13243
rect 19794 13240 19800 13252
rect 18617 13203 18675 13209
rect 18708 13212 19800 13240
rect 8803 13144 9352 13172
rect 10781 13175 10839 13181
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 10781 13141 10793 13175
rect 10827 13172 10839 13175
rect 13814 13172 13820 13184
rect 10827 13144 13820 13172
rect 10827 13141 10839 13144
rect 10781 13135 10839 13141
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 18138 13132 18144 13184
rect 18196 13172 18202 13184
rect 18708 13172 18736 13212
rect 19794 13200 19800 13212
rect 19852 13200 19858 13252
rect 21361 13243 21419 13249
rect 21361 13209 21373 13243
rect 21407 13240 21419 13243
rect 22370 13240 22376 13252
rect 21407 13212 22376 13240
rect 21407 13209 21419 13212
rect 21361 13203 21419 13209
rect 22370 13200 22376 13212
rect 22428 13200 22434 13252
rect 23477 13243 23535 13249
rect 23477 13209 23489 13243
rect 23523 13209 23535 13243
rect 23477 13203 23535 13209
rect 18196 13144 18736 13172
rect 18785 13175 18843 13181
rect 18196 13132 18202 13144
rect 18785 13141 18797 13175
rect 18831 13172 18843 13175
rect 19058 13172 19064 13184
rect 18831 13144 19064 13172
rect 18831 13141 18843 13144
rect 18785 13135 18843 13141
rect 19058 13132 19064 13144
rect 19116 13132 19122 13184
rect 19429 13175 19487 13181
rect 19429 13141 19441 13175
rect 19475 13172 19487 13175
rect 20714 13172 20720 13184
rect 19475 13144 20720 13172
rect 19475 13141 19487 13144
rect 19429 13135 19487 13141
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 21450 13132 21456 13184
rect 21508 13172 21514 13184
rect 21566 13175 21624 13181
rect 21566 13172 21578 13175
rect 21508 13144 21578 13172
rect 21508 13132 21514 13144
rect 21566 13141 21578 13144
rect 21612 13141 21624 13175
rect 23492 13172 23520 13203
rect 25038 13200 25044 13252
rect 25096 13240 25102 13252
rect 27798 13240 27804 13252
rect 25096 13212 27804 13240
rect 25096 13200 25102 13212
rect 27798 13200 27804 13212
rect 27856 13200 27862 13252
rect 27890 13200 27896 13252
rect 27948 13240 27954 13252
rect 27985 13243 28043 13249
rect 27985 13240 27997 13243
rect 27948 13212 27997 13240
rect 27948 13200 27954 13212
rect 27985 13209 27997 13212
rect 28031 13209 28043 13243
rect 27985 13203 28043 13209
rect 23937 13175 23995 13181
rect 23937 13172 23949 13175
rect 23492 13144 23949 13172
rect 21566 13135 21624 13141
rect 23937 13141 23949 13144
rect 23983 13172 23995 13175
rect 24394 13172 24400 13184
rect 23983 13144 24400 13172
rect 23983 13141 23995 13144
rect 23937 13135 23995 13141
rect 24394 13132 24400 13144
rect 24452 13132 24458 13184
rect 26421 13175 26479 13181
rect 26421 13141 26433 13175
rect 26467 13172 26479 13175
rect 26786 13172 26792 13184
rect 26467 13144 26792 13172
rect 26467 13141 26479 13144
rect 26421 13135 26479 13141
rect 26786 13132 26792 13144
rect 26844 13132 26850 13184
rect 28276 13172 28304 13271
rect 28350 13200 28356 13252
rect 28408 13240 28414 13252
rect 28460 13240 28488 13271
rect 28718 13268 28724 13320
rect 28776 13268 28782 13320
rect 29089 13311 29147 13317
rect 29089 13308 29101 13311
rect 28828 13280 29101 13308
rect 28828 13240 28856 13280
rect 29089 13277 29101 13280
rect 29135 13277 29147 13311
rect 29089 13271 29147 13277
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13277 30159 13311
rect 30101 13271 30159 13277
rect 28408 13212 28856 13240
rect 28905 13243 28963 13249
rect 28408 13200 28414 13212
rect 28905 13209 28917 13243
rect 28951 13209 28963 13243
rect 30116 13240 30144 13271
rect 30374 13268 30380 13320
rect 30432 13268 30438 13320
rect 31726 13308 31754 13348
rect 34146 13336 34152 13388
rect 34204 13376 34210 13388
rect 35253 13379 35311 13385
rect 35253 13376 35265 13379
rect 34204 13348 35265 13376
rect 34204 13336 34210 13348
rect 35253 13345 35265 13348
rect 35299 13345 35311 13379
rect 35253 13339 35311 13345
rect 31938 13308 31944 13320
rect 31726 13280 31944 13308
rect 31938 13268 31944 13280
rect 31996 13268 32002 13320
rect 35069 13311 35127 13317
rect 35069 13277 35081 13311
rect 35115 13277 35127 13311
rect 35069 13271 35127 13277
rect 35345 13311 35403 13317
rect 35345 13277 35357 13311
rect 35391 13308 35403 13311
rect 35805 13311 35863 13317
rect 35805 13308 35817 13311
rect 35391 13280 35817 13308
rect 35391 13277 35403 13280
rect 35345 13271 35403 13277
rect 35805 13277 35817 13280
rect 35851 13277 35863 13311
rect 35805 13271 35863 13277
rect 30282 13240 30288 13252
rect 30116 13212 30288 13240
rect 28905 13203 28963 13209
rect 28920 13172 28948 13203
rect 30282 13200 30288 13212
rect 30340 13200 30346 13252
rect 32401 13243 32459 13249
rect 32401 13209 32413 13243
rect 32447 13209 32459 13243
rect 35084 13240 35112 13271
rect 35434 13240 35440 13252
rect 35084 13212 35440 13240
rect 32401 13203 32459 13209
rect 28276 13144 28948 13172
rect 31938 13132 31944 13184
rect 31996 13172 32002 13184
rect 32125 13175 32183 13181
rect 32125 13172 32137 13175
rect 31996 13144 32137 13172
rect 31996 13132 32002 13144
rect 32125 13141 32137 13144
rect 32171 13172 32183 13175
rect 32416 13172 32444 13203
rect 35434 13200 35440 13212
rect 35492 13200 35498 13252
rect 35912 13240 35940 13416
rect 36814 13404 36820 13456
rect 36872 13444 36878 13456
rect 37185 13447 37243 13453
rect 37185 13444 37197 13447
rect 36872 13416 37197 13444
rect 36872 13404 36878 13416
rect 37185 13413 37197 13416
rect 37231 13413 37243 13447
rect 37553 13447 37611 13453
rect 37553 13444 37565 13447
rect 37185 13407 37243 13413
rect 37384 13416 37565 13444
rect 37384 13376 37412 13416
rect 37553 13413 37565 13416
rect 37599 13413 37611 13447
rect 37553 13407 37611 13413
rect 38749 13447 38807 13453
rect 38749 13413 38761 13447
rect 38795 13444 38807 13447
rect 39503 13447 39561 13453
rect 39503 13444 39515 13447
rect 38795 13416 39515 13444
rect 38795 13413 38807 13416
rect 38749 13407 38807 13413
rect 39503 13413 39515 13416
rect 39549 13413 39561 13447
rect 39503 13407 39561 13413
rect 39758 13404 39764 13456
rect 39816 13444 39822 13456
rect 40034 13444 40040 13456
rect 39816 13416 40040 13444
rect 39816 13404 39822 13416
rect 40034 13404 40040 13416
rect 40092 13444 40098 13456
rect 40770 13444 40776 13456
rect 40092 13416 40776 13444
rect 40092 13404 40098 13416
rect 40770 13404 40776 13416
rect 40828 13404 40834 13456
rect 42518 13404 42524 13456
rect 42576 13444 42582 13456
rect 43533 13447 43591 13453
rect 43533 13444 43545 13447
rect 42576 13416 43545 13444
rect 42576 13404 42582 13416
rect 43533 13413 43545 13416
rect 43579 13444 43591 13447
rect 44542 13444 44548 13456
rect 43579 13416 44548 13444
rect 43579 13413 43591 13416
rect 43533 13407 43591 13413
rect 44542 13404 44548 13416
rect 44600 13404 44606 13456
rect 44634 13404 44640 13456
rect 44692 13444 44698 13456
rect 50617 13447 50675 13453
rect 44692 13416 45513 13444
rect 44692 13404 44698 13416
rect 36740 13348 37412 13376
rect 37461 13379 37519 13385
rect 36740 13320 36768 13348
rect 37461 13345 37473 13379
rect 37507 13376 37519 13379
rect 39301 13379 39359 13385
rect 39301 13376 39313 13379
rect 37507 13348 39313 13376
rect 37507 13345 37519 13348
rect 37461 13339 37519 13345
rect 39301 13345 39313 13348
rect 39347 13345 39359 13379
rect 40957 13379 41015 13385
rect 40957 13376 40969 13379
rect 39301 13339 39359 13345
rect 39684 13348 40969 13376
rect 36354 13268 36360 13320
rect 36412 13268 36418 13320
rect 36722 13268 36728 13320
rect 36780 13268 36786 13320
rect 36998 13268 37004 13320
rect 37056 13268 37062 13320
rect 37826 13268 37832 13320
rect 37884 13308 37890 13320
rect 38105 13311 38163 13317
rect 38105 13308 38117 13311
rect 37884 13280 38117 13308
rect 37884 13268 37890 13280
rect 38105 13277 38117 13280
rect 38151 13277 38163 13311
rect 38105 13271 38163 13277
rect 38194 13268 38200 13320
rect 38252 13308 38258 13320
rect 38252 13280 38297 13308
rect 38252 13268 38258 13280
rect 38378 13268 38384 13320
rect 38436 13268 38442 13320
rect 38570 13311 38628 13317
rect 38570 13277 38582 13311
rect 38616 13277 38628 13311
rect 38570 13271 38628 13277
rect 35912 13212 36952 13240
rect 32171 13144 32444 13172
rect 32171 13141 32183 13144
rect 32125 13135 32183 13141
rect 34698 13132 34704 13184
rect 34756 13172 34762 13184
rect 34885 13175 34943 13181
rect 34885 13172 34897 13175
rect 34756 13144 34897 13172
rect 34756 13132 34762 13144
rect 34885 13141 34897 13144
rect 34931 13141 34943 13175
rect 34885 13135 34943 13141
rect 36538 13132 36544 13184
rect 36596 13172 36602 13184
rect 36817 13175 36875 13181
rect 36817 13172 36829 13175
rect 36596 13144 36829 13172
rect 36596 13132 36602 13144
rect 36817 13141 36829 13144
rect 36863 13141 36875 13175
rect 36924 13172 36952 13212
rect 37090 13200 37096 13252
rect 37148 13240 37154 13252
rect 38010 13240 38016 13252
rect 37148 13212 38016 13240
rect 37148 13200 37154 13212
rect 38010 13200 38016 13212
rect 38068 13200 38074 13252
rect 38473 13243 38531 13249
rect 38473 13240 38485 13243
rect 38120 13212 38485 13240
rect 38120 13172 38148 13212
rect 38473 13209 38485 13212
rect 38519 13209 38531 13243
rect 38473 13203 38531 13209
rect 36924 13144 38148 13172
rect 36817 13135 36875 13141
rect 38286 13132 38292 13184
rect 38344 13172 38350 13184
rect 38580 13172 38608 13271
rect 39114 13268 39120 13320
rect 39172 13268 39178 13320
rect 39684 13317 39712 13348
rect 40957 13345 40969 13348
rect 41003 13345 41015 13379
rect 40957 13339 41015 13345
rect 41325 13379 41383 13385
rect 41325 13345 41337 13379
rect 41371 13376 41383 13379
rect 41506 13376 41512 13388
rect 41371 13348 41512 13376
rect 41371 13345 41383 13348
rect 41325 13339 41383 13345
rect 41506 13336 41512 13348
rect 41564 13376 41570 13388
rect 45485 13376 45513 13416
rect 50617 13413 50629 13447
rect 50663 13444 50675 13447
rect 51166 13444 51172 13456
rect 50663 13416 51172 13444
rect 50663 13413 50675 13416
rect 50617 13407 50675 13413
rect 51166 13404 51172 13416
rect 51224 13404 51230 13456
rect 52362 13404 52368 13456
rect 52420 13444 52426 13456
rect 54205 13447 54263 13453
rect 54205 13444 54217 13447
rect 52420 13416 54217 13444
rect 52420 13404 52426 13416
rect 54205 13413 54217 13416
rect 54251 13413 54263 13447
rect 54205 13407 54263 13413
rect 48038 13376 48044 13388
rect 41564 13348 45232 13376
rect 41564 13336 41570 13348
rect 39669 13311 39727 13317
rect 39669 13277 39681 13311
rect 39715 13277 39727 13311
rect 39669 13271 39727 13277
rect 39850 13268 39856 13320
rect 39908 13268 39914 13320
rect 40034 13268 40040 13320
rect 40092 13268 40098 13320
rect 40221 13311 40279 13317
rect 40221 13277 40233 13311
rect 40267 13308 40279 13311
rect 40494 13308 40500 13320
rect 40267 13280 40500 13308
rect 40267 13277 40279 13280
rect 40221 13271 40279 13277
rect 40494 13268 40500 13280
rect 40552 13308 40558 13320
rect 40770 13308 40776 13320
rect 40552 13280 40776 13308
rect 40552 13268 40558 13280
rect 40770 13268 40776 13280
rect 40828 13268 40834 13320
rect 41141 13311 41199 13317
rect 41141 13277 41153 13311
rect 41187 13308 41199 13311
rect 41690 13308 41696 13320
rect 41187 13280 41696 13308
rect 41187 13277 41199 13280
rect 41141 13271 41199 13277
rect 41690 13268 41696 13280
rect 41748 13268 41754 13320
rect 42886 13268 42892 13320
rect 42944 13308 42950 13320
rect 42981 13311 43039 13317
rect 42981 13308 42993 13311
rect 42944 13280 42993 13308
rect 42944 13268 42950 13280
rect 42981 13277 42993 13280
rect 43027 13277 43039 13311
rect 42981 13271 43039 13277
rect 43257 13311 43315 13317
rect 43257 13277 43269 13311
rect 43303 13308 43315 13311
rect 43901 13311 43959 13317
rect 43901 13308 43913 13311
rect 43303 13280 43913 13308
rect 43303 13277 43315 13280
rect 43257 13271 43315 13277
rect 43901 13277 43913 13280
rect 43947 13277 43959 13311
rect 43901 13271 43959 13277
rect 44450 13268 44456 13320
rect 44508 13268 44514 13320
rect 44910 13268 44916 13320
rect 44968 13308 44974 13320
rect 45005 13311 45063 13317
rect 45005 13308 45017 13311
rect 44968 13280 45017 13308
rect 44968 13268 44974 13280
rect 45005 13277 45017 13280
rect 45051 13277 45063 13311
rect 45005 13271 45063 13277
rect 45098 13311 45156 13317
rect 45098 13277 45110 13311
rect 45144 13277 45156 13311
rect 45098 13271 45156 13277
rect 40126 13200 40132 13252
rect 40184 13200 40190 13252
rect 43717 13243 43775 13249
rect 43717 13209 43729 13243
rect 43763 13209 43775 13243
rect 44468 13240 44496 13268
rect 45112 13240 45140 13271
rect 44468 13212 45140 13240
rect 45204 13240 45232 13348
rect 45485 13348 48044 13376
rect 45278 13268 45284 13320
rect 45336 13268 45342 13320
rect 45485 13317 45513 13348
rect 48038 13336 48044 13348
rect 48096 13336 48102 13388
rect 50246 13336 50252 13388
rect 50304 13376 50310 13388
rect 50304 13348 50476 13376
rect 50304 13336 50310 13348
rect 45470 13311 45528 13317
rect 45470 13277 45482 13311
rect 45516 13277 45528 13311
rect 45470 13271 45528 13277
rect 47762 13268 47768 13320
rect 47820 13308 47826 13320
rect 50448 13317 50476 13348
rect 53834 13336 53840 13388
rect 53892 13376 53898 13388
rect 54297 13379 54355 13385
rect 54297 13376 54309 13379
rect 53892 13348 54309 13376
rect 53892 13336 53898 13348
rect 54297 13345 54309 13348
rect 54343 13376 54355 13379
rect 55398 13376 55404 13388
rect 54343 13348 55404 13376
rect 54343 13345 54355 13348
rect 54297 13339 54355 13345
rect 55398 13336 55404 13348
rect 55456 13336 55462 13388
rect 50341 13311 50399 13317
rect 50341 13308 50353 13311
rect 47820 13280 50353 13308
rect 47820 13268 47826 13280
rect 50341 13277 50353 13280
rect 50387 13277 50399 13311
rect 50341 13271 50399 13277
rect 50433 13311 50491 13317
rect 50433 13277 50445 13311
rect 50479 13277 50491 13311
rect 50433 13271 50491 13277
rect 50614 13268 50620 13320
rect 50672 13308 50678 13320
rect 50709 13311 50767 13317
rect 50709 13308 50721 13311
rect 50672 13280 50721 13308
rect 50672 13268 50678 13280
rect 50709 13277 50721 13280
rect 50755 13277 50767 13311
rect 50709 13271 50767 13277
rect 54021 13311 54079 13317
rect 54021 13277 54033 13311
rect 54067 13308 54079 13311
rect 54110 13308 54116 13320
rect 54067 13280 54116 13308
rect 54067 13277 54079 13280
rect 54021 13271 54079 13277
rect 54110 13268 54116 13280
rect 54168 13268 54174 13320
rect 45370 13240 45376 13252
rect 45204 13212 45376 13240
rect 43717 13203 43775 13209
rect 38344 13144 38608 13172
rect 39117 13175 39175 13181
rect 38344 13132 38350 13144
rect 39117 13141 39129 13175
rect 39163 13172 39175 13175
rect 40402 13172 40408 13184
rect 39163 13144 40408 13172
rect 39163 13141 39175 13144
rect 39117 13135 39175 13141
rect 40402 13132 40408 13144
rect 40460 13132 40466 13184
rect 42797 13175 42855 13181
rect 42797 13141 42809 13175
rect 42843 13172 42855 13175
rect 42978 13172 42984 13184
rect 42843 13144 42984 13172
rect 42843 13141 42855 13144
rect 42797 13135 42855 13141
rect 42978 13132 42984 13144
rect 43036 13132 43042 13184
rect 43732 13172 43760 13203
rect 45370 13200 45376 13212
rect 45428 13200 45434 13252
rect 44634 13172 44640 13184
rect 43732 13144 44640 13172
rect 44634 13132 44640 13144
rect 44692 13132 44698 13184
rect 45554 13132 45560 13184
rect 45612 13172 45618 13184
rect 45649 13175 45707 13181
rect 45649 13172 45661 13175
rect 45612 13144 45661 13172
rect 45612 13132 45618 13144
rect 45649 13141 45661 13144
rect 45695 13141 45707 13175
rect 45649 13135 45707 13141
rect 1104 13082 78844 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 66314 13082
rect 66366 13030 66378 13082
rect 66430 13030 66442 13082
rect 66494 13030 66506 13082
rect 66558 13030 66570 13082
rect 66622 13030 78844 13082
rect 1104 13008 78844 13030
rect 13814 12928 13820 12980
rect 13872 12928 13878 12980
rect 14458 12928 14464 12980
rect 14516 12968 14522 12980
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 14516 12940 15025 12968
rect 14516 12928 14522 12940
rect 15013 12937 15025 12940
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 18414 12928 18420 12980
rect 18472 12968 18478 12980
rect 19150 12968 19156 12980
rect 18472 12940 19156 12968
rect 18472 12928 18478 12940
rect 19150 12928 19156 12940
rect 19208 12968 19214 12980
rect 19208 12940 19840 12968
rect 19208 12928 19214 12940
rect 13832 12900 13860 12928
rect 18506 12900 18512 12912
rect 13832 12872 18512 12900
rect 15396 12841 15424 12872
rect 18506 12860 18512 12872
rect 18564 12860 18570 12912
rect 19613 12903 19671 12909
rect 19613 12900 19625 12903
rect 18616 12872 19625 12900
rect 13909 12835 13967 12841
rect 13909 12801 13921 12835
rect 13955 12832 13967 12835
rect 14277 12835 14335 12841
rect 14277 12832 14289 12835
rect 13955 12804 14289 12832
rect 13955 12801 13967 12804
rect 13909 12795 13967 12801
rect 14277 12801 14289 12804
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 17129 12835 17187 12841
rect 17129 12801 17141 12835
rect 17175 12832 17187 12835
rect 17310 12832 17316 12844
rect 17175 12804 17316 12832
rect 17175 12801 17187 12804
rect 17129 12795 17187 12801
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 18325 12835 18383 12841
rect 18325 12801 18337 12835
rect 18371 12832 18383 12835
rect 18414 12832 18420 12844
rect 18371 12804 18420 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 18616 12841 18644 12872
rect 19613 12869 19625 12872
rect 19659 12869 19671 12903
rect 19812 12900 19840 12940
rect 22186 12928 22192 12980
rect 22244 12968 22250 12980
rect 22370 12968 22376 12980
rect 22244 12940 22376 12968
rect 22244 12928 22250 12940
rect 22370 12928 22376 12940
rect 22428 12928 22434 12980
rect 22465 12971 22523 12977
rect 22465 12937 22477 12971
rect 22511 12968 22523 12971
rect 23934 12968 23940 12980
rect 22511 12940 23940 12968
rect 22511 12937 22523 12940
rect 22465 12931 22523 12937
rect 23934 12928 23940 12940
rect 23992 12968 23998 12980
rect 25038 12968 25044 12980
rect 23992 12940 25044 12968
rect 23992 12928 23998 12940
rect 25038 12928 25044 12940
rect 25096 12968 25102 12980
rect 25498 12968 25504 12980
rect 25096 12940 25504 12968
rect 25096 12928 25102 12940
rect 25498 12928 25504 12940
rect 25556 12928 25562 12980
rect 27890 12928 27896 12980
rect 27948 12968 27954 12980
rect 28534 12968 28540 12980
rect 27948 12940 28540 12968
rect 27948 12928 27954 12940
rect 28534 12928 28540 12940
rect 28592 12928 28598 12980
rect 31662 12968 31668 12980
rect 31036 12940 31668 12968
rect 19812 12872 19932 12900
rect 19613 12863 19671 12869
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 18782 12792 18788 12844
rect 18840 12792 18846 12844
rect 18874 12792 18880 12844
rect 18932 12792 18938 12844
rect 19058 12792 19064 12844
rect 19116 12792 19122 12844
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12832 19395 12835
rect 19383 12804 19748 12832
rect 19383 12801 19395 12804
rect 19337 12795 19395 12801
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12733 14151 12767
rect 14093 12727 14151 12733
rect 14108 12696 14136 12727
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14884 12736 14933 12764
rect 14884 12724 14890 12736
rect 14921 12733 14933 12736
rect 14967 12764 14979 12767
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 14967 12736 15301 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 15289 12733 15301 12736
rect 15335 12733 15347 12767
rect 15289 12727 15347 12733
rect 16942 12724 16948 12776
rect 17000 12764 17006 12776
rect 17865 12767 17923 12773
rect 17865 12764 17877 12767
rect 17000 12736 17877 12764
rect 17000 12724 17006 12736
rect 17865 12733 17877 12736
rect 17911 12733 17923 12767
rect 18800 12764 18828 12792
rect 17865 12727 17923 12733
rect 18248 12736 18828 12764
rect 19521 12767 19579 12773
rect 15010 12696 15016 12708
rect 14108 12668 15016 12696
rect 15010 12656 15016 12668
rect 15068 12696 15074 12708
rect 16390 12696 16396 12708
rect 15068 12668 16396 12696
rect 15068 12656 15074 12668
rect 16390 12656 16396 12668
rect 16448 12656 16454 12708
rect 17880 12696 17908 12727
rect 18248 12696 18276 12736
rect 19521 12733 19533 12767
rect 19567 12733 19579 12767
rect 19720 12764 19748 12804
rect 19794 12792 19800 12844
rect 19852 12792 19858 12844
rect 19904 12841 19932 12872
rect 21450 12860 21456 12912
rect 21508 12900 21514 12912
rect 22097 12903 22155 12909
rect 22097 12900 22109 12903
rect 21508 12872 22109 12900
rect 21508 12860 21514 12872
rect 22097 12869 22109 12872
rect 22143 12869 22155 12903
rect 26694 12900 26700 12912
rect 22097 12863 22155 12869
rect 25516 12872 26700 12900
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12801 19947 12835
rect 19889 12795 19947 12801
rect 20070 12792 20076 12844
rect 20128 12792 20134 12844
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12832 20867 12835
rect 21542 12832 21548 12844
rect 20855 12804 21548 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 20824 12764 20852 12795
rect 21542 12792 21548 12804
rect 21600 12832 21606 12844
rect 22306 12835 22364 12841
rect 22306 12832 22318 12835
rect 21600 12804 22318 12832
rect 21600 12792 21606 12804
rect 22306 12801 22318 12804
rect 22352 12801 22364 12835
rect 22306 12795 22364 12801
rect 25222 12792 25228 12844
rect 25280 12832 25286 12844
rect 25516 12841 25544 12872
rect 26694 12860 26700 12872
rect 26752 12860 26758 12912
rect 31036 12909 31064 12940
rect 31662 12928 31668 12940
rect 31720 12928 31726 12980
rect 32306 12968 32312 12980
rect 31772 12940 32312 12968
rect 31021 12903 31079 12909
rect 31021 12869 31033 12903
rect 31067 12869 31079 12903
rect 31021 12863 31079 12869
rect 31237 12903 31295 12909
rect 31237 12869 31249 12903
rect 31283 12900 31295 12903
rect 31772 12900 31800 12940
rect 32306 12928 32312 12940
rect 32364 12928 32370 12980
rect 33229 12971 33287 12977
rect 33229 12937 33241 12971
rect 33275 12968 33287 12971
rect 33318 12968 33324 12980
rect 33275 12940 33324 12968
rect 33275 12937 33287 12940
rect 33229 12931 33287 12937
rect 33318 12928 33324 12940
rect 33376 12928 33382 12980
rect 36265 12971 36323 12977
rect 36265 12968 36277 12971
rect 35085 12940 36277 12968
rect 31283 12872 31800 12900
rect 31849 12903 31907 12909
rect 31283 12869 31295 12872
rect 31237 12863 31295 12869
rect 31849 12869 31861 12903
rect 31895 12900 31907 12903
rect 32401 12903 32459 12909
rect 32401 12900 32413 12903
rect 31895 12872 32413 12900
rect 31895 12869 31907 12872
rect 31849 12863 31907 12869
rect 32401 12869 32413 12872
rect 32447 12869 32459 12903
rect 32401 12863 32459 12869
rect 33336 12900 33364 12928
rect 33870 12900 33876 12912
rect 33336 12872 33876 12900
rect 25409 12835 25467 12841
rect 25409 12832 25421 12835
rect 25280 12804 25421 12832
rect 25280 12792 25286 12804
rect 25409 12801 25421 12804
rect 25455 12801 25467 12835
rect 25409 12795 25467 12801
rect 25501 12835 25559 12841
rect 25501 12801 25513 12835
rect 25547 12801 25559 12835
rect 25501 12795 25559 12801
rect 19720 12736 20852 12764
rect 21821 12767 21879 12773
rect 19521 12727 19579 12733
rect 21821 12733 21833 12767
rect 21867 12733 21879 12767
rect 21821 12727 21879 12733
rect 17880 12668 18276 12696
rect 18509 12699 18567 12705
rect 18509 12665 18521 12699
rect 18555 12696 18567 12699
rect 19334 12696 19340 12708
rect 18555 12668 19340 12696
rect 18555 12665 18567 12668
rect 18509 12659 18567 12665
rect 19334 12656 19340 12668
rect 19392 12656 19398 12708
rect 19536 12696 19564 12727
rect 20165 12699 20223 12705
rect 20165 12696 20177 12699
rect 19536 12668 20177 12696
rect 20165 12665 20177 12668
rect 20211 12665 20223 12699
rect 20165 12659 20223 12665
rect 20714 12656 20720 12708
rect 20772 12696 20778 12708
rect 21836 12696 21864 12727
rect 23934 12724 23940 12776
rect 23992 12764 23998 12776
rect 25516 12764 25544 12795
rect 25682 12792 25688 12844
rect 25740 12792 25746 12844
rect 25774 12792 25780 12844
rect 25832 12792 25838 12844
rect 31665 12835 31723 12841
rect 31665 12832 31677 12835
rect 31404 12804 31677 12832
rect 23992 12736 25544 12764
rect 23992 12724 23998 12736
rect 20772 12668 21864 12696
rect 20772 12656 20778 12668
rect 26970 12656 26976 12708
rect 27028 12696 27034 12708
rect 27890 12696 27896 12708
rect 27028 12668 27896 12696
rect 27028 12656 27034 12668
rect 27890 12656 27896 12668
rect 27948 12656 27954 12708
rect 31404 12705 31432 12804
rect 31665 12801 31677 12804
rect 31711 12801 31723 12835
rect 31665 12795 31723 12801
rect 31941 12835 31999 12841
rect 31941 12801 31953 12835
rect 31987 12832 31999 12835
rect 32030 12832 32036 12844
rect 31987 12804 32036 12832
rect 31987 12801 31999 12804
rect 31941 12795 31999 12801
rect 32030 12792 32036 12804
rect 32088 12832 32094 12844
rect 32766 12832 32772 12844
rect 32088 12804 32772 12832
rect 32088 12792 32094 12804
rect 32766 12792 32772 12804
rect 32824 12792 32830 12844
rect 33336 12841 33364 12872
rect 33870 12860 33876 12872
rect 33928 12860 33934 12912
rect 34698 12860 34704 12912
rect 34756 12860 34762 12912
rect 34790 12860 34796 12912
rect 34848 12900 34854 12912
rect 35085 12900 35113 12940
rect 36265 12937 36277 12940
rect 36311 12937 36323 12971
rect 36265 12931 36323 12937
rect 36906 12928 36912 12980
rect 36964 12928 36970 12980
rect 36998 12928 37004 12980
rect 37056 12968 37062 12980
rect 37093 12971 37151 12977
rect 37093 12968 37105 12971
rect 37056 12940 37105 12968
rect 37056 12928 37062 12940
rect 37093 12937 37105 12940
rect 37139 12937 37151 12971
rect 37093 12931 37151 12937
rect 37826 12928 37832 12980
rect 37884 12928 37890 12980
rect 37918 12928 37924 12980
rect 37976 12968 37982 12980
rect 38286 12968 38292 12980
rect 37976 12940 38292 12968
rect 37976 12928 37982 12940
rect 38286 12928 38292 12940
rect 38344 12968 38350 12980
rect 38841 12971 38899 12977
rect 38841 12968 38853 12971
rect 38344 12940 38853 12968
rect 38344 12928 38350 12940
rect 38841 12937 38853 12940
rect 38887 12937 38899 12971
rect 45094 12968 45100 12980
rect 38841 12931 38899 12937
rect 42720 12940 45100 12968
rect 34848 12872 35190 12900
rect 34848 12860 34854 12872
rect 36354 12860 36360 12912
rect 36412 12900 36418 12912
rect 36924 12900 36952 12928
rect 36412 12872 37320 12900
rect 36412 12860 36418 12872
rect 33321 12835 33379 12841
rect 33321 12801 33333 12835
rect 33367 12801 33379 12835
rect 33321 12795 33379 12801
rect 33594 12792 33600 12844
rect 33652 12792 33658 12844
rect 36633 12835 36691 12841
rect 36633 12801 36645 12835
rect 36679 12832 36691 12835
rect 36814 12832 36820 12844
rect 36679 12804 36820 12832
rect 36679 12801 36691 12804
rect 36633 12795 36691 12801
rect 36814 12792 36820 12804
rect 36872 12832 36878 12844
rect 36909 12835 36967 12841
rect 36909 12832 36921 12835
rect 36872 12804 36921 12832
rect 36872 12792 36878 12804
rect 36909 12801 36921 12804
rect 36955 12832 36967 12835
rect 37090 12832 37096 12844
rect 36955 12804 37096 12832
rect 36955 12801 36967 12804
rect 36909 12795 36967 12801
rect 37090 12792 37096 12804
rect 37148 12792 37154 12844
rect 37292 12841 37320 12872
rect 37458 12860 37464 12912
rect 37516 12860 37522 12912
rect 37553 12903 37611 12909
rect 37553 12869 37565 12903
rect 37599 12900 37611 12903
rect 37734 12900 37740 12912
rect 37599 12872 37740 12900
rect 37599 12869 37611 12872
rect 37553 12863 37611 12869
rect 37734 12860 37740 12872
rect 37792 12860 37798 12912
rect 38013 12903 38071 12909
rect 38013 12869 38025 12903
rect 38059 12900 38071 12903
rect 38102 12900 38108 12912
rect 38059 12872 38108 12900
rect 38059 12869 38071 12872
rect 38013 12863 38071 12869
rect 37277 12835 37335 12841
rect 37277 12801 37289 12835
rect 37323 12801 37335 12835
rect 37277 12795 37335 12801
rect 37642 12792 37648 12844
rect 37700 12832 37706 12844
rect 38028 12832 38056 12863
rect 38102 12860 38108 12872
rect 38160 12860 38166 12912
rect 40126 12860 40132 12912
rect 40184 12900 40190 12912
rect 40184 12872 42656 12900
rect 40184 12860 40190 12872
rect 37700 12804 38056 12832
rect 38197 12835 38255 12841
rect 37700 12792 37706 12804
rect 38197 12801 38209 12835
rect 38243 12832 38255 12835
rect 38286 12832 38292 12844
rect 38243 12804 38292 12832
rect 38243 12801 38255 12804
rect 38197 12795 38255 12801
rect 38286 12792 38292 12804
rect 38344 12792 38350 12844
rect 38562 12792 38568 12844
rect 38620 12832 38626 12844
rect 38620 12804 40080 12832
rect 38620 12792 38626 12804
rect 33045 12767 33103 12773
rect 33045 12733 33057 12767
rect 33091 12733 33103 12767
rect 33045 12727 33103 12733
rect 31389 12699 31447 12705
rect 31389 12665 31401 12699
rect 31435 12665 31447 12699
rect 31389 12659 31447 12665
rect 32858 12656 32864 12708
rect 32916 12696 32922 12708
rect 33060 12696 33088 12727
rect 34422 12724 34428 12776
rect 34480 12724 34486 12776
rect 36725 12767 36783 12773
rect 36725 12764 36737 12767
rect 34532 12736 36737 12764
rect 34532 12696 34560 12736
rect 36725 12733 36737 12736
rect 36771 12733 36783 12767
rect 39850 12764 39856 12776
rect 36725 12727 36783 12733
rect 36832 12736 39856 12764
rect 32916 12668 34560 12696
rect 32916 12656 32922 12668
rect 35710 12656 35716 12708
rect 35768 12696 35774 12708
rect 36832 12696 36860 12736
rect 39850 12724 39856 12736
rect 39908 12724 39914 12776
rect 40052 12764 40080 12804
rect 40586 12792 40592 12844
rect 40644 12792 40650 12844
rect 41414 12832 41420 12844
rect 40788 12804 41420 12832
rect 40788 12773 40816 12804
rect 41414 12792 41420 12804
rect 41472 12832 41478 12844
rect 42242 12832 42248 12844
rect 41472 12804 42248 12832
rect 41472 12792 41478 12804
rect 42242 12792 42248 12804
rect 42300 12792 42306 12844
rect 40773 12767 40831 12773
rect 40773 12764 40785 12767
rect 40052 12736 40785 12764
rect 40773 12733 40785 12736
rect 40819 12733 40831 12767
rect 40773 12727 40831 12733
rect 40865 12767 40923 12773
rect 40865 12733 40877 12767
rect 40911 12764 40923 12767
rect 41325 12767 41383 12773
rect 41325 12764 41337 12767
rect 40911 12736 41337 12764
rect 40911 12733 40923 12736
rect 40865 12727 40923 12733
rect 41325 12733 41337 12736
rect 41371 12733 41383 12767
rect 41325 12727 41383 12733
rect 41969 12767 42027 12773
rect 41969 12733 41981 12767
rect 42015 12764 42027 12767
rect 42150 12764 42156 12776
rect 42015 12736 42156 12764
rect 42015 12733 42027 12736
rect 41969 12727 42027 12733
rect 35768 12668 36860 12696
rect 35768 12656 35774 12668
rect 38194 12656 38200 12708
rect 38252 12696 38258 12708
rect 41984 12696 42012 12727
rect 42150 12724 42156 12736
rect 42208 12724 42214 12776
rect 42628 12764 42656 12872
rect 42720 12841 42748 12940
rect 45094 12928 45100 12940
rect 45152 12928 45158 12980
rect 42978 12860 42984 12912
rect 43036 12860 43042 12912
rect 44266 12900 44272 12912
rect 44206 12872 44272 12900
rect 44266 12860 44272 12872
rect 44324 12900 44330 12912
rect 45005 12903 45063 12909
rect 45005 12900 45017 12903
rect 44324 12872 45017 12900
rect 44324 12860 44330 12872
rect 45005 12869 45017 12872
rect 45051 12869 45063 12903
rect 46750 12900 46756 12912
rect 46598 12872 46756 12900
rect 45005 12863 45063 12869
rect 46750 12860 46756 12872
rect 46808 12860 46814 12912
rect 42705 12835 42763 12841
rect 42705 12801 42717 12835
rect 42751 12801 42763 12835
rect 42705 12795 42763 12801
rect 44542 12792 44548 12844
rect 44600 12832 44606 12844
rect 44637 12835 44695 12841
rect 44637 12832 44649 12835
rect 44600 12804 44649 12832
rect 44600 12792 44606 12804
rect 44637 12801 44649 12804
rect 44683 12801 44695 12835
rect 44637 12795 44695 12801
rect 45094 12792 45100 12844
rect 45152 12792 45158 12844
rect 50338 12792 50344 12844
rect 50396 12832 50402 12844
rect 50801 12835 50859 12841
rect 50801 12832 50813 12835
rect 50396 12804 50813 12832
rect 50396 12792 50402 12804
rect 50801 12801 50813 12804
rect 50847 12832 50859 12835
rect 51169 12835 51227 12841
rect 51169 12832 51181 12835
rect 50847 12804 51181 12832
rect 50847 12801 50859 12804
rect 50801 12795 50859 12801
rect 51169 12801 51181 12804
rect 51215 12832 51227 12835
rect 54478 12832 54484 12844
rect 51215 12804 54484 12832
rect 51215 12801 51227 12804
rect 51169 12795 51227 12801
rect 54478 12792 54484 12804
rect 54536 12792 54542 12844
rect 44450 12764 44456 12776
rect 42628 12736 44456 12764
rect 44450 12724 44456 12736
rect 44508 12724 44514 12776
rect 45370 12724 45376 12776
rect 45428 12724 45434 12776
rect 38252 12668 42012 12696
rect 38252 12656 38258 12668
rect 44266 12656 44272 12708
rect 44324 12696 44330 12708
rect 44910 12696 44916 12708
rect 44324 12668 44916 12696
rect 44324 12656 44330 12668
rect 44910 12656 44916 12668
rect 44968 12656 44974 12708
rect 12986 12588 12992 12640
rect 13044 12628 13050 12640
rect 13449 12631 13507 12637
rect 13449 12628 13461 12631
rect 13044 12600 13461 12628
rect 13044 12588 13050 12600
rect 13449 12597 13461 12600
rect 13495 12597 13507 12631
rect 13449 12591 13507 12597
rect 17678 12588 17684 12640
rect 17736 12588 17742 12640
rect 18414 12588 18420 12640
rect 18472 12628 18478 12640
rect 19242 12628 19248 12640
rect 18472 12600 19248 12628
rect 18472 12588 18478 12600
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 20901 12631 20959 12637
rect 20901 12597 20913 12631
rect 20947 12628 20959 12631
rect 21174 12628 21180 12640
rect 20947 12600 21180 12628
rect 20947 12597 20959 12600
rect 20901 12591 20959 12597
rect 21174 12588 21180 12600
rect 21232 12588 21238 12640
rect 25225 12631 25283 12637
rect 25225 12597 25237 12631
rect 25271 12628 25283 12631
rect 27338 12628 27344 12640
rect 25271 12600 27344 12628
rect 25271 12597 25283 12600
rect 25225 12591 25283 12597
rect 27338 12588 27344 12600
rect 27396 12588 27402 12640
rect 31018 12588 31024 12640
rect 31076 12628 31082 12640
rect 31205 12631 31263 12637
rect 31205 12628 31217 12631
rect 31076 12600 31217 12628
rect 31076 12588 31082 12600
rect 31205 12597 31217 12600
rect 31251 12597 31263 12631
rect 31205 12591 31263 12597
rect 31478 12588 31484 12640
rect 31536 12588 31542 12640
rect 33410 12588 33416 12640
rect 33468 12628 33474 12640
rect 36173 12631 36231 12637
rect 36173 12628 36185 12631
rect 33468 12600 36185 12628
rect 33468 12588 33474 12600
rect 36173 12597 36185 12600
rect 36219 12628 36231 12631
rect 36354 12628 36360 12640
rect 36219 12600 36360 12628
rect 36219 12597 36231 12600
rect 36173 12591 36231 12597
rect 36354 12588 36360 12600
rect 36412 12588 36418 12640
rect 40405 12631 40463 12637
rect 40405 12597 40417 12631
rect 40451 12628 40463 12631
rect 40678 12628 40684 12640
rect 40451 12600 40684 12628
rect 40451 12597 40463 12600
rect 40405 12591 40463 12597
rect 40678 12588 40684 12600
rect 40736 12588 40742 12640
rect 46842 12588 46848 12640
rect 46900 12588 46906 12640
rect 50982 12588 50988 12640
rect 51040 12588 51046 12640
rect 1104 12538 78844 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 78844 12538
rect 1104 12464 78844 12486
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 14185 12427 14243 12433
rect 14185 12424 14197 12427
rect 14056 12396 14197 12424
rect 14056 12384 14062 12396
rect 14185 12393 14197 12396
rect 14231 12393 14243 12427
rect 14185 12387 14243 12393
rect 16991 12427 17049 12433
rect 16991 12393 17003 12427
rect 17037 12424 17049 12427
rect 17310 12424 17316 12436
rect 17037 12396 17316 12424
rect 17037 12393 17049 12396
rect 16991 12387 17049 12393
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 19797 12427 19855 12433
rect 19797 12393 19809 12427
rect 19843 12424 19855 12427
rect 20070 12424 20076 12436
rect 19843 12396 20076 12424
rect 19843 12393 19855 12396
rect 19797 12387 19855 12393
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 23661 12427 23719 12433
rect 23661 12393 23673 12427
rect 23707 12424 23719 12427
rect 24210 12424 24216 12436
rect 23707 12396 24216 12424
rect 23707 12393 23719 12396
rect 23661 12387 23719 12393
rect 24210 12384 24216 12396
rect 24268 12384 24274 12436
rect 24302 12384 24308 12436
rect 24360 12424 24366 12436
rect 24489 12427 24547 12433
rect 24489 12424 24501 12427
rect 24360 12396 24501 12424
rect 24360 12384 24366 12396
rect 24489 12393 24501 12396
rect 24535 12393 24547 12427
rect 24489 12387 24547 12393
rect 25685 12427 25743 12433
rect 25685 12393 25697 12427
rect 25731 12424 25743 12427
rect 25774 12424 25780 12436
rect 25731 12396 25780 12424
rect 25731 12393 25743 12396
rect 25685 12387 25743 12393
rect 25774 12384 25780 12396
rect 25832 12384 25838 12436
rect 28534 12424 28540 12436
rect 26068 12396 28540 12424
rect 18322 12356 18328 12368
rect 17972 12328 18328 12356
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 15197 12291 15255 12297
rect 15197 12288 15209 12291
rect 12768 12260 15209 12288
rect 12768 12248 12774 12260
rect 15197 12257 15209 12260
rect 15243 12288 15255 12291
rect 17126 12288 17132 12300
rect 15243 12260 17132 12288
rect 15243 12257 15255 12260
rect 15197 12251 15255 12257
rect 17126 12248 17132 12260
rect 17184 12288 17190 12300
rect 17865 12291 17923 12297
rect 17865 12288 17877 12291
rect 17184 12260 17877 12288
rect 17184 12248 17190 12260
rect 17865 12257 17877 12260
rect 17911 12257 17923 12291
rect 17865 12251 17923 12257
rect 17972 12232 18000 12328
rect 18322 12316 18328 12328
rect 18380 12316 18386 12368
rect 24578 12356 24584 12368
rect 23492 12328 24584 12356
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 21450 12288 21456 12300
rect 19392 12260 21456 12288
rect 19392 12248 19398 12260
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12220 14519 12223
rect 14918 12220 14924 12232
rect 14507 12192 14924 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 14918 12180 14924 12192
rect 14976 12180 14982 12232
rect 15562 12180 15568 12232
rect 15620 12180 15626 12232
rect 17954 12220 17960 12232
rect 16592 12192 17960 12220
rect 16592 12138 16620 12192
rect 17954 12180 17960 12192
rect 18012 12180 18018 12232
rect 18046 12180 18052 12232
rect 18104 12220 18110 12232
rect 18141 12223 18199 12229
rect 18141 12220 18153 12223
rect 18104 12192 18153 12220
rect 18104 12180 18110 12192
rect 18141 12189 18153 12192
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12220 18383 12223
rect 19150 12220 19156 12232
rect 18371 12192 19156 12220
rect 18371 12189 18383 12192
rect 18325 12183 18383 12189
rect 19150 12180 19156 12192
rect 19208 12180 19214 12232
rect 19426 12180 19432 12232
rect 19484 12220 19490 12232
rect 19705 12223 19763 12229
rect 19705 12220 19717 12223
rect 19484 12192 19717 12220
rect 19484 12180 19490 12192
rect 19705 12189 19717 12192
rect 19751 12189 19763 12223
rect 19705 12183 19763 12189
rect 19886 12180 19892 12232
rect 19944 12180 19950 12232
rect 21192 12229 21220 12260
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 23492 12229 23520 12328
rect 24578 12316 24584 12328
rect 24636 12316 24642 12368
rect 23584 12260 24624 12288
rect 21177 12223 21235 12229
rect 21177 12189 21189 12223
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 23477 12223 23535 12229
rect 23477 12189 23489 12223
rect 23523 12189 23535 12223
rect 23477 12183 23535 12189
rect 17129 12155 17187 12161
rect 17129 12121 17141 12155
rect 17175 12152 17187 12155
rect 17494 12152 17500 12164
rect 17175 12124 17500 12152
rect 17175 12121 17187 12124
rect 17129 12115 17187 12121
rect 17494 12112 17500 12124
rect 17552 12152 17558 12164
rect 18417 12155 18475 12161
rect 18417 12152 18429 12155
rect 17552 12124 18429 12152
rect 17552 12112 17558 12124
rect 18417 12121 18429 12124
rect 18463 12121 18475 12155
rect 18417 12115 18475 12121
rect 17402 12044 17408 12096
rect 17460 12084 17466 12096
rect 18233 12087 18291 12093
rect 18233 12084 18245 12087
rect 17460 12056 18245 12084
rect 17460 12044 17466 12056
rect 18233 12053 18245 12056
rect 18279 12053 18291 12087
rect 18233 12047 18291 12053
rect 20530 12044 20536 12096
rect 20588 12084 20594 12096
rect 21085 12087 21143 12093
rect 21085 12084 21097 12087
rect 20588 12056 21097 12084
rect 20588 12044 20594 12056
rect 21085 12053 21097 12056
rect 21131 12053 21143 12087
rect 21085 12047 21143 12053
rect 23290 12044 23296 12096
rect 23348 12044 23354 12096
rect 23382 12044 23388 12096
rect 23440 12084 23446 12096
rect 23584 12084 23612 12260
rect 23753 12223 23811 12229
rect 23753 12189 23765 12223
rect 23799 12220 23811 12223
rect 24026 12220 24032 12232
rect 23799 12192 24032 12220
rect 23799 12189 23811 12192
rect 23753 12183 23811 12189
rect 24026 12180 24032 12192
rect 24084 12180 24090 12232
rect 24118 12180 24124 12232
rect 24176 12180 24182 12232
rect 24302 12180 24308 12232
rect 24360 12220 24366 12232
rect 24596 12229 24624 12260
rect 25038 12248 25044 12300
rect 25096 12248 25102 12300
rect 25222 12248 25228 12300
rect 25280 12288 25286 12300
rect 25961 12291 26019 12297
rect 25961 12288 25973 12291
rect 25280 12260 25973 12288
rect 25280 12248 25286 12260
rect 25961 12257 25973 12260
rect 26007 12257 26019 12291
rect 25961 12251 26019 12257
rect 24397 12223 24455 12229
rect 24397 12220 24409 12223
rect 24360 12192 24409 12220
rect 24360 12180 24366 12192
rect 24397 12189 24409 12192
rect 24443 12189 24455 12223
rect 24397 12183 24455 12189
rect 24581 12223 24639 12229
rect 24581 12189 24593 12223
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 25774 12180 25780 12232
rect 25832 12220 25838 12232
rect 25869 12223 25927 12229
rect 25869 12220 25881 12223
rect 25832 12192 25881 12220
rect 25832 12180 25838 12192
rect 25869 12189 25881 12192
rect 25915 12220 25927 12223
rect 26068 12220 26096 12396
rect 28534 12384 28540 12396
rect 28592 12384 28598 12436
rect 32858 12384 32864 12436
rect 32916 12384 32922 12436
rect 34514 12424 34520 12436
rect 32968 12396 34520 12424
rect 26142 12316 26148 12368
rect 26200 12356 26206 12368
rect 26200 12328 27384 12356
rect 26200 12316 26206 12328
rect 26694 12248 26700 12300
rect 26752 12288 26758 12300
rect 27356 12297 27384 12328
rect 27706 12316 27712 12368
rect 27764 12316 27770 12368
rect 32766 12316 32772 12368
rect 32824 12356 32830 12368
rect 32968 12356 32996 12396
rect 34514 12384 34520 12396
rect 34572 12384 34578 12436
rect 35434 12384 35440 12436
rect 35492 12424 35498 12436
rect 35621 12427 35679 12433
rect 35621 12424 35633 12427
rect 35492 12396 35633 12424
rect 35492 12384 35498 12396
rect 35621 12393 35633 12396
rect 35667 12393 35679 12427
rect 35621 12387 35679 12393
rect 35986 12384 35992 12436
rect 36044 12424 36050 12436
rect 36044 12396 37872 12424
rect 36044 12384 36050 12396
rect 32824 12328 32996 12356
rect 32824 12316 32830 12328
rect 27249 12291 27307 12297
rect 27249 12288 27261 12291
rect 26752 12260 27261 12288
rect 26752 12248 26758 12260
rect 27249 12257 27261 12260
rect 27295 12257 27307 12291
rect 27249 12251 27307 12257
rect 27341 12291 27399 12297
rect 27341 12257 27353 12291
rect 27387 12257 27399 12291
rect 27341 12251 27399 12257
rect 27525 12291 27583 12297
rect 27525 12257 27537 12291
rect 27571 12288 27583 12291
rect 27724 12288 27752 12316
rect 27571 12260 28488 12288
rect 27571 12257 27583 12260
rect 27525 12251 27583 12257
rect 25915 12192 26096 12220
rect 25915 12189 25927 12192
rect 25869 12183 25927 12189
rect 26142 12180 26148 12232
rect 26200 12180 26206 12232
rect 26234 12180 26240 12232
rect 26292 12180 26298 12232
rect 27433 12223 27491 12229
rect 27433 12189 27445 12223
rect 27479 12220 27491 12223
rect 27706 12220 27712 12232
rect 27479 12192 27712 12220
rect 27479 12189 27491 12192
rect 27433 12183 27491 12189
rect 27706 12180 27712 12192
rect 27764 12180 27770 12232
rect 27890 12180 27896 12232
rect 27948 12180 27954 12232
rect 27982 12180 27988 12232
rect 28040 12180 28046 12232
rect 28077 12223 28135 12229
rect 28077 12189 28089 12223
rect 28123 12220 28135 12223
rect 28258 12220 28264 12232
rect 28123 12192 28264 12220
rect 28123 12189 28135 12192
rect 28077 12183 28135 12189
rect 28258 12180 28264 12192
rect 28316 12180 28322 12232
rect 28460 12229 28488 12260
rect 28626 12248 28632 12300
rect 28684 12288 28690 12300
rect 31389 12291 31447 12297
rect 28684 12260 28856 12288
rect 28684 12248 28690 12260
rect 28828 12229 28856 12260
rect 31389 12257 31401 12291
rect 31435 12288 31447 12291
rect 31478 12288 31484 12300
rect 31435 12260 31484 12288
rect 31435 12257 31447 12260
rect 31389 12251 31447 12257
rect 31478 12248 31484 12260
rect 31536 12248 31542 12300
rect 28445 12223 28503 12229
rect 28445 12189 28457 12223
rect 28491 12189 28503 12223
rect 28445 12183 28503 12189
rect 28537 12223 28595 12229
rect 28537 12189 28549 12223
rect 28583 12189 28595 12223
rect 28537 12183 28595 12189
rect 28721 12223 28779 12229
rect 28721 12189 28733 12223
rect 28767 12189 28779 12223
rect 28721 12183 28779 12189
rect 28813 12223 28871 12229
rect 28813 12189 28825 12223
rect 28859 12189 28871 12223
rect 28813 12183 28871 12189
rect 24210 12112 24216 12164
rect 24268 12152 24274 12164
rect 25317 12155 25375 12161
rect 25317 12152 25329 12155
rect 24268 12124 25329 12152
rect 24268 12112 24274 12124
rect 25317 12121 25329 12124
rect 25363 12121 25375 12155
rect 25317 12115 25375 12121
rect 26421 12155 26479 12161
rect 26421 12121 26433 12155
rect 26467 12152 26479 12155
rect 28166 12152 28172 12164
rect 26467 12124 28172 12152
rect 26467 12121 26479 12124
rect 26421 12115 26479 12121
rect 28166 12112 28172 12124
rect 28224 12112 28230 12164
rect 28353 12155 28411 12161
rect 28353 12121 28365 12155
rect 28399 12152 28411 12155
rect 28552 12152 28580 12183
rect 28399 12124 28580 12152
rect 28736 12152 28764 12183
rect 29454 12180 29460 12232
rect 29512 12220 29518 12232
rect 31113 12223 31171 12229
rect 31113 12220 31125 12223
rect 29512 12192 31125 12220
rect 29512 12180 29518 12192
rect 31113 12189 31125 12192
rect 31159 12189 31171 12223
rect 32968 12220 32996 12328
rect 33226 12316 33232 12368
rect 33284 12356 33290 12368
rect 34238 12356 34244 12368
rect 33284 12328 34244 12356
rect 33284 12316 33290 12328
rect 34238 12316 34244 12328
rect 34296 12356 34302 12368
rect 35710 12356 35716 12368
rect 34296 12328 35716 12356
rect 34296 12316 34302 12328
rect 33594 12288 33600 12300
rect 33336 12260 33600 12288
rect 33336 12229 33364 12260
rect 33594 12248 33600 12260
rect 33652 12248 33658 12300
rect 33045 12223 33103 12229
rect 33045 12220 33057 12223
rect 32968 12192 33057 12220
rect 31113 12183 31171 12189
rect 33045 12189 33057 12192
rect 33091 12189 33103 12223
rect 33045 12183 33103 12189
rect 33138 12223 33196 12229
rect 33138 12189 33150 12223
rect 33184 12189 33196 12223
rect 33138 12183 33196 12189
rect 33321 12223 33379 12229
rect 33321 12189 33333 12223
rect 33367 12189 33379 12223
rect 33321 12183 33379 12189
rect 28736 12124 29224 12152
rect 28399 12121 28411 12124
rect 28353 12115 28411 12121
rect 23937 12087 23995 12093
rect 23937 12084 23949 12087
rect 23440 12056 23949 12084
rect 23440 12044 23446 12056
rect 23937 12053 23949 12056
rect 23983 12053 23995 12087
rect 23937 12047 23995 12053
rect 24026 12044 24032 12096
rect 24084 12084 24090 12096
rect 25225 12087 25283 12093
rect 25225 12084 25237 12087
rect 24084 12056 25237 12084
rect 24084 12044 24090 12056
rect 25225 12053 25237 12056
rect 25271 12084 25283 12087
rect 25866 12084 25872 12096
rect 25271 12056 25872 12084
rect 25271 12053 25283 12056
rect 25225 12047 25283 12053
rect 25866 12044 25872 12056
rect 25924 12044 25930 12096
rect 26602 12044 26608 12096
rect 26660 12084 26666 12096
rect 27062 12084 27068 12096
rect 26660 12056 27068 12084
rect 26660 12044 26666 12056
rect 27062 12044 27068 12056
rect 27120 12044 27126 12096
rect 27890 12044 27896 12096
rect 27948 12084 27954 12096
rect 29196 12093 29224 12124
rect 31846 12112 31852 12164
rect 31904 12112 31910 12164
rect 32858 12112 32864 12164
rect 32916 12152 32922 12164
rect 33152 12152 33180 12183
rect 33410 12180 33416 12232
rect 33468 12180 33474 12232
rect 33502 12180 33508 12232
rect 33560 12229 33566 12232
rect 33560 12220 33568 12229
rect 33965 12223 34023 12229
rect 33965 12220 33977 12223
rect 33560 12192 33605 12220
rect 33704 12192 33977 12220
rect 33560 12183 33568 12192
rect 33560 12180 33566 12183
rect 32916 12124 33180 12152
rect 32916 12112 32922 12124
rect 28997 12087 29055 12093
rect 28997 12084 29009 12087
rect 27948 12056 29009 12084
rect 27948 12044 27954 12056
rect 28997 12053 29009 12056
rect 29043 12053 29055 12087
rect 28997 12047 29055 12053
rect 29181 12087 29239 12093
rect 29181 12053 29193 12087
rect 29227 12084 29239 12087
rect 29822 12084 29828 12096
rect 29227 12056 29828 12084
rect 29227 12053 29239 12056
rect 29181 12047 29239 12053
rect 29822 12044 29828 12056
rect 29880 12044 29886 12096
rect 33704 12093 33732 12192
rect 33965 12189 33977 12192
rect 34011 12189 34023 12223
rect 33965 12183 34023 12189
rect 34146 12180 34152 12232
rect 34204 12180 34210 12232
rect 34238 12180 34244 12232
rect 34296 12180 34302 12232
rect 35084 12229 35112 12328
rect 35710 12316 35716 12328
rect 35768 12316 35774 12368
rect 36630 12316 36636 12368
rect 36688 12356 36694 12368
rect 37366 12356 37372 12368
rect 36688 12328 37372 12356
rect 36688 12316 36694 12328
rect 37366 12316 37372 12328
rect 37424 12356 37430 12368
rect 37461 12359 37519 12365
rect 37461 12356 37473 12359
rect 37424 12328 37473 12356
rect 37424 12316 37430 12328
rect 37461 12325 37473 12328
rect 37507 12325 37519 12359
rect 37461 12319 37519 12325
rect 35342 12288 35348 12300
rect 35268 12260 35348 12288
rect 35268 12229 35296 12260
rect 35342 12248 35348 12260
rect 35400 12248 35406 12300
rect 37550 12288 37556 12300
rect 37200 12260 37556 12288
rect 34977 12223 35035 12229
rect 34977 12189 34989 12223
rect 35023 12189 35035 12223
rect 34977 12183 35035 12189
rect 35070 12223 35128 12229
rect 35070 12189 35082 12223
rect 35116 12189 35128 12223
rect 35070 12183 35128 12189
rect 35253 12223 35311 12229
rect 35253 12189 35265 12223
rect 35299 12189 35311 12223
rect 35253 12183 35311 12189
rect 35483 12223 35541 12229
rect 35483 12189 35495 12223
rect 35529 12220 35541 12223
rect 37200 12220 37228 12260
rect 37550 12248 37556 12260
rect 37608 12248 37614 12300
rect 37844 12232 37872 12396
rect 42150 12384 42156 12436
rect 42208 12384 42214 12436
rect 42886 12384 42892 12436
rect 42944 12384 42950 12436
rect 44453 12427 44511 12433
rect 44453 12393 44465 12427
rect 44499 12424 44511 12427
rect 44542 12424 44548 12436
rect 44499 12396 44548 12424
rect 44499 12393 44511 12396
rect 44453 12387 44511 12393
rect 44542 12384 44548 12396
rect 44600 12384 44606 12436
rect 45281 12427 45339 12433
rect 45281 12393 45293 12427
rect 45327 12424 45339 12427
rect 45370 12424 45376 12436
rect 45327 12396 45376 12424
rect 45327 12393 45339 12396
rect 45281 12387 45339 12393
rect 45370 12384 45376 12396
rect 45428 12384 45434 12436
rect 45649 12427 45707 12433
rect 45649 12393 45661 12427
rect 45695 12424 45707 12427
rect 46934 12424 46940 12436
rect 45695 12396 46940 12424
rect 45695 12393 45707 12396
rect 45649 12387 45707 12393
rect 42794 12356 42800 12368
rect 42725 12328 42800 12356
rect 40678 12248 40684 12300
rect 40736 12248 40742 12300
rect 42150 12248 42156 12300
rect 42208 12288 42214 12300
rect 42725 12288 42753 12328
rect 42794 12316 42800 12328
rect 42852 12356 42858 12368
rect 42852 12328 43898 12356
rect 42852 12316 42858 12328
rect 42208 12260 42380 12288
rect 42208 12248 42214 12260
rect 35529 12192 37228 12220
rect 35529 12189 35541 12192
rect 35483 12183 35541 12189
rect 33781 12155 33839 12161
rect 33781 12121 33793 12155
rect 33827 12152 33839 12155
rect 33827 12124 33962 12152
rect 33827 12121 33839 12124
rect 33781 12115 33839 12121
rect 33934 12096 33962 12124
rect 34514 12112 34520 12164
rect 34572 12152 34578 12164
rect 34992 12152 35020 12183
rect 37274 12180 37280 12232
rect 37332 12180 37338 12232
rect 37737 12223 37795 12229
rect 37737 12189 37749 12223
rect 37783 12189 37795 12223
rect 37737 12183 37795 12189
rect 35345 12155 35403 12161
rect 34572 12124 35112 12152
rect 34572 12112 34578 12124
rect 33689 12087 33747 12093
rect 33689 12053 33701 12087
rect 33735 12053 33747 12087
rect 33934 12056 33968 12096
rect 33689 12047 33747 12053
rect 33962 12044 33968 12056
rect 34020 12044 34026 12096
rect 35084 12084 35112 12124
rect 35345 12121 35357 12155
rect 35391 12152 35403 12155
rect 35986 12152 35992 12164
rect 35391 12124 35992 12152
rect 35391 12121 35403 12124
rect 35345 12115 35403 12121
rect 35986 12112 35992 12124
rect 36044 12112 36050 12164
rect 37752 12084 37780 12183
rect 37826 12180 37832 12232
rect 37884 12180 37890 12232
rect 38102 12180 38108 12232
rect 38160 12180 38166 12232
rect 38202 12223 38260 12229
rect 38202 12189 38214 12223
rect 38248 12220 38260 12223
rect 38470 12220 38476 12232
rect 38248 12192 38476 12220
rect 38248 12189 38260 12192
rect 38202 12183 38260 12189
rect 38470 12180 38476 12192
rect 38528 12180 38534 12232
rect 40218 12180 40224 12232
rect 40276 12220 40282 12232
rect 42352 12229 42380 12260
rect 42628 12260 42753 12288
rect 43870 12288 43898 12328
rect 44174 12316 44180 12368
rect 44232 12356 44238 12368
rect 45664 12356 45692 12387
rect 46934 12384 46940 12396
rect 46992 12384 46998 12436
rect 50338 12384 50344 12436
rect 50396 12424 50402 12436
rect 50396 12396 55996 12424
rect 50396 12384 50402 12396
rect 44232 12328 45692 12356
rect 44232 12316 44238 12328
rect 46842 12288 46848 12300
rect 43870 12260 46848 12288
rect 42628 12229 42656 12260
rect 46842 12248 46848 12260
rect 46900 12288 46906 12300
rect 46937 12291 46995 12297
rect 46937 12288 46949 12291
rect 46900 12260 46949 12288
rect 46900 12248 46906 12260
rect 46937 12257 46949 12260
rect 46983 12257 46995 12291
rect 50341 12291 50399 12297
rect 50341 12288 50353 12291
rect 46937 12251 46995 12257
rect 47136 12260 50353 12288
rect 47136 12232 47164 12260
rect 50341 12257 50353 12260
rect 50387 12288 50399 12291
rect 51810 12288 51816 12300
rect 50387 12260 51816 12288
rect 50387 12257 50399 12260
rect 50341 12251 50399 12257
rect 51810 12248 51816 12260
rect 51868 12248 51874 12300
rect 52457 12291 52515 12297
rect 52457 12257 52469 12291
rect 52503 12288 52515 12291
rect 54018 12288 54024 12300
rect 52503 12260 54024 12288
rect 52503 12257 52515 12260
rect 52457 12251 52515 12257
rect 54018 12248 54024 12260
rect 54076 12288 54082 12300
rect 54202 12288 54208 12300
rect 54076 12260 54208 12288
rect 54076 12248 54082 12260
rect 54202 12248 54208 12260
rect 54260 12248 54266 12300
rect 40405 12223 40463 12229
rect 40405 12220 40417 12223
rect 40276 12192 40417 12220
rect 40276 12180 40282 12192
rect 40405 12189 40417 12192
rect 40451 12189 40463 12223
rect 40405 12183 40463 12189
rect 42245 12223 42303 12229
rect 42245 12189 42257 12223
rect 42291 12189 42303 12223
rect 42245 12183 42303 12189
rect 42338 12223 42396 12229
rect 42338 12189 42350 12223
rect 42384 12189 42396 12223
rect 42338 12183 42396 12189
rect 42613 12223 42671 12229
rect 42613 12189 42625 12223
rect 42659 12189 42671 12223
rect 42613 12183 42671 12189
rect 42710 12223 42768 12229
rect 42710 12189 42722 12223
rect 42756 12189 42768 12223
rect 43622 12220 43628 12232
rect 42710 12183 42768 12189
rect 42904 12192 43628 12220
rect 38013 12155 38071 12161
rect 38013 12121 38025 12155
rect 38059 12121 38071 12155
rect 38013 12115 38071 12121
rect 35084 12056 37780 12084
rect 38028 12084 38056 12115
rect 39114 12112 39120 12164
rect 39172 12152 39178 12164
rect 39172 12124 41170 12152
rect 39172 12112 39178 12124
rect 38102 12084 38108 12096
rect 38028 12056 38108 12084
rect 38102 12044 38108 12056
rect 38160 12044 38166 12096
rect 38378 12044 38384 12096
rect 38436 12044 38442 12096
rect 42260 12084 42288 12183
rect 42518 12112 42524 12164
rect 42576 12112 42582 12164
rect 42725 12152 42753 12183
rect 42904 12152 42932 12192
rect 43622 12180 43628 12192
rect 43680 12180 43686 12232
rect 45465 12223 45523 12229
rect 45465 12189 45477 12223
rect 45511 12220 45523 12223
rect 45554 12220 45560 12232
rect 45511 12192 45560 12220
rect 45511 12189 45523 12192
rect 45465 12183 45523 12189
rect 45554 12180 45560 12192
rect 45612 12180 45618 12232
rect 45741 12223 45799 12229
rect 45741 12189 45753 12223
rect 45787 12220 45799 12223
rect 46385 12223 46443 12229
rect 46385 12220 46397 12223
rect 45787 12192 46397 12220
rect 45787 12189 45799 12192
rect 45741 12183 45799 12189
rect 46385 12189 46397 12192
rect 46431 12189 46443 12223
rect 46385 12183 46443 12189
rect 47118 12180 47124 12232
rect 47176 12180 47182 12232
rect 55398 12180 55404 12232
rect 55456 12220 55462 12232
rect 55968 12229 55996 12396
rect 55585 12223 55643 12229
rect 55585 12220 55597 12223
rect 55456 12192 55597 12220
rect 55456 12180 55462 12192
rect 55585 12189 55597 12192
rect 55631 12189 55643 12223
rect 55585 12183 55643 12189
rect 55953 12223 56011 12229
rect 55953 12189 55965 12223
rect 55999 12220 56011 12223
rect 56137 12223 56195 12229
rect 56137 12220 56149 12223
rect 55999 12192 56149 12220
rect 55999 12189 56011 12192
rect 55953 12183 56011 12189
rect 56137 12189 56149 12192
rect 56183 12189 56195 12223
rect 56137 12183 56195 12189
rect 42725 12124 42932 12152
rect 47397 12155 47455 12161
rect 47397 12121 47409 12155
rect 47443 12152 47455 12155
rect 47670 12152 47676 12164
rect 47443 12124 47676 12152
rect 47443 12121 47455 12124
rect 47397 12115 47455 12121
rect 47670 12112 47676 12124
rect 47728 12112 47734 12164
rect 49234 12152 49240 12164
rect 48622 12124 49240 12152
rect 49234 12112 49240 12124
rect 49292 12152 49298 12164
rect 50338 12152 50344 12164
rect 49292 12124 50344 12152
rect 49292 12112 49298 12124
rect 50338 12112 50344 12124
rect 50396 12112 50402 12164
rect 50617 12155 50675 12161
rect 50617 12121 50629 12155
rect 50663 12152 50675 12155
rect 50706 12152 50712 12164
rect 50663 12124 50712 12152
rect 50663 12121 50675 12124
rect 50617 12115 50675 12121
rect 50706 12112 50712 12124
rect 50764 12112 50770 12164
rect 51842 12124 52592 12152
rect 44266 12084 44272 12096
rect 42260 12056 44272 12084
rect 44266 12044 44272 12056
rect 44324 12044 44330 12096
rect 48314 12044 48320 12096
rect 48372 12084 48378 12096
rect 48869 12087 48927 12093
rect 48869 12084 48881 12087
rect 48372 12056 48881 12084
rect 48372 12044 48378 12056
rect 48869 12053 48881 12056
rect 48915 12053 48927 12087
rect 48869 12047 48927 12053
rect 51534 12044 51540 12096
rect 51592 12084 51598 12096
rect 51920 12084 51948 12124
rect 51592 12056 51948 12084
rect 52089 12087 52147 12093
rect 51592 12044 51598 12056
rect 52089 12053 52101 12087
rect 52135 12084 52147 12087
rect 52270 12084 52276 12096
rect 52135 12056 52276 12084
rect 52135 12053 52147 12056
rect 52089 12047 52147 12053
rect 52270 12044 52276 12056
rect 52328 12044 52334 12096
rect 52564 12084 52592 12124
rect 52638 12112 52644 12164
rect 52696 12152 52702 12164
rect 52733 12155 52791 12161
rect 52733 12152 52745 12155
rect 52696 12124 52745 12152
rect 52696 12112 52702 12124
rect 52733 12121 52745 12124
rect 52779 12121 52791 12155
rect 55600 12152 55628 12183
rect 55858 12152 55864 12164
rect 52733 12115 52791 12121
rect 53116 12124 53222 12152
rect 55600 12124 55864 12152
rect 53116 12084 53144 12124
rect 55858 12112 55864 12124
rect 55916 12112 55922 12164
rect 52564 12056 53144 12084
rect 54110 12044 54116 12096
rect 54168 12084 54174 12096
rect 54205 12087 54263 12093
rect 54205 12084 54217 12087
rect 54168 12056 54217 12084
rect 54168 12044 54174 12056
rect 54205 12053 54217 12056
rect 54251 12053 54263 12087
rect 54205 12047 54263 12053
rect 54938 12044 54944 12096
rect 54996 12084 55002 12096
rect 56229 12087 56287 12093
rect 56229 12084 56241 12087
rect 54996 12056 56241 12084
rect 54996 12044 55002 12056
rect 56229 12053 56241 12056
rect 56275 12053 56287 12087
rect 56229 12047 56287 12053
rect 1104 11994 78844 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 66314 11994
rect 66366 11942 66378 11994
rect 66430 11942 66442 11994
rect 66494 11942 66506 11994
rect 66558 11942 66570 11994
rect 66622 11942 78844 11994
rect 1104 11920 78844 11942
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11880 14519 11883
rect 14826 11880 14832 11892
rect 14507 11852 14832 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 15562 11840 15568 11892
rect 15620 11880 15626 11892
rect 17037 11883 17095 11889
rect 17037 11880 17049 11883
rect 15620 11852 17049 11880
rect 15620 11840 15626 11852
rect 17037 11849 17049 11852
rect 17083 11849 17095 11883
rect 18874 11880 18880 11892
rect 17037 11843 17095 11849
rect 17328 11852 18880 11880
rect 12986 11772 12992 11824
rect 13044 11772 13050 11824
rect 13998 11772 14004 11824
rect 14056 11772 14062 11824
rect 17328 11821 17356 11852
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 22925 11883 22983 11889
rect 22925 11849 22937 11883
rect 22971 11880 22983 11883
rect 22971 11852 23980 11880
rect 22971 11849 22983 11852
rect 22925 11843 22983 11849
rect 17313 11815 17371 11821
rect 17313 11781 17325 11815
rect 17359 11781 17371 11815
rect 17313 11775 17371 11781
rect 17402 11772 17408 11824
rect 17460 11772 17466 11824
rect 17543 11815 17601 11821
rect 17543 11781 17555 11815
rect 17589 11812 17601 11815
rect 18138 11812 18144 11824
rect 17589 11784 18144 11812
rect 17589 11781 17601 11784
rect 17543 11775 17601 11781
rect 18138 11772 18144 11784
rect 18196 11772 18202 11824
rect 22186 11772 22192 11824
rect 22244 11812 22250 11824
rect 23382 11812 23388 11824
rect 22244 11784 23388 11812
rect 22244 11772 22250 11784
rect 12710 11704 12716 11756
rect 12768 11704 12774 11756
rect 16942 11704 16948 11756
rect 17000 11744 17006 11756
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 17000 11716 17233 11744
rect 17000 11704 17006 11716
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 17678 11704 17684 11756
rect 17736 11704 17742 11756
rect 21174 11704 21180 11756
rect 21232 11744 21238 11756
rect 22646 11744 22652 11756
rect 21232 11716 22652 11744
rect 21232 11704 21238 11716
rect 22646 11704 22652 11716
rect 22704 11704 22710 11756
rect 22833 11747 22891 11753
rect 22833 11713 22845 11747
rect 22879 11744 22891 11747
rect 22922 11744 22928 11756
rect 22879 11716 22928 11744
rect 22879 11713 22891 11716
rect 22833 11707 22891 11713
rect 22922 11704 22928 11716
rect 22980 11704 22986 11756
rect 23216 11753 23244 11784
rect 23382 11772 23388 11784
rect 23440 11772 23446 11824
rect 23952 11812 23980 11852
rect 24118 11840 24124 11892
rect 24176 11880 24182 11892
rect 34333 11883 34391 11889
rect 34333 11880 34345 11883
rect 24176 11852 28304 11880
rect 24176 11840 24182 11852
rect 24946 11812 24952 11824
rect 23584 11784 23796 11812
rect 23952 11784 24952 11812
rect 23201 11747 23259 11753
rect 23201 11713 23213 11747
rect 23247 11713 23259 11747
rect 23201 11707 23259 11713
rect 23290 11704 23296 11756
rect 23348 11704 23354 11756
rect 20530 11636 20536 11688
rect 20588 11676 20594 11688
rect 22741 11679 22799 11685
rect 20588 11648 22094 11676
rect 20588 11636 20594 11648
rect 22066 11608 22094 11648
rect 22741 11645 22753 11679
rect 22787 11676 22799 11679
rect 23584 11676 23612 11784
rect 23658 11704 23664 11756
rect 23716 11704 23722 11756
rect 22787 11648 23612 11676
rect 22787 11645 22799 11648
rect 22741 11639 22799 11645
rect 23308 11620 23336 11648
rect 22922 11608 22928 11620
rect 22066 11580 22928 11608
rect 22922 11568 22928 11580
rect 22980 11568 22986 11620
rect 23290 11568 23296 11620
rect 23348 11568 23354 11620
rect 23676 11608 23704 11704
rect 23768 11676 23796 11784
rect 24946 11772 24952 11784
rect 25004 11772 25010 11824
rect 25866 11772 25872 11824
rect 25924 11812 25930 11824
rect 26053 11815 26111 11821
rect 26053 11812 26065 11815
rect 25924 11784 26065 11812
rect 25924 11772 25930 11784
rect 26053 11781 26065 11784
rect 26099 11781 26111 11815
rect 26053 11775 26111 11781
rect 26234 11772 26240 11824
rect 26292 11812 26298 11824
rect 27982 11812 27988 11824
rect 26292 11784 27568 11812
rect 26292 11772 26298 11784
rect 27540 11756 27568 11784
rect 27632 11784 27988 11812
rect 27632 11756 27660 11784
rect 27982 11772 27988 11784
rect 28040 11772 28046 11824
rect 23934 11704 23940 11756
rect 23992 11704 23998 11756
rect 24302 11744 24308 11756
rect 24044 11716 24308 11744
rect 24044 11676 24072 11716
rect 24302 11704 24308 11716
rect 24360 11704 24366 11756
rect 24486 11704 24492 11756
rect 24544 11704 24550 11756
rect 25222 11704 25228 11756
rect 25280 11704 25286 11756
rect 25314 11704 25320 11756
rect 25372 11744 25378 11756
rect 25409 11747 25467 11753
rect 25409 11744 25421 11747
rect 25372 11716 25421 11744
rect 25372 11704 25378 11716
rect 25409 11713 25421 11716
rect 25455 11713 25467 11747
rect 25409 11707 25467 11713
rect 25593 11747 25651 11753
rect 25593 11713 25605 11747
rect 25639 11744 25651 11747
rect 27433 11747 27491 11753
rect 27433 11744 27445 11747
rect 25639 11716 26096 11744
rect 25639 11713 25651 11716
rect 25593 11707 25651 11713
rect 23768 11648 24072 11676
rect 24210 11636 24216 11688
rect 24268 11636 24274 11688
rect 24397 11679 24455 11685
rect 24397 11645 24409 11679
rect 24443 11676 24455 11679
rect 24578 11676 24584 11688
rect 24443 11648 24584 11676
rect 24443 11645 24455 11648
rect 24397 11639 24455 11645
rect 24578 11636 24584 11648
rect 24636 11636 24642 11688
rect 25424 11676 25452 11707
rect 26068 11688 26096 11716
rect 27356 11716 27445 11744
rect 25866 11676 25872 11688
rect 25424 11648 25872 11676
rect 25866 11636 25872 11648
rect 25924 11636 25930 11688
rect 25961 11679 26019 11685
rect 25961 11645 25973 11679
rect 26007 11645 26019 11679
rect 25961 11639 26019 11645
rect 25976 11608 26004 11639
rect 26050 11636 26056 11688
rect 26108 11636 26114 11688
rect 26510 11636 26516 11688
rect 26568 11676 26574 11688
rect 27356 11676 27384 11716
rect 27433 11713 27445 11716
rect 27479 11713 27491 11747
rect 27433 11707 27491 11713
rect 27522 11704 27528 11756
rect 27580 11704 27586 11756
rect 27614 11704 27620 11756
rect 27672 11704 27678 11756
rect 27706 11704 27712 11756
rect 27764 11744 27770 11756
rect 28169 11747 28227 11753
rect 28169 11744 28181 11747
rect 27764 11716 28181 11744
rect 27764 11704 27770 11716
rect 28169 11713 28181 11716
rect 28215 11713 28227 11747
rect 28169 11707 28227 11713
rect 26568 11648 27384 11676
rect 26568 11636 26574 11648
rect 27356 11608 27384 11648
rect 27893 11679 27951 11685
rect 27893 11645 27905 11679
rect 27939 11676 27951 11679
rect 28276 11676 28304 11852
rect 33888 11852 34345 11880
rect 31846 11812 31852 11824
rect 30958 11784 31852 11812
rect 31846 11772 31852 11784
rect 31904 11812 31910 11824
rect 32122 11812 32128 11824
rect 31904 11784 32128 11812
rect 31904 11772 31910 11784
rect 32122 11772 32128 11784
rect 32180 11772 32186 11824
rect 33888 11812 33916 11852
rect 34333 11849 34345 11852
rect 34379 11880 34391 11883
rect 34790 11880 34796 11892
rect 34379 11852 34796 11880
rect 34379 11849 34391 11852
rect 34333 11843 34391 11849
rect 34790 11840 34796 11852
rect 34848 11840 34854 11892
rect 36538 11840 36544 11892
rect 36596 11880 36602 11892
rect 37090 11880 37096 11892
rect 36596 11852 37096 11880
rect 36596 11840 36602 11852
rect 37090 11840 37096 11852
rect 37148 11840 37154 11892
rect 37458 11840 37464 11892
rect 37516 11880 37522 11892
rect 40405 11883 40463 11889
rect 37516 11852 40361 11880
rect 37516 11840 37522 11852
rect 33534 11784 33916 11812
rect 33962 11772 33968 11824
rect 34020 11772 34026 11824
rect 36280 11784 37136 11812
rect 29454 11704 29460 11756
rect 29512 11704 29518 11756
rect 34241 11747 34299 11753
rect 34241 11713 34253 11747
rect 34287 11744 34299 11747
rect 34514 11744 34520 11756
rect 34287 11716 34520 11744
rect 34287 11713 34299 11716
rect 34241 11707 34299 11713
rect 34514 11704 34520 11716
rect 34572 11704 34578 11756
rect 27939 11648 28304 11676
rect 27939 11645 27951 11648
rect 27893 11639 27951 11645
rect 29730 11636 29736 11688
rect 29788 11636 29794 11688
rect 31386 11636 31392 11688
rect 31444 11676 31450 11688
rect 36280 11685 36308 11784
rect 36630 11753 36636 11756
rect 36628 11707 36636 11753
rect 36630 11704 36636 11707
rect 36688 11704 36694 11756
rect 36725 11747 36783 11753
rect 36725 11713 36737 11747
rect 36771 11713 36783 11747
rect 36725 11707 36783 11713
rect 36817 11747 36875 11753
rect 36817 11713 36829 11747
rect 36863 11713 36875 11747
rect 36817 11707 36875 11713
rect 36265 11679 36323 11685
rect 36265 11676 36277 11679
rect 31444 11648 36277 11676
rect 31444 11636 31450 11648
rect 36265 11645 36277 11648
rect 36311 11645 36323 11679
rect 36265 11639 36323 11645
rect 36538 11636 36544 11688
rect 36596 11676 36602 11688
rect 36740 11676 36768 11707
rect 36596 11648 36768 11676
rect 36832 11676 36860 11707
rect 36906 11704 36912 11756
rect 36964 11753 36970 11756
rect 37108 11753 37136 11784
rect 37550 11772 37556 11824
rect 37608 11812 37614 11824
rect 38470 11812 38476 11824
rect 37608 11784 38476 11812
rect 37608 11772 37614 11784
rect 38470 11772 38476 11784
rect 38528 11812 38534 11824
rect 38528 11784 40269 11812
rect 38528 11772 38534 11784
rect 36964 11747 37003 11753
rect 36991 11713 37003 11747
rect 36964 11707 37003 11713
rect 37093 11747 37151 11753
rect 37093 11713 37105 11747
rect 37139 11713 37151 11747
rect 37093 11707 37151 11713
rect 36964 11704 36970 11707
rect 37826 11704 37832 11756
rect 37884 11704 37890 11756
rect 38378 11704 38384 11756
rect 38436 11704 38442 11756
rect 39482 11704 39488 11756
rect 39540 11744 39546 11756
rect 40241 11753 40269 11784
rect 39761 11747 39819 11753
rect 39761 11744 39773 11747
rect 39540 11716 39773 11744
rect 39540 11704 39546 11716
rect 39761 11713 39773 11716
rect 39807 11713 39819 11747
rect 39761 11707 39819 11713
rect 39854 11747 39912 11753
rect 39854 11713 39866 11747
rect 39900 11713 39912 11747
rect 39854 11707 39912 11713
rect 40037 11747 40095 11753
rect 40037 11713 40049 11747
rect 40083 11713 40095 11747
rect 40037 11707 40095 11713
rect 40126 11747 40184 11753
rect 40126 11713 40138 11747
rect 40172 11713 40184 11747
rect 40126 11707 40184 11713
rect 40226 11747 40284 11753
rect 40226 11713 40238 11747
rect 40272 11713 40284 11747
rect 40226 11707 40284 11713
rect 36832 11648 36952 11676
rect 36596 11636 36602 11648
rect 28258 11608 28264 11620
rect 23676 11580 26004 11608
rect 26068 11580 27292 11608
rect 27356 11580 28264 11608
rect 17865 11543 17923 11549
rect 17865 11509 17877 11543
rect 17911 11540 17923 11543
rect 17954 11540 17960 11552
rect 17911 11512 17960 11540
rect 17911 11509 17923 11512
rect 17865 11503 17923 11509
rect 17954 11500 17960 11512
rect 18012 11540 18018 11552
rect 18690 11540 18696 11552
rect 18012 11512 18696 11540
rect 18012 11500 18018 11512
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 23382 11500 23388 11552
rect 23440 11500 23446 11552
rect 23477 11543 23535 11549
rect 23477 11509 23489 11543
rect 23523 11540 23535 11543
rect 23753 11543 23811 11549
rect 23753 11540 23765 11543
rect 23523 11512 23765 11540
rect 23523 11509 23535 11512
rect 23477 11503 23535 11509
rect 23753 11509 23765 11512
rect 23799 11509 23811 11543
rect 23753 11503 23811 11509
rect 24118 11500 24124 11552
rect 24176 11500 24182 11552
rect 25866 11500 25872 11552
rect 25924 11540 25930 11552
rect 26068 11540 26096 11580
rect 27264 11552 27292 11580
rect 28258 11568 28264 11580
rect 28316 11568 28322 11620
rect 25924 11512 26096 11540
rect 25924 11500 25930 11512
rect 26418 11500 26424 11552
rect 26476 11500 26482 11552
rect 27246 11500 27252 11552
rect 27304 11500 27310 11552
rect 31202 11500 31208 11552
rect 31260 11500 31266 11552
rect 31662 11500 31668 11552
rect 31720 11540 31726 11552
rect 32493 11543 32551 11549
rect 32493 11540 32505 11543
rect 31720 11512 32505 11540
rect 31720 11500 31726 11512
rect 32493 11509 32505 11512
rect 32539 11540 32551 11543
rect 33226 11540 33232 11552
rect 32539 11512 33232 11540
rect 32539 11509 32551 11512
rect 32493 11503 32551 11509
rect 33226 11500 33232 11512
rect 33284 11500 33290 11552
rect 33594 11500 33600 11552
rect 33652 11540 33658 11552
rect 34422 11540 34428 11552
rect 33652 11512 34428 11540
rect 33652 11500 33658 11512
rect 34422 11500 34428 11512
rect 34480 11500 34486 11552
rect 36449 11543 36507 11549
rect 36449 11509 36461 11543
rect 36495 11540 36507 11543
rect 36538 11540 36544 11552
rect 36495 11512 36544 11540
rect 36495 11509 36507 11512
rect 36449 11503 36507 11509
rect 36538 11500 36544 11512
rect 36596 11500 36602 11552
rect 36924 11540 36952 11648
rect 37274 11636 37280 11688
rect 37332 11636 37338 11688
rect 38657 11679 38715 11685
rect 38657 11645 38669 11679
rect 38703 11676 38715 11679
rect 39025 11679 39083 11685
rect 39025 11676 39037 11679
rect 38703 11648 39037 11676
rect 38703 11645 38715 11648
rect 38657 11639 38715 11645
rect 39025 11645 39037 11648
rect 39071 11645 39083 11679
rect 39025 11639 39083 11645
rect 39577 11679 39635 11685
rect 39577 11645 39589 11679
rect 39623 11676 39635 11679
rect 39868 11676 39896 11707
rect 39623 11648 39896 11676
rect 39623 11645 39635 11648
rect 39577 11639 39635 11645
rect 37090 11568 37096 11620
rect 37148 11608 37154 11620
rect 39592 11608 39620 11639
rect 39666 11608 39672 11620
rect 37148 11580 39672 11608
rect 37148 11568 37154 11580
rect 39666 11568 39672 11580
rect 39724 11568 39730 11620
rect 38102 11540 38108 11552
rect 36924 11512 38108 11540
rect 38102 11500 38108 11512
rect 38160 11500 38166 11552
rect 38194 11500 38200 11552
rect 38252 11500 38258 11552
rect 38562 11500 38568 11552
rect 38620 11500 38626 11552
rect 40052 11540 40080 11707
rect 40144 11620 40172 11707
rect 40333 11676 40361 11852
rect 40405 11849 40417 11883
rect 40451 11880 40463 11883
rect 40586 11880 40592 11892
rect 40451 11852 40592 11880
rect 40451 11849 40463 11852
rect 40405 11843 40463 11849
rect 40586 11840 40592 11852
rect 40644 11840 40650 11892
rect 47670 11840 47676 11892
rect 47728 11840 47734 11892
rect 47946 11840 47952 11892
rect 48004 11880 48010 11892
rect 48317 11883 48375 11889
rect 48317 11880 48329 11883
rect 48004 11852 48329 11880
rect 48004 11840 48010 11852
rect 48317 11849 48329 11852
rect 48363 11849 48375 11883
rect 48317 11843 48375 11849
rect 49697 11883 49755 11889
rect 49697 11849 49709 11883
rect 49743 11880 49755 11883
rect 49743 11852 49832 11880
rect 49743 11849 49755 11852
rect 49697 11843 49755 11849
rect 42518 11772 42524 11824
rect 42576 11812 42582 11824
rect 45830 11812 45836 11824
rect 42576 11784 45836 11812
rect 42576 11772 42582 11784
rect 45830 11772 45836 11784
rect 45888 11812 45894 11824
rect 49804 11821 49832 11852
rect 50706 11840 50712 11892
rect 50764 11840 50770 11892
rect 50982 11840 50988 11892
rect 51040 11880 51046 11892
rect 51040 11840 51074 11880
rect 48685 11815 48743 11821
rect 48685 11812 48697 11815
rect 45888 11784 48697 11812
rect 45888 11772 45894 11784
rect 48685 11781 48697 11784
rect 48731 11781 48743 11815
rect 49421 11815 49479 11821
rect 49421 11812 49433 11815
rect 48685 11775 48743 11781
rect 48976 11784 49433 11812
rect 47854 11704 47860 11756
rect 47912 11704 47918 11756
rect 47946 11704 47952 11756
rect 48004 11704 48010 11756
rect 48225 11747 48283 11753
rect 48225 11713 48237 11747
rect 48271 11713 48283 11747
rect 48225 11707 48283 11713
rect 48240 11676 48268 11707
rect 48498 11704 48504 11756
rect 48556 11704 48562 11756
rect 48590 11704 48596 11756
rect 48648 11704 48654 11756
rect 48866 11704 48872 11756
rect 48924 11704 48930 11756
rect 48314 11676 48320 11688
rect 40333 11648 48320 11676
rect 48314 11636 48320 11648
rect 48372 11636 48378 11688
rect 48608 11676 48636 11704
rect 48976 11685 49004 11784
rect 49421 11781 49433 11784
rect 49467 11781 49479 11815
rect 49421 11775 49479 11781
rect 49789 11815 49847 11821
rect 49789 11781 49801 11815
rect 49835 11781 49847 11815
rect 51046 11812 51074 11840
rect 52822 11812 52828 11824
rect 49789 11775 49847 11781
rect 50908 11784 52828 11812
rect 49145 11747 49203 11753
rect 49145 11713 49157 11747
rect 49191 11713 49203 11747
rect 49145 11707 49203 11713
rect 48961 11679 49019 11685
rect 48961 11676 48973 11679
rect 48608 11648 48973 11676
rect 48961 11645 48973 11648
rect 49007 11645 49019 11679
rect 48961 11639 49019 11645
rect 40126 11568 40132 11620
rect 40184 11568 40190 11620
rect 46566 11568 46572 11620
rect 46624 11608 46630 11620
rect 49160 11608 49188 11707
rect 49326 11704 49332 11756
rect 49384 11704 49390 11756
rect 49513 11747 49571 11753
rect 49513 11713 49525 11747
rect 49559 11744 49571 11747
rect 49694 11744 49700 11756
rect 49559 11716 49700 11744
rect 49559 11713 49571 11716
rect 49513 11707 49571 11713
rect 49694 11704 49700 11716
rect 49752 11704 49758 11756
rect 49970 11704 49976 11756
rect 50028 11744 50034 11756
rect 50908 11753 50936 11784
rect 52822 11772 52828 11784
rect 52880 11812 52886 11824
rect 54386 11812 54392 11824
rect 52880 11784 54392 11812
rect 52880 11772 52886 11784
rect 54386 11772 54392 11784
rect 54444 11772 54450 11824
rect 54938 11772 54944 11824
rect 54996 11772 55002 11824
rect 50065 11747 50123 11753
rect 50065 11744 50077 11747
rect 50028 11716 50077 11744
rect 50028 11704 50034 11716
rect 50065 11713 50077 11716
rect 50111 11713 50123 11747
rect 50065 11707 50123 11713
rect 50893 11747 50951 11753
rect 50893 11713 50905 11747
rect 50939 11713 50951 11747
rect 50893 11707 50951 11713
rect 50982 11704 50988 11756
rect 51040 11704 51046 11756
rect 51261 11747 51319 11753
rect 51261 11713 51273 11747
rect 51307 11744 51319 11747
rect 51721 11747 51779 11753
rect 51721 11744 51733 11747
rect 51307 11716 51733 11744
rect 51307 11713 51319 11716
rect 51261 11707 51319 11713
rect 51721 11713 51733 11716
rect 51767 11713 51779 11747
rect 51721 11707 51779 11713
rect 51994 11704 52000 11756
rect 52052 11744 52058 11756
rect 52270 11744 52276 11756
rect 52052 11716 52276 11744
rect 52052 11704 52058 11716
rect 52270 11704 52276 11716
rect 52328 11704 52334 11756
rect 53006 11704 53012 11756
rect 53064 11704 53070 11756
rect 54202 11704 54208 11756
rect 54260 11704 54266 11756
rect 49878 11636 49884 11688
rect 49936 11636 49942 11688
rect 52733 11679 52791 11685
rect 52733 11676 52745 11679
rect 52472 11648 52745 11676
rect 51994 11608 52000 11620
rect 46624 11580 48268 11608
rect 49160 11580 52000 11608
rect 46624 11568 46630 11580
rect 41690 11540 41696 11552
rect 40052 11512 41696 11540
rect 41690 11500 41696 11512
rect 41748 11500 41754 11552
rect 46934 11500 46940 11552
rect 46992 11540 46998 11552
rect 48130 11540 48136 11552
rect 46992 11512 48136 11540
rect 46992 11500 46998 11512
rect 48130 11500 48136 11512
rect 48188 11500 48194 11552
rect 48240 11540 48268 11580
rect 51994 11568 52000 11580
rect 52052 11568 52058 11620
rect 52472 11552 52500 11648
rect 52733 11645 52745 11648
rect 52779 11645 52791 11679
rect 52733 11639 52791 11645
rect 54478 11636 54484 11688
rect 54536 11636 54542 11688
rect 49789 11543 49847 11549
rect 49789 11540 49801 11543
rect 48240 11512 49801 11540
rect 49789 11509 49801 11512
rect 49835 11509 49847 11543
rect 49789 11503 49847 11509
rect 50249 11543 50307 11549
rect 50249 11509 50261 11543
rect 50295 11540 50307 11543
rect 51074 11540 51080 11552
rect 50295 11512 51080 11540
rect 50295 11509 50307 11512
rect 50249 11503 50307 11509
rect 51074 11500 51080 11512
rect 51132 11500 51138 11552
rect 51166 11500 51172 11552
rect 51224 11540 51230 11552
rect 51902 11540 51908 11552
rect 51224 11512 51908 11540
rect 51224 11500 51230 11512
rect 51902 11500 51908 11512
rect 51960 11500 51966 11552
rect 52454 11500 52460 11552
rect 52512 11500 52518 11552
rect 55030 11500 55036 11552
rect 55088 11540 55094 11552
rect 55953 11543 56011 11549
rect 55953 11540 55965 11543
rect 55088 11512 55965 11540
rect 55088 11500 55094 11512
rect 55953 11509 55965 11512
rect 55999 11509 56011 11543
rect 55953 11503 56011 11509
rect 1104 11450 78844 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 78844 11450
rect 1104 11376 78844 11398
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 19150 11336 19156 11348
rect 18923 11308 19156 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 19150 11296 19156 11308
rect 19208 11296 19214 11348
rect 22462 11296 22468 11348
rect 22520 11336 22526 11348
rect 23293 11339 23351 11345
rect 23293 11336 23305 11339
rect 22520 11308 23305 11336
rect 22520 11296 22526 11308
rect 23293 11305 23305 11308
rect 23339 11305 23351 11339
rect 23293 11299 23351 11305
rect 23382 11296 23388 11348
rect 23440 11336 23446 11348
rect 23477 11339 23535 11345
rect 23477 11336 23489 11339
rect 23440 11308 23489 11336
rect 23440 11296 23446 11308
rect 23477 11305 23489 11308
rect 23523 11305 23535 11339
rect 23477 11299 23535 11305
rect 24394 11296 24400 11348
rect 24452 11336 24458 11348
rect 24452 11308 26096 11336
rect 24452 11296 24458 11308
rect 22373 11271 22431 11277
rect 22373 11237 22385 11271
rect 22419 11268 22431 11271
rect 24026 11268 24032 11280
rect 22419 11240 24032 11268
rect 22419 11237 22431 11240
rect 22373 11231 22431 11237
rect 24026 11228 24032 11240
rect 24084 11228 24090 11280
rect 26068 11268 26096 11308
rect 26142 11296 26148 11348
rect 26200 11336 26206 11348
rect 26789 11339 26847 11345
rect 26789 11336 26801 11339
rect 26200 11308 26801 11336
rect 26200 11296 26206 11308
rect 26789 11305 26801 11308
rect 26835 11305 26847 11339
rect 26789 11299 26847 11305
rect 27798 11296 27804 11348
rect 27856 11296 27862 11348
rect 29730 11296 29736 11348
rect 29788 11296 29794 11348
rect 29822 11296 29828 11348
rect 29880 11336 29886 11348
rect 41782 11336 41788 11348
rect 29880 11308 41788 11336
rect 29880 11296 29886 11308
rect 41782 11296 41788 11308
rect 41840 11296 41846 11348
rect 42242 11296 42248 11348
rect 42300 11296 42306 11348
rect 43993 11339 44051 11345
rect 43993 11305 44005 11339
rect 44039 11336 44051 11339
rect 44174 11336 44180 11348
rect 44039 11308 44180 11336
rect 44039 11305 44051 11308
rect 43993 11299 44051 11305
rect 44174 11296 44180 11308
rect 44232 11296 44238 11348
rect 45646 11296 45652 11348
rect 45704 11336 45710 11348
rect 46290 11336 46296 11348
rect 45704 11308 46296 11336
rect 45704 11296 45710 11308
rect 46290 11296 46296 11308
rect 46348 11296 46354 11348
rect 48314 11296 48320 11348
rect 48372 11296 48378 11348
rect 49053 11339 49111 11345
rect 49053 11305 49065 11339
rect 49099 11336 49111 11339
rect 49694 11336 49700 11348
rect 49099 11308 49700 11336
rect 49099 11305 49111 11308
rect 49053 11299 49111 11305
rect 49694 11296 49700 11308
rect 49752 11296 49758 11348
rect 50982 11296 50988 11348
rect 51040 11336 51046 11348
rect 51353 11339 51411 11345
rect 51353 11336 51365 11339
rect 51040 11308 51365 11336
rect 51040 11296 51046 11308
rect 51353 11305 51365 11308
rect 51399 11305 51411 11339
rect 51353 11299 51411 11305
rect 52380 11308 54437 11336
rect 37461 11271 37519 11277
rect 26068 11240 33824 11268
rect 17126 11160 17132 11212
rect 17184 11160 17190 11212
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11200 17463 11203
rect 20530 11200 20536 11212
rect 17451 11172 20536 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 20530 11160 20536 11172
rect 20588 11160 20594 11212
rect 20625 11203 20683 11209
rect 20625 11169 20637 11203
rect 20671 11200 20683 11203
rect 21450 11200 21456 11212
rect 20671 11172 21456 11200
rect 20671 11169 20683 11172
rect 20625 11163 20683 11169
rect 21450 11160 21456 11172
rect 21508 11160 21514 11212
rect 22922 11160 22928 11212
rect 22980 11200 22986 11212
rect 24118 11200 24124 11212
rect 22980 11172 24124 11200
rect 22980 11160 22986 11172
rect 24118 11160 24124 11172
rect 24176 11200 24182 11212
rect 25501 11203 25559 11209
rect 25501 11200 25513 11203
rect 24176 11172 25513 11200
rect 24176 11160 24182 11172
rect 25501 11169 25513 11172
rect 25547 11200 25559 11203
rect 27614 11200 27620 11212
rect 25547 11172 27620 11200
rect 25547 11169 25559 11172
rect 25501 11163 25559 11169
rect 27614 11160 27620 11172
rect 27672 11160 27678 11212
rect 27890 11160 27896 11212
rect 27948 11160 27954 11212
rect 29454 11160 29460 11212
rect 29512 11200 29518 11212
rect 30282 11200 30288 11212
rect 29512 11172 30288 11200
rect 29512 11160 29518 11172
rect 30282 11160 30288 11172
rect 30340 11160 30346 11212
rect 22002 11092 22008 11144
rect 22060 11132 22066 11144
rect 22465 11135 22523 11141
rect 22465 11132 22477 11135
rect 22060 11104 22477 11132
rect 22060 11092 22066 11104
rect 22465 11101 22477 11104
rect 22511 11101 22523 11135
rect 24486 11132 24492 11144
rect 22465 11095 22523 11101
rect 23124 11104 24492 11132
rect 18690 11064 18696 11076
rect 18630 11036 18696 11064
rect 18690 11024 18696 11036
rect 18748 11064 18754 11076
rect 19061 11067 19119 11073
rect 19061 11064 19073 11067
rect 18748 11036 19073 11064
rect 18748 11024 18754 11036
rect 19061 11033 19073 11036
rect 19107 11064 19119 11067
rect 19242 11064 19248 11076
rect 19107 11036 19248 11064
rect 19107 11033 19119 11036
rect 19061 11027 19119 11033
rect 19242 11024 19248 11036
rect 19300 11024 19306 11076
rect 20898 11024 20904 11076
rect 20956 11024 20962 11076
rect 23124 11073 23152 11104
rect 24486 11092 24492 11104
rect 24544 11132 24550 11144
rect 25777 11135 25835 11141
rect 25777 11132 25789 11135
rect 24544 11104 25789 11132
rect 24544 11092 24550 11104
rect 25777 11101 25789 11104
rect 25823 11132 25835 11135
rect 26234 11132 26240 11144
rect 25823 11104 26240 11132
rect 25823 11101 25835 11104
rect 25777 11095 25835 11101
rect 26234 11092 26240 11104
rect 26292 11092 26298 11144
rect 26329 11135 26387 11141
rect 26329 11101 26341 11135
rect 26375 11101 26387 11135
rect 26329 11095 26387 11101
rect 23109 11067 23167 11073
rect 23109 11064 23121 11067
rect 22204 11036 23121 11064
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 22204 10996 22232 11036
rect 23109 11033 23121 11036
rect 23155 11033 23167 11067
rect 23109 11027 23167 11033
rect 23290 11024 23296 11076
rect 23348 11073 23354 11076
rect 23348 11067 23367 11073
rect 23355 11033 23367 11067
rect 24210 11064 24216 11076
rect 23348 11027 23367 11033
rect 23400 11036 24216 11064
rect 23348 11024 23354 11027
rect 20772 10968 22232 10996
rect 20772 10956 20778 10968
rect 22646 10956 22652 11008
rect 22704 10996 22710 11008
rect 23400 10996 23428 11036
rect 24210 11024 24216 11036
rect 24268 11064 24274 11076
rect 26344 11064 26372 11095
rect 26418 11092 26424 11144
rect 26476 11092 26482 11144
rect 26602 11092 26608 11144
rect 26660 11092 26666 11144
rect 27338 11092 27344 11144
rect 27396 11132 27402 11144
rect 27801 11135 27859 11141
rect 27801 11132 27813 11135
rect 27396 11104 27813 11132
rect 27396 11092 27402 11104
rect 27801 11101 27813 11104
rect 27847 11101 27859 11135
rect 27801 11095 27859 11101
rect 28166 11092 28172 11144
rect 28224 11132 28230 11144
rect 30101 11135 30159 11141
rect 28224 11104 28580 11132
rect 28224 11092 28230 11104
rect 26510 11064 26516 11076
rect 24268 11036 26516 11064
rect 24268 11024 24274 11036
rect 26510 11024 26516 11036
rect 26568 11024 26574 11076
rect 27246 11024 27252 11076
rect 27304 11064 27310 11076
rect 28261 11067 28319 11073
rect 28261 11064 28273 11067
rect 27304 11036 28273 11064
rect 27304 11024 27310 11036
rect 28261 11033 28273 11036
rect 28307 11033 28319 11067
rect 28261 11027 28319 11033
rect 28442 11024 28448 11076
rect 28500 11024 28506 11076
rect 28552 11064 28580 11104
rect 30101 11101 30113 11135
rect 30147 11132 30159 11135
rect 30653 11135 30711 11141
rect 30653 11132 30665 11135
rect 30147 11104 30665 11132
rect 30147 11101 30159 11104
rect 30101 11095 30159 11101
rect 30653 11101 30665 11104
rect 30699 11132 30711 11135
rect 31202 11132 31208 11144
rect 30699 11104 31208 11132
rect 30699 11101 30711 11104
rect 30653 11095 30711 11101
rect 31202 11092 31208 11104
rect 31260 11092 31266 11144
rect 30193 11067 30251 11073
rect 30193 11064 30205 11067
rect 28552 11036 30205 11064
rect 30193 11033 30205 11036
rect 30239 11033 30251 11067
rect 30193 11027 30251 11033
rect 22704 10968 23428 10996
rect 22704 10956 22710 10968
rect 26050 10956 26056 11008
rect 26108 10996 26114 11008
rect 26237 10999 26295 11005
rect 26237 10996 26249 10999
rect 26108 10968 26249 10996
rect 26108 10956 26114 10968
rect 26237 10965 26249 10968
rect 26283 10965 26295 10999
rect 26237 10959 26295 10965
rect 28166 10956 28172 11008
rect 28224 10956 28230 11008
rect 28626 10956 28632 11008
rect 28684 10956 28690 11008
rect 33796 10996 33824 11240
rect 37461 11237 37473 11271
rect 37507 11268 37519 11271
rect 37826 11268 37832 11280
rect 37507 11240 37832 11268
rect 37507 11237 37519 11240
rect 37461 11231 37519 11237
rect 37826 11228 37832 11240
rect 37884 11228 37890 11280
rect 39666 11228 39672 11280
rect 39724 11228 39730 11280
rect 34422 11160 34428 11212
rect 34480 11200 34486 11212
rect 35713 11203 35771 11209
rect 35713 11200 35725 11203
rect 34480 11172 35725 11200
rect 34480 11160 34486 11172
rect 35713 11169 35725 11172
rect 35759 11200 35771 11203
rect 37642 11200 37648 11212
rect 35759 11172 37648 11200
rect 35759 11169 35771 11172
rect 35713 11163 35771 11169
rect 37642 11160 37648 11172
rect 37700 11200 37706 11212
rect 37921 11203 37979 11209
rect 37921 11200 37933 11203
rect 37700 11172 37933 11200
rect 37700 11160 37706 11172
rect 37921 11169 37933 11172
rect 37967 11169 37979 11203
rect 37921 11163 37979 11169
rect 38194 11160 38200 11212
rect 38252 11160 38258 11212
rect 41782 11160 41788 11212
rect 41840 11200 41846 11212
rect 47854 11200 47860 11212
rect 41840 11172 43944 11200
rect 41840 11160 41846 11172
rect 42058 11092 42064 11144
rect 42116 11092 42122 11144
rect 42337 11135 42395 11141
rect 42337 11101 42349 11135
rect 42383 11132 42395 11135
rect 42981 11135 43039 11141
rect 42981 11132 42993 11135
rect 42383 11104 42993 11132
rect 42383 11101 42395 11104
rect 42337 11095 42395 11101
rect 42981 11101 42993 11104
rect 43027 11101 43039 11135
rect 42981 11095 43039 11101
rect 43346 11092 43352 11144
rect 43404 11132 43410 11144
rect 43916 11141 43944 11172
rect 44284 11172 47860 11200
rect 43533 11135 43591 11141
rect 43533 11132 43545 11135
rect 43404 11104 43545 11132
rect 43404 11092 43410 11104
rect 43533 11101 43545 11104
rect 43579 11101 43591 11135
rect 43533 11095 43591 11101
rect 43901 11135 43959 11141
rect 43901 11101 43913 11135
rect 43947 11101 43959 11135
rect 43901 11095 43959 11101
rect 35986 11024 35992 11076
rect 36044 11024 36050 11076
rect 37214 11036 38608 11064
rect 37458 10996 37464 11008
rect 33796 10968 37464 10996
rect 37458 10956 37464 10968
rect 37516 10956 37522 11008
rect 38580 10996 38608 11036
rect 38654 11024 38660 11076
rect 38712 11024 38718 11076
rect 43916 11064 43944 11095
rect 44174 11092 44180 11144
rect 44232 11092 44238 11144
rect 44284 11141 44312 11172
rect 47854 11160 47860 11172
rect 47912 11160 47918 11212
rect 48498 11160 48504 11212
rect 48556 11200 48562 11212
rect 50430 11200 50436 11212
rect 48556 11172 50436 11200
rect 48556 11160 48562 11172
rect 50430 11160 50436 11172
rect 50488 11200 50494 11212
rect 50488 11172 50568 11200
rect 50488 11160 50494 11172
rect 44269 11135 44327 11141
rect 44269 11101 44281 11135
rect 44315 11101 44327 11135
rect 44269 11095 44327 11101
rect 44818 11092 44824 11144
rect 44876 11132 44882 11144
rect 46566 11132 46572 11144
rect 44876 11104 46572 11132
rect 44876 11092 44882 11104
rect 46566 11092 46572 11104
rect 46624 11092 46630 11144
rect 48590 11092 48596 11144
rect 48648 11092 48654 11144
rect 50540 11132 50568 11172
rect 50614 11160 50620 11212
rect 50672 11200 50678 11212
rect 50890 11200 50896 11212
rect 50672 11172 50896 11200
rect 50672 11160 50678 11172
rect 50890 11160 50896 11172
rect 50948 11160 50954 11212
rect 52380 11200 52408 11308
rect 52549 11271 52607 11277
rect 52549 11237 52561 11271
rect 52595 11237 52607 11271
rect 54409 11268 54437 11308
rect 54478 11296 54484 11348
rect 54536 11296 54542 11348
rect 54941 11339 54999 11345
rect 54941 11305 54953 11339
rect 54987 11336 54999 11339
rect 55766 11336 55772 11348
rect 54987 11308 55772 11336
rect 54987 11305 54999 11308
rect 54941 11299 54999 11305
rect 54570 11268 54576 11280
rect 54409 11240 54576 11268
rect 52549 11231 52607 11237
rect 51552 11172 52408 11200
rect 52564 11200 52592 11231
rect 54570 11228 54576 11240
rect 54628 11228 54634 11280
rect 53101 11203 53159 11209
rect 52564 11172 52960 11200
rect 51552 11141 51580 11172
rect 51537 11135 51595 11141
rect 51537 11132 51549 11135
rect 50540 11104 51549 11132
rect 51537 11101 51549 11104
rect 51583 11101 51595 11135
rect 51537 11095 51595 11101
rect 51629 11135 51687 11141
rect 51629 11101 51641 11135
rect 51675 11101 51687 11135
rect 51629 11095 51687 11101
rect 44545 11067 44603 11073
rect 44545 11064 44557 11067
rect 43916 11036 44557 11064
rect 44545 11033 44557 11036
rect 44591 11064 44603 11067
rect 45373 11067 45431 11073
rect 45373 11064 45385 11067
rect 44591 11036 45385 11064
rect 44591 11033 44603 11036
rect 44545 11027 44603 11033
rect 45373 11033 45385 11036
rect 45419 11064 45431 11067
rect 45646 11064 45652 11076
rect 45419 11036 45652 11064
rect 45419 11033 45431 11036
rect 45373 11027 45431 11033
rect 45646 11024 45652 11036
rect 45704 11024 45710 11076
rect 48774 11024 48780 11076
rect 48832 11064 48838 11076
rect 49326 11064 49332 11076
rect 48832 11036 49332 11064
rect 48832 11024 48838 11036
rect 49326 11024 49332 11036
rect 49384 11024 49390 11076
rect 50890 11024 50896 11076
rect 50948 11064 50954 11076
rect 51644 11064 51672 11095
rect 51994 11092 52000 11144
rect 52052 11092 52058 11144
rect 52380 11141 52408 11172
rect 52273 11135 52331 11141
rect 52273 11132 52285 11135
rect 52104 11104 52285 11132
rect 51718 11064 51724 11076
rect 50948 11036 51724 11064
rect 50948 11024 50954 11036
rect 51718 11024 51724 11036
rect 51776 11024 51782 11076
rect 39022 10996 39028 11008
rect 38580 10968 39028 10996
rect 39022 10956 39028 10968
rect 39080 10956 39086 11008
rect 41877 10999 41935 11005
rect 41877 10965 41889 10999
rect 41923 10996 41935 10999
rect 41966 10996 41972 11008
rect 41923 10968 41972 10996
rect 41923 10965 41935 10968
rect 41877 10959 41935 10965
rect 41966 10956 41972 10968
rect 42024 10956 42030 11008
rect 42242 10956 42248 11008
rect 42300 10996 42306 11008
rect 42429 10999 42487 11005
rect 42429 10996 42441 10999
rect 42300 10968 42441 10996
rect 42300 10956 42306 10968
rect 42429 10965 42441 10968
rect 42475 10965 42487 10999
rect 42429 10959 42487 10965
rect 44266 10956 44272 11008
rect 44324 10996 44330 11008
rect 44453 10999 44511 11005
rect 44453 10996 44465 10999
rect 44324 10968 44465 10996
rect 44324 10956 44330 10968
rect 44453 10965 44465 10968
rect 44499 10965 44511 10999
rect 44453 10959 44511 10965
rect 45738 10956 45744 11008
rect 45796 10996 45802 11008
rect 45833 10999 45891 11005
rect 45833 10996 45845 10999
rect 45796 10968 45845 10996
rect 45796 10956 45802 10968
rect 45833 10965 45845 10968
rect 45879 10996 45891 10999
rect 46106 10996 46112 11008
rect 45879 10968 46112 10996
rect 45879 10965 45891 10968
rect 45833 10959 45891 10965
rect 46106 10956 46112 10968
rect 46164 10956 46170 11008
rect 50706 10956 50712 11008
rect 50764 10996 50770 11008
rect 52104 10996 52132 11104
rect 52273 11101 52285 11104
rect 52319 11101 52331 11135
rect 52273 11095 52331 11101
rect 52365 11135 52423 11141
rect 52365 11101 52377 11135
rect 52411 11101 52423 11135
rect 52365 11095 52423 11101
rect 52638 11092 52644 11144
rect 52696 11092 52702 11144
rect 52822 11092 52828 11144
rect 52880 11092 52886 11144
rect 52932 11141 52960 11172
rect 53101 11169 53113 11203
rect 53147 11200 53159 11203
rect 53558 11200 53564 11212
rect 53147 11172 53564 11200
rect 53147 11169 53159 11172
rect 53101 11163 53159 11169
rect 53558 11160 53564 11172
rect 53616 11200 53622 11212
rect 53616 11172 53788 11200
rect 53616 11160 53622 11172
rect 52917 11135 52975 11141
rect 52917 11101 52929 11135
rect 52963 11101 52975 11135
rect 52917 11095 52975 11101
rect 53193 11135 53251 11141
rect 53193 11101 53205 11135
rect 53239 11132 53251 11135
rect 53653 11135 53711 11141
rect 53653 11132 53665 11135
rect 53239 11104 53665 11132
rect 53239 11101 53251 11104
rect 53193 11095 53251 11101
rect 53653 11101 53665 11104
rect 53699 11101 53711 11135
rect 53760 11132 53788 11172
rect 54202 11160 54208 11212
rect 54260 11160 54266 11212
rect 54956 11200 54984 11299
rect 55766 11296 55772 11308
rect 55824 11296 55830 11348
rect 54312 11172 54984 11200
rect 54312 11132 54340 11172
rect 53760 11104 54340 11132
rect 53653 11095 53711 11101
rect 54386 11092 54392 11144
rect 54444 11132 54450 11144
rect 54665 11135 54723 11141
rect 54665 11132 54677 11135
rect 54444 11104 54677 11132
rect 54444 11092 54450 11104
rect 54665 11101 54677 11104
rect 54711 11101 54723 11135
rect 54665 11095 54723 11101
rect 52181 11067 52239 11073
rect 52181 11033 52193 11067
rect 52227 11064 52239 11067
rect 53006 11064 53012 11076
rect 52227 11036 53012 11064
rect 52227 11033 52239 11036
rect 52181 11027 52239 11033
rect 53006 11024 53012 11036
rect 53064 11064 53070 11076
rect 54294 11064 54300 11076
rect 53064 11036 54300 11064
rect 53064 11024 53070 11036
rect 54294 11024 54300 11036
rect 54352 11024 54358 11076
rect 54680 11064 54708 11095
rect 54754 11092 54760 11144
rect 54812 11092 54818 11144
rect 55030 11092 55036 11144
rect 55088 11092 55094 11144
rect 54938 11064 54944 11076
rect 54680 11036 54944 11064
rect 54938 11024 54944 11036
rect 54996 11024 55002 11076
rect 55030 10996 55036 11008
rect 50764 10968 55036 10996
rect 50764 10956 50770 10968
rect 55030 10956 55036 10968
rect 55088 10956 55094 11008
rect 1104 10906 78844 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 66314 10906
rect 66366 10854 66378 10906
rect 66430 10854 66442 10906
rect 66494 10854 66506 10906
rect 66558 10854 66570 10906
rect 66622 10854 78844 10906
rect 1104 10832 78844 10854
rect 19150 10752 19156 10804
rect 19208 10792 19214 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 19208 10764 19625 10792
rect 19208 10752 19214 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 19613 10755 19671 10761
rect 19705 10795 19763 10801
rect 19705 10761 19717 10795
rect 19751 10792 19763 10795
rect 19886 10792 19892 10804
rect 19751 10764 19892 10792
rect 19751 10761 19763 10764
rect 19705 10755 19763 10761
rect 19886 10752 19892 10764
rect 19944 10752 19950 10804
rect 32769 10795 32827 10801
rect 32769 10761 32781 10795
rect 32815 10792 32827 10795
rect 32950 10792 32956 10804
rect 32815 10764 32956 10792
rect 32815 10761 32827 10764
rect 32769 10755 32827 10761
rect 22002 10724 22008 10736
rect 20746 10696 22008 10724
rect 22002 10684 22008 10696
rect 22060 10684 22066 10736
rect 26970 10724 26976 10736
rect 26620 10696 26976 10724
rect 17126 10616 17132 10668
rect 17184 10656 17190 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17184 10628 17877 10656
rect 17184 10616 17190 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 19242 10616 19248 10668
rect 19300 10656 19306 10668
rect 19702 10656 19708 10668
rect 19300 10628 19708 10656
rect 19300 10616 19306 10628
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 25774 10616 25780 10668
rect 25832 10656 25838 10668
rect 26145 10659 26203 10665
rect 26145 10656 26157 10659
rect 25832 10628 26157 10656
rect 25832 10616 25838 10628
rect 26145 10625 26157 10628
rect 26191 10625 26203 10659
rect 26145 10619 26203 10625
rect 26326 10616 26332 10668
rect 26384 10616 26390 10668
rect 26620 10665 26648 10696
rect 26970 10684 26976 10696
rect 27028 10724 27034 10736
rect 32493 10727 32551 10733
rect 27028 10696 29592 10724
rect 27028 10684 27034 10696
rect 29564 10668 29592 10696
rect 32493 10693 32505 10727
rect 32539 10724 32551 10727
rect 32784 10724 32812 10755
rect 32950 10752 32956 10764
rect 33008 10752 33014 10804
rect 35986 10752 35992 10804
rect 36044 10792 36050 10804
rect 36265 10795 36323 10801
rect 36265 10792 36277 10795
rect 36044 10764 36277 10792
rect 36044 10752 36050 10764
rect 36265 10761 36277 10764
rect 36311 10761 36323 10795
rect 36265 10755 36323 10761
rect 38838 10752 38844 10804
rect 38896 10792 38902 10804
rect 39485 10795 39543 10801
rect 39485 10792 39497 10795
rect 38896 10764 39497 10792
rect 38896 10752 38902 10764
rect 39485 10761 39497 10764
rect 39531 10792 39543 10795
rect 39574 10792 39580 10804
rect 39531 10764 39580 10792
rect 39531 10761 39543 10764
rect 39485 10755 39543 10761
rect 39574 10752 39580 10764
rect 39632 10752 39638 10804
rect 42058 10752 42064 10804
rect 42116 10752 42122 10804
rect 43901 10795 43959 10801
rect 43901 10761 43913 10795
rect 43947 10792 43959 10795
rect 44174 10792 44180 10804
rect 43947 10764 44180 10792
rect 43947 10761 43959 10764
rect 43901 10755 43959 10761
rect 44174 10752 44180 10764
rect 44232 10752 44238 10804
rect 45646 10752 45652 10804
rect 45704 10792 45710 10804
rect 45741 10795 45799 10801
rect 45741 10792 45753 10795
rect 45704 10764 45753 10792
rect 45704 10752 45710 10764
rect 45741 10761 45753 10764
rect 45787 10792 45799 10795
rect 45787 10764 46244 10792
rect 45787 10761 45799 10764
rect 45741 10755 45799 10761
rect 33778 10724 33784 10736
rect 32539 10696 32812 10724
rect 33336 10696 33784 10724
rect 32539 10693 32551 10696
rect 32493 10687 32551 10693
rect 33336 10668 33364 10696
rect 33778 10684 33784 10696
rect 33836 10684 33842 10736
rect 34422 10684 34428 10736
rect 34480 10684 34486 10736
rect 38562 10724 38568 10736
rect 36648 10696 38568 10724
rect 26605 10659 26663 10665
rect 26605 10625 26617 10659
rect 26651 10625 26663 10659
rect 26605 10619 26663 10625
rect 28626 10616 28632 10668
rect 28684 10616 28690 10668
rect 28813 10659 28871 10665
rect 28813 10625 28825 10659
rect 28859 10656 28871 10659
rect 29454 10656 29460 10668
rect 28859 10628 29460 10656
rect 28859 10625 28871 10628
rect 28813 10619 28871 10625
rect 29454 10616 29460 10628
rect 29512 10616 29518 10668
rect 29546 10616 29552 10668
rect 29604 10616 29610 10668
rect 32950 10616 32956 10668
rect 33008 10616 33014 10668
rect 33137 10659 33195 10665
rect 33137 10625 33149 10659
rect 33183 10625 33195 10659
rect 33137 10619 33195 10625
rect 18141 10591 18199 10597
rect 18141 10557 18153 10591
rect 18187 10588 18199 10591
rect 20714 10588 20720 10600
rect 18187 10560 20720 10588
rect 18187 10557 18199 10560
rect 18141 10551 18199 10557
rect 20714 10548 20720 10560
rect 20772 10548 20778 10600
rect 21174 10548 21180 10600
rect 21232 10548 21238 10600
rect 21450 10548 21456 10600
rect 21508 10548 21514 10600
rect 28166 10548 28172 10600
rect 28224 10588 28230 10600
rect 28721 10591 28779 10597
rect 28721 10588 28733 10591
rect 28224 10560 28733 10588
rect 28224 10548 28230 10560
rect 28721 10557 28733 10560
rect 28767 10557 28779 10591
rect 28721 10551 28779 10557
rect 28905 10591 28963 10597
rect 28905 10557 28917 10591
rect 28951 10588 28963 10591
rect 29365 10591 29423 10597
rect 29365 10588 29377 10591
rect 28951 10560 29377 10588
rect 28951 10557 28963 10560
rect 28905 10551 28963 10557
rect 29365 10557 29377 10560
rect 29411 10557 29423 10591
rect 29365 10551 29423 10557
rect 29733 10591 29791 10597
rect 29733 10557 29745 10591
rect 29779 10588 29791 10591
rect 29822 10588 29828 10600
rect 29779 10560 29828 10588
rect 29779 10557 29791 10560
rect 29733 10551 29791 10557
rect 29822 10548 29828 10560
rect 29880 10548 29886 10600
rect 32122 10548 32128 10600
rect 32180 10588 32186 10600
rect 33152 10588 33180 10619
rect 33226 10616 33232 10668
rect 33284 10616 33290 10668
rect 33318 10616 33324 10668
rect 33376 10616 33382 10668
rect 36449 10659 36507 10665
rect 36449 10625 36461 10659
rect 36495 10656 36507 10659
rect 36538 10656 36544 10668
rect 36495 10628 36544 10656
rect 36495 10625 36507 10628
rect 36449 10619 36507 10625
rect 36538 10616 36544 10628
rect 36596 10616 36602 10668
rect 36648 10665 36676 10696
rect 38562 10684 38568 10696
rect 38620 10684 38626 10736
rect 38654 10684 38660 10736
rect 38712 10724 38718 10736
rect 39022 10724 39028 10736
rect 38712 10696 39028 10724
rect 38712 10684 38718 10696
rect 39022 10684 39028 10696
rect 39080 10684 39086 10736
rect 41690 10684 41696 10736
rect 41748 10724 41754 10736
rect 41748 10696 42748 10724
rect 41748 10684 41754 10696
rect 36633 10659 36691 10665
rect 36633 10625 36645 10659
rect 36679 10625 36691 10659
rect 36633 10619 36691 10625
rect 36725 10659 36783 10665
rect 36725 10625 36737 10659
rect 36771 10656 36783 10659
rect 37274 10656 37280 10668
rect 36771 10628 37280 10656
rect 36771 10625 36783 10628
rect 36725 10619 36783 10625
rect 37274 10616 37280 10628
rect 37332 10616 37338 10668
rect 37826 10616 37832 10668
rect 37884 10656 37890 10668
rect 38746 10656 38752 10668
rect 37884 10628 38752 10656
rect 37884 10616 37890 10628
rect 38746 10616 38752 10628
rect 38804 10656 38810 10668
rect 38841 10659 38899 10665
rect 38841 10656 38853 10659
rect 38804 10628 38853 10656
rect 38804 10616 38810 10628
rect 38841 10625 38853 10628
rect 38887 10625 38899 10659
rect 38841 10619 38899 10625
rect 41414 10616 41420 10668
rect 41472 10616 41478 10668
rect 41565 10659 41623 10665
rect 41565 10625 41577 10659
rect 41611 10656 41623 10659
rect 41611 10628 41736 10656
rect 41611 10625 41623 10628
rect 41565 10619 41623 10625
rect 41708 10600 41736 10628
rect 41782 10616 41788 10668
rect 41840 10616 41846 10668
rect 41923 10659 41981 10665
rect 41923 10625 41935 10659
rect 41969 10656 41981 10659
rect 42058 10656 42064 10668
rect 41969 10628 42064 10656
rect 41969 10625 41981 10628
rect 41923 10619 41981 10625
rect 42058 10616 42064 10628
rect 42116 10656 42122 10668
rect 42720 10665 42748 10696
rect 43272 10696 43760 10724
rect 42705 10659 42763 10665
rect 42116 10628 42656 10656
rect 42116 10616 42122 10628
rect 32180 10560 33180 10588
rect 32180 10548 32186 10560
rect 33594 10548 33600 10600
rect 33652 10548 33658 10600
rect 33870 10548 33876 10600
rect 33928 10548 33934 10600
rect 34882 10548 34888 10600
rect 34940 10588 34946 10600
rect 35345 10591 35403 10597
rect 35345 10588 35357 10591
rect 34940 10560 35357 10588
rect 34940 10548 34946 10560
rect 35345 10557 35357 10560
rect 35391 10557 35403 10591
rect 35345 10551 35403 10557
rect 37642 10548 37648 10600
rect 37700 10588 37706 10600
rect 38565 10591 38623 10597
rect 38565 10588 38577 10591
rect 37700 10560 38577 10588
rect 37700 10548 37706 10560
rect 38565 10557 38577 10560
rect 38611 10588 38623 10591
rect 40218 10588 40224 10600
rect 38611 10560 40224 10588
rect 38611 10557 38623 10560
rect 38565 10551 38623 10557
rect 40218 10548 40224 10560
rect 40276 10548 40282 10600
rect 41690 10548 41696 10600
rect 41748 10548 41754 10600
rect 41800 10588 41828 10616
rect 42153 10591 42211 10597
rect 42153 10588 42165 10591
rect 41800 10560 42165 10588
rect 42153 10557 42165 10560
rect 42199 10557 42211 10591
rect 42153 10551 42211 10557
rect 42242 10548 42248 10600
rect 42300 10588 42306 10600
rect 42429 10591 42487 10597
rect 42429 10588 42441 10591
rect 42300 10560 42441 10588
rect 42300 10548 42306 10560
rect 42429 10557 42441 10560
rect 42475 10557 42487 10591
rect 42628 10588 42656 10628
rect 42705 10625 42717 10659
rect 42751 10625 42763 10659
rect 42705 10619 42763 10625
rect 43272 10588 43300 10696
rect 43732 10668 43760 10696
rect 44266 10684 44272 10736
rect 44324 10684 44330 10736
rect 46216 10733 46244 10764
rect 48866 10752 48872 10804
rect 48924 10792 48930 10804
rect 49234 10792 49240 10804
rect 48924 10764 49240 10792
rect 48924 10752 48930 10764
rect 49234 10752 49240 10764
rect 49292 10792 49298 10804
rect 49329 10795 49387 10801
rect 49329 10792 49341 10795
rect 49292 10764 49341 10792
rect 49292 10752 49298 10764
rect 49329 10761 49341 10764
rect 49375 10761 49387 10795
rect 49329 10755 49387 10761
rect 50249 10795 50307 10801
rect 50249 10761 50261 10795
rect 50295 10792 50307 10795
rect 51350 10792 51356 10804
rect 50295 10764 51356 10792
rect 50295 10761 50307 10764
rect 50249 10755 50307 10761
rect 46201 10727 46259 10733
rect 46201 10693 46213 10727
rect 46247 10693 46259 10727
rect 46201 10687 46259 10693
rect 46290 10684 46296 10736
rect 46348 10684 46354 10736
rect 46658 10684 46664 10736
rect 46716 10724 46722 10736
rect 46716 10696 48346 10724
rect 46716 10684 46722 10696
rect 43346 10616 43352 10668
rect 43404 10616 43410 10668
rect 43533 10659 43591 10665
rect 43533 10625 43545 10659
rect 43579 10625 43591 10659
rect 43533 10619 43591 10625
rect 42628 10560 43300 10588
rect 43548 10588 43576 10619
rect 43622 10616 43628 10668
rect 43680 10616 43686 10668
rect 43714 10616 43720 10668
rect 43772 10616 43778 10668
rect 46106 10665 46112 10668
rect 46104 10656 46112 10665
rect 43548 10560 43668 10588
rect 42429 10551 42487 10557
rect 21637 10455 21695 10461
rect 21637 10421 21649 10455
rect 21683 10452 21695 10455
rect 22002 10452 22008 10464
rect 21683 10424 22008 10452
rect 21683 10421 21695 10424
rect 21637 10415 21695 10421
rect 22002 10412 22008 10424
rect 22060 10412 22066 10464
rect 26602 10412 26608 10464
rect 26660 10452 26666 10464
rect 26789 10455 26847 10461
rect 26789 10452 26801 10455
rect 26660 10424 26801 10452
rect 26660 10412 26666 10424
rect 26789 10421 26801 10424
rect 26835 10421 26847 10455
rect 26789 10415 26847 10421
rect 28442 10412 28448 10464
rect 28500 10412 28506 10464
rect 32398 10412 32404 10464
rect 32456 10412 32462 10464
rect 33505 10455 33563 10461
rect 33505 10421 33517 10455
rect 33551 10452 33563 10455
rect 34606 10452 34612 10464
rect 33551 10424 34612 10452
rect 33551 10421 33563 10424
rect 33505 10415 33563 10421
rect 34606 10412 34612 10424
rect 34664 10412 34670 10464
rect 43640 10452 43668 10560
rect 43990 10548 43996 10600
rect 44048 10548 44054 10600
rect 45388 10588 45416 10642
rect 46067 10628 46112 10656
rect 46104 10619 46112 10628
rect 46106 10616 46112 10619
rect 46164 10616 46170 10668
rect 46476 10659 46534 10665
rect 46476 10625 46488 10659
rect 46522 10625 46534 10659
rect 46476 10619 46534 10625
rect 46492 10588 46520 10619
rect 46566 10616 46572 10668
rect 46624 10616 46630 10668
rect 47118 10616 47124 10668
rect 47176 10656 47182 10668
rect 47581 10659 47639 10665
rect 47581 10656 47593 10659
rect 47176 10628 47593 10656
rect 47176 10616 47182 10628
rect 47581 10625 47593 10628
rect 47627 10625 47639 10659
rect 49344 10656 49372 10755
rect 51350 10752 51356 10764
rect 51408 10752 51414 10804
rect 51718 10752 51724 10804
rect 51776 10792 51782 10804
rect 51776 10764 53512 10792
rect 51776 10752 51782 10764
rect 50798 10684 50804 10736
rect 50856 10724 50862 10736
rect 51442 10724 51448 10736
rect 50856 10696 51448 10724
rect 50856 10684 50862 10696
rect 51442 10684 51448 10696
rect 51500 10684 51506 10736
rect 51810 10684 51816 10736
rect 51868 10684 51874 10736
rect 49973 10659 50031 10665
rect 49973 10656 49985 10659
rect 49344 10628 49985 10656
rect 47581 10619 47639 10625
rect 49973 10625 49985 10628
rect 50019 10625 50031 10659
rect 49973 10619 50031 10625
rect 51077 10659 51135 10665
rect 51077 10625 51089 10659
rect 51123 10656 51135 10659
rect 53098 10656 53104 10668
rect 51123 10628 53104 10656
rect 51123 10625 51135 10628
rect 51077 10619 51135 10625
rect 47026 10588 47032 10600
rect 45388 10560 46428 10588
rect 46492 10560 47032 10588
rect 45278 10480 45284 10532
rect 45336 10520 45342 10532
rect 45925 10523 45983 10529
rect 45925 10520 45937 10523
rect 45336 10492 45937 10520
rect 45336 10480 45342 10492
rect 45925 10489 45937 10492
rect 45971 10489 45983 10523
rect 46400 10520 46428 10560
rect 47026 10548 47032 10560
rect 47084 10548 47090 10600
rect 47857 10591 47915 10597
rect 47857 10557 47869 10591
rect 47903 10588 47915 10591
rect 47946 10588 47952 10600
rect 47903 10560 47952 10588
rect 47903 10557 47915 10560
rect 47857 10551 47915 10557
rect 47946 10548 47952 10560
rect 48004 10548 48010 10600
rect 49418 10548 49424 10600
rect 49476 10588 49482 10600
rect 49476 10560 49648 10588
rect 49476 10548 49482 10560
rect 46661 10523 46719 10529
rect 46661 10520 46673 10523
rect 46400 10492 46673 10520
rect 45925 10483 45983 10489
rect 46661 10489 46673 10492
rect 46707 10489 46719 10523
rect 46661 10483 46719 10489
rect 44266 10452 44272 10464
rect 43640 10424 44272 10452
rect 44266 10412 44272 10424
rect 44324 10412 44330 10464
rect 46676 10452 46704 10483
rect 49620 10464 49648 10560
rect 48222 10452 48228 10464
rect 46676 10424 48228 10452
rect 48222 10412 48228 10424
rect 48280 10412 48286 10464
rect 49418 10412 49424 10464
rect 49476 10412 49482 10464
rect 49602 10412 49608 10464
rect 49660 10452 49666 10464
rect 50341 10455 50399 10461
rect 50341 10452 50353 10455
rect 49660 10424 50353 10452
rect 49660 10412 49666 10424
rect 50341 10421 50353 10424
rect 50387 10452 50399 10455
rect 50798 10452 50804 10464
rect 50387 10424 50804 10452
rect 50387 10421 50399 10424
rect 50341 10415 50399 10421
rect 50798 10412 50804 10424
rect 50856 10412 50862 10464
rect 50985 10455 51043 10461
rect 50985 10421 50997 10455
rect 51031 10452 51043 10455
rect 51092 10452 51120 10619
rect 53098 10616 53104 10628
rect 53156 10656 53162 10668
rect 53374 10656 53380 10668
rect 53156 10628 53380 10656
rect 53156 10616 53162 10628
rect 53374 10616 53380 10628
rect 53432 10616 53438 10668
rect 53484 10656 53512 10764
rect 54754 10752 54760 10804
rect 54812 10752 54818 10804
rect 54294 10684 54300 10736
rect 54352 10724 54358 10736
rect 54389 10727 54447 10733
rect 54389 10724 54401 10727
rect 54352 10696 54401 10724
rect 54352 10684 54358 10696
rect 54389 10693 54401 10696
rect 54435 10693 54447 10727
rect 54389 10687 54447 10693
rect 54202 10656 54208 10668
rect 53484 10628 54208 10656
rect 54202 10616 54208 10628
rect 54260 10616 54266 10668
rect 54481 10659 54539 10665
rect 54481 10625 54493 10659
rect 54527 10625 54539 10659
rect 54481 10619 54539 10625
rect 52086 10548 52092 10600
rect 52144 10588 52150 10600
rect 54496 10588 54524 10619
rect 54570 10616 54576 10668
rect 54628 10616 54634 10668
rect 56594 10588 56600 10600
rect 52144 10560 56600 10588
rect 52144 10548 52150 10560
rect 56594 10548 56600 10560
rect 56652 10548 56658 10600
rect 51031 10424 51120 10452
rect 51031 10421 51043 10424
rect 50985 10415 51043 10421
rect 54846 10412 54852 10464
rect 54904 10452 54910 10464
rect 55766 10452 55772 10464
rect 54904 10424 55772 10452
rect 54904 10412 54910 10424
rect 55766 10412 55772 10424
rect 55824 10412 55830 10464
rect 1104 10362 78844 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 78844 10362
rect 1104 10288 78844 10310
rect 25406 10208 25412 10260
rect 25464 10248 25470 10260
rect 30098 10248 30104 10260
rect 25464 10220 30104 10248
rect 25464 10208 25470 10220
rect 30098 10208 30104 10220
rect 30156 10208 30162 10260
rect 32674 10208 32680 10260
rect 32732 10248 32738 10260
rect 32769 10251 32827 10257
rect 32769 10248 32781 10251
rect 32732 10220 32781 10248
rect 32732 10208 32738 10220
rect 32769 10217 32781 10220
rect 32815 10217 32827 10251
rect 32769 10211 32827 10217
rect 32950 10208 32956 10260
rect 33008 10208 33014 10260
rect 33870 10208 33876 10260
rect 33928 10208 33934 10260
rect 39666 10208 39672 10260
rect 39724 10208 39730 10260
rect 43346 10208 43352 10260
rect 43404 10248 43410 10260
rect 43530 10248 43536 10260
rect 43404 10220 43536 10248
rect 43404 10208 43410 10220
rect 43530 10208 43536 10220
rect 43588 10208 43594 10260
rect 47946 10208 47952 10260
rect 48004 10208 48010 10260
rect 48130 10208 48136 10260
rect 48188 10248 48194 10260
rect 48409 10251 48467 10257
rect 48409 10248 48421 10251
rect 48188 10220 48421 10248
rect 48188 10208 48194 10220
rect 48409 10217 48421 10220
rect 48455 10217 48467 10251
rect 48409 10211 48467 10217
rect 48593 10251 48651 10257
rect 48593 10217 48605 10251
rect 48639 10217 48651 10251
rect 48593 10211 48651 10217
rect 39485 10183 39543 10189
rect 39485 10149 39497 10183
rect 39531 10180 39543 10183
rect 39758 10180 39764 10192
rect 39531 10152 39764 10180
rect 39531 10149 39543 10152
rect 39485 10143 39543 10149
rect 21450 10072 21456 10124
rect 21508 10112 21514 10124
rect 26329 10115 26387 10121
rect 26329 10112 26341 10115
rect 21508 10084 26341 10112
rect 21508 10072 21514 10084
rect 26329 10081 26341 10084
rect 26375 10112 26387 10115
rect 26510 10112 26516 10124
rect 26375 10084 26516 10112
rect 26375 10081 26387 10084
rect 26329 10075 26387 10081
rect 26510 10072 26516 10084
rect 26568 10072 26574 10124
rect 32677 10115 32735 10121
rect 32677 10081 32689 10115
rect 32723 10081 32735 10115
rect 32677 10075 32735 10081
rect 25406 10004 25412 10056
rect 25464 10044 25470 10056
rect 25593 10047 25651 10053
rect 25593 10044 25605 10047
rect 25464 10016 25605 10044
rect 25464 10004 25470 10016
rect 25593 10013 25605 10016
rect 25639 10013 25651 10047
rect 25593 10007 25651 10013
rect 26602 10004 26608 10056
rect 26660 10004 26666 10056
rect 26786 10004 26792 10056
rect 26844 10004 26850 10056
rect 26970 10004 26976 10056
rect 27028 10004 27034 10056
rect 30926 10004 30932 10056
rect 30984 10004 30990 10056
rect 32490 10004 32496 10056
rect 32548 10044 32554 10056
rect 32692 10044 32720 10075
rect 34606 10072 34612 10124
rect 34664 10112 34670 10124
rect 35253 10115 35311 10121
rect 35253 10112 35265 10115
rect 34664 10084 35265 10112
rect 34664 10072 34670 10084
rect 35253 10081 35265 10084
rect 35299 10081 35311 10115
rect 39500 10112 39528 10143
rect 39758 10140 39764 10152
rect 39816 10140 39822 10192
rect 48608 10180 48636 10211
rect 48682 10208 48688 10260
rect 48740 10248 48746 10260
rect 49326 10248 49332 10260
rect 48740 10220 49332 10248
rect 48740 10208 48746 10220
rect 49326 10208 49332 10220
rect 49384 10248 49390 10260
rect 50062 10248 50068 10260
rect 49384 10220 50068 10248
rect 49384 10208 49390 10220
rect 50062 10208 50068 10220
rect 50120 10248 50126 10260
rect 50157 10251 50215 10257
rect 50157 10248 50169 10251
rect 50120 10220 50169 10248
rect 50120 10208 50126 10220
rect 50157 10217 50169 10220
rect 50203 10217 50215 10251
rect 50157 10211 50215 10217
rect 51810 10208 51816 10260
rect 51868 10248 51874 10260
rect 51868 10220 52408 10248
rect 51868 10208 51874 10220
rect 48240 10152 48636 10180
rect 35253 10075 35311 10081
rect 39040 10084 39528 10112
rect 33042 10044 33048 10056
rect 32548 10016 33048 10044
rect 32548 10004 32554 10016
rect 33042 10004 33048 10016
rect 33100 10044 33106 10056
rect 33505 10047 33563 10053
rect 33505 10044 33517 10047
rect 33100 10016 33517 10044
rect 33100 10004 33106 10016
rect 33505 10013 33517 10016
rect 33551 10013 33563 10047
rect 33505 10007 33563 10013
rect 34514 10004 34520 10056
rect 34572 10004 34578 10056
rect 38838 10053 38844 10056
rect 38836 10044 38844 10053
rect 38799 10016 38844 10044
rect 38836 10007 38844 10016
rect 38838 10004 38844 10007
rect 38896 10004 38902 10056
rect 39040 10053 39068 10084
rect 39850 10072 39856 10124
rect 39908 10112 39914 10124
rect 39945 10115 40003 10121
rect 39945 10112 39957 10115
rect 39908 10084 39957 10112
rect 39908 10072 39914 10084
rect 39945 10081 39957 10084
rect 39991 10112 40003 10115
rect 40218 10112 40224 10124
rect 39991 10084 40224 10112
rect 39991 10081 40003 10084
rect 39945 10075 40003 10081
rect 40218 10072 40224 10084
rect 40276 10112 40282 10124
rect 41785 10115 41843 10121
rect 41785 10112 41797 10115
rect 40276 10084 41797 10112
rect 40276 10072 40282 10084
rect 41785 10081 41797 10084
rect 41831 10112 41843 10115
rect 43990 10112 43996 10124
rect 41831 10084 43996 10112
rect 41831 10081 41843 10084
rect 41785 10075 41843 10081
rect 43990 10072 43996 10084
rect 44048 10072 44054 10124
rect 45281 10115 45339 10121
rect 45281 10081 45293 10115
rect 45327 10112 45339 10115
rect 46934 10112 46940 10124
rect 45327 10084 46940 10112
rect 45327 10081 45339 10084
rect 45281 10075 45339 10081
rect 46934 10072 46940 10084
rect 46992 10072 46998 10124
rect 47026 10072 47032 10124
rect 47084 10072 47090 10124
rect 47210 10072 47216 10124
rect 47268 10112 47274 10124
rect 47854 10112 47860 10124
rect 47268 10084 47860 10112
rect 47268 10072 47274 10084
rect 47854 10072 47860 10084
rect 47912 10112 47918 10124
rect 47912 10084 48176 10112
rect 47912 10072 47918 10084
rect 39025 10047 39083 10053
rect 39025 10013 39037 10047
rect 39071 10013 39083 10047
rect 39206 10044 39212 10056
rect 39167 10016 39212 10044
rect 39025 10007 39083 10013
rect 39206 10004 39212 10016
rect 39264 10004 39270 10056
rect 39301 10047 39359 10053
rect 39301 10013 39313 10047
rect 39347 10044 39359 10047
rect 39666 10044 39672 10056
rect 39347 10016 39672 10044
rect 39347 10013 39359 10016
rect 39301 10007 39359 10013
rect 39666 10004 39672 10016
rect 39724 10004 39730 10056
rect 43346 10004 43352 10056
rect 43404 10044 43410 10056
rect 43809 10047 43867 10053
rect 43809 10044 43821 10047
rect 43404 10016 43821 10044
rect 43404 10004 43410 10016
rect 43809 10013 43821 10016
rect 43855 10044 43867 10047
rect 43898 10044 43904 10056
rect 43855 10016 43904 10044
rect 43855 10013 43867 10016
rect 43809 10007 43867 10013
rect 43898 10004 43904 10016
rect 43956 10044 43962 10056
rect 44085 10047 44143 10053
rect 44085 10044 44097 10047
rect 43956 10016 44097 10044
rect 43956 10004 43962 10016
rect 44085 10013 44097 10016
rect 44131 10013 44143 10047
rect 47044 10044 47072 10072
rect 47670 10044 47676 10056
rect 47044 10016 47676 10044
rect 44085 10007 44143 10013
rect 47670 10004 47676 10016
rect 47728 10004 47734 10056
rect 48148 10053 48176 10084
rect 48240 10053 48268 10152
rect 48866 10140 48872 10192
rect 48924 10180 48930 10192
rect 49881 10183 49939 10189
rect 49881 10180 49893 10183
rect 48924 10152 49893 10180
rect 48924 10140 48930 10152
rect 49418 10112 49424 10124
rect 48516 10084 49424 10112
rect 48516 10053 48544 10084
rect 49418 10072 49424 10084
rect 49476 10072 49482 10124
rect 48133 10047 48191 10053
rect 48133 10013 48145 10047
rect 48179 10013 48191 10047
rect 48133 10007 48191 10013
rect 48225 10047 48283 10053
rect 48225 10013 48237 10047
rect 48271 10013 48283 10047
rect 48225 10007 48283 10013
rect 48501 10047 48559 10053
rect 48501 10013 48513 10047
rect 48547 10013 48559 10047
rect 48501 10007 48559 10013
rect 48590 10004 48596 10056
rect 48648 10044 48654 10056
rect 48777 10047 48835 10053
rect 48777 10044 48789 10047
rect 48648 10016 48789 10044
rect 48648 10004 48654 10016
rect 48777 10013 48789 10016
rect 48823 10013 48835 10047
rect 48777 10007 48835 10013
rect 48866 10004 48872 10056
rect 48924 10004 48930 10056
rect 49145 10047 49203 10053
rect 49145 10013 49157 10047
rect 49191 10013 49203 10047
rect 49145 10007 49203 10013
rect 26878 9936 26884 9988
rect 26936 9936 26942 9988
rect 31202 9936 31208 9988
rect 31260 9936 31266 9988
rect 32674 9976 32680 9988
rect 32430 9948 32680 9976
rect 32674 9936 32680 9948
rect 32732 9936 32738 9988
rect 34790 9936 34796 9988
rect 34848 9976 34854 9988
rect 38933 9979 38991 9985
rect 38933 9976 38945 9979
rect 34848 9948 38945 9976
rect 34848 9936 34854 9948
rect 38933 9945 38945 9948
rect 38979 9945 38991 9979
rect 38933 9939 38991 9945
rect 40218 9936 40224 9988
rect 40276 9936 40282 9988
rect 41446 9948 41828 9976
rect 19702 9868 19708 9920
rect 19760 9868 19766 9920
rect 27154 9868 27160 9920
rect 27212 9868 27218 9920
rect 33870 9868 33876 9920
rect 33928 9908 33934 9920
rect 34330 9908 34336 9920
rect 33928 9880 34336 9908
rect 33928 9868 33934 9880
rect 34330 9868 34336 9880
rect 34388 9868 34394 9920
rect 34698 9868 34704 9920
rect 34756 9868 34762 9920
rect 37274 9868 37280 9920
rect 37332 9908 37338 9920
rect 38657 9911 38715 9917
rect 38657 9908 38669 9911
rect 37332 9880 38669 9908
rect 37332 9868 37338 9880
rect 38657 9877 38669 9880
rect 38703 9877 38715 9911
rect 38657 9871 38715 9877
rect 41230 9868 41236 9920
rect 41288 9908 41294 9920
rect 41524 9908 41552 9948
rect 41288 9880 41552 9908
rect 41288 9868 41294 9880
rect 41690 9868 41696 9920
rect 41748 9868 41754 9920
rect 41800 9908 41828 9948
rect 41966 9936 41972 9988
rect 42024 9976 42030 9988
rect 42061 9979 42119 9985
rect 42061 9976 42073 9979
rect 42024 9948 42073 9976
rect 42024 9936 42030 9948
rect 42061 9945 42073 9948
rect 42107 9945 42119 9979
rect 43993 9979 44051 9985
rect 42061 9939 42119 9945
rect 42168 9948 42550 9976
rect 42168 9908 42196 9948
rect 43993 9945 44005 9979
rect 44039 9976 44051 9979
rect 44266 9976 44272 9988
rect 44039 9948 44272 9976
rect 44039 9945 44051 9948
rect 43993 9939 44051 9945
rect 44266 9936 44272 9948
rect 44324 9976 44330 9988
rect 45186 9976 45192 9988
rect 44324 9948 45192 9976
rect 44324 9936 44330 9948
rect 45186 9936 45192 9948
rect 45244 9976 45250 9988
rect 45244 9948 45416 9976
rect 45244 9936 45250 9948
rect 41800 9880 42196 9908
rect 45388 9908 45416 9948
rect 45554 9936 45560 9988
rect 45612 9936 45618 9988
rect 46566 9936 46572 9988
rect 46624 9936 46630 9988
rect 46860 9948 47256 9976
rect 46860 9908 46888 9948
rect 45388 9880 46888 9908
rect 47118 9868 47124 9920
rect 47176 9868 47182 9920
rect 47228 9908 47256 9948
rect 48314 9936 48320 9988
rect 48372 9976 48378 9988
rect 48884 9976 48912 10004
rect 48372 9948 48912 9976
rect 48961 9979 49019 9985
rect 48372 9936 48378 9948
rect 48961 9945 48973 9979
rect 49007 9945 49019 9979
rect 48961 9939 49019 9945
rect 48976 9908 49004 9939
rect 47228 9880 49004 9908
rect 49160 9908 49188 10007
rect 49234 10004 49240 10056
rect 49292 10004 49298 10056
rect 49528 10053 49556 10152
rect 49881 10149 49893 10152
rect 49927 10149 49939 10183
rect 51350 10180 51356 10192
rect 49881 10143 49939 10149
rect 51046 10152 51356 10180
rect 49896 10112 49924 10143
rect 50154 10112 50160 10124
rect 49896 10084 50160 10112
rect 50154 10072 50160 10084
rect 50212 10072 50218 10124
rect 51046 10112 51074 10152
rect 51350 10140 51356 10152
rect 51408 10140 51414 10192
rect 51626 10140 51632 10192
rect 51684 10140 51690 10192
rect 51994 10180 52000 10192
rect 51920 10152 52000 10180
rect 51644 10112 51672 10140
rect 50632 10084 51074 10112
rect 51271 10084 51672 10112
rect 49513 10047 49571 10053
rect 49513 10013 49525 10047
rect 49559 10013 49571 10047
rect 49513 10007 49571 10013
rect 49605 10047 49663 10053
rect 49605 10013 49617 10047
rect 49651 10044 49663 10047
rect 49970 10044 49976 10056
rect 49651 10016 49976 10044
rect 49651 10013 49663 10016
rect 49605 10007 49663 10013
rect 49970 10004 49976 10016
rect 50028 10004 50034 10056
rect 50338 10004 50344 10056
rect 50396 10004 50402 10056
rect 50430 10004 50436 10056
rect 50488 10044 50494 10056
rect 50632 10053 50660 10084
rect 51271 10056 51299 10084
rect 50617 10047 50675 10053
rect 50488 10016 50533 10044
rect 50488 10004 50494 10016
rect 50617 10013 50629 10047
rect 50663 10013 50675 10047
rect 50617 10007 50675 10013
rect 50706 10004 50712 10056
rect 50764 10004 50770 10056
rect 50798 10004 50804 10056
rect 50856 10053 50862 10056
rect 51258 10053 51264 10056
rect 50856 10044 50864 10053
rect 50856 10016 50901 10044
rect 50856 10007 50864 10016
rect 51256 10007 51264 10053
rect 50856 10004 50862 10007
rect 51258 10004 51264 10007
rect 51316 10004 51322 10056
rect 51442 10004 51448 10056
rect 51500 10004 51506 10056
rect 51534 10004 51540 10056
rect 51592 10053 51598 10056
rect 51592 10047 51631 10053
rect 51619 10013 51631 10047
rect 51592 10007 51631 10013
rect 51592 10004 51598 10007
rect 51718 10004 51724 10056
rect 51776 10004 51782 10056
rect 51920 10053 51948 10152
rect 51994 10140 52000 10152
rect 52052 10180 52058 10192
rect 52178 10180 52184 10192
rect 52052 10152 52184 10180
rect 52052 10140 52058 10152
rect 52178 10140 52184 10152
rect 52236 10140 52242 10192
rect 52380 10112 52408 10220
rect 52641 10115 52699 10121
rect 52641 10112 52653 10115
rect 52380 10084 52653 10112
rect 52641 10081 52653 10084
rect 52687 10112 52699 10115
rect 55309 10115 55367 10121
rect 55309 10112 55321 10115
rect 52687 10084 55321 10112
rect 52687 10081 52699 10084
rect 52641 10075 52699 10081
rect 55309 10081 55321 10084
rect 55355 10081 55367 10115
rect 55309 10075 55367 10081
rect 56594 10072 56600 10124
rect 56652 10112 56658 10124
rect 57057 10115 57115 10121
rect 57057 10112 57069 10115
rect 56652 10084 57069 10112
rect 56652 10072 56658 10084
rect 57057 10081 57069 10084
rect 57103 10081 57115 10115
rect 57057 10075 57115 10081
rect 51905 10047 51963 10053
rect 51905 10013 51917 10047
rect 51951 10013 51963 10047
rect 51905 10007 51963 10013
rect 51998 10047 52056 10053
rect 51998 10013 52010 10047
rect 52044 10044 52056 10047
rect 52086 10044 52092 10056
rect 52044 10016 52092 10044
rect 52044 10013 52056 10016
rect 51998 10007 52056 10013
rect 49326 9936 49332 9988
rect 49384 9976 49390 9988
rect 49421 9979 49479 9985
rect 49421 9976 49433 9979
rect 49384 9948 49433 9976
rect 49384 9936 49390 9948
rect 49421 9945 49433 9948
rect 49467 9945 49479 9979
rect 49421 9939 49479 9945
rect 51353 9979 51411 9985
rect 51353 9945 51365 9979
rect 51399 9976 51411 9979
rect 52012 9976 52040 10007
rect 52086 10004 52092 10016
rect 52144 10004 52150 10056
rect 52362 10004 52368 10056
rect 52420 10053 52426 10056
rect 52420 10044 52428 10053
rect 54846 10044 54852 10056
rect 52420 10016 52465 10044
rect 54050 10016 54852 10044
rect 52420 10007 52428 10016
rect 52420 10004 52426 10007
rect 54846 10004 54852 10016
rect 54904 10004 54910 10056
rect 55033 10047 55091 10053
rect 55033 10044 55045 10047
rect 54956 10016 55045 10044
rect 51399 9948 52040 9976
rect 51399 9945 51411 9948
rect 51353 9939 51411 9945
rect 52178 9936 52184 9988
rect 52236 9936 52242 9988
rect 52273 9979 52331 9985
rect 52273 9945 52285 9979
rect 52319 9945 52331 9979
rect 52273 9939 52331 9945
rect 49694 9908 49700 9920
rect 49160 9880 49700 9908
rect 49694 9868 49700 9880
rect 49752 9868 49758 9920
rect 49786 9868 49792 9920
rect 49844 9868 49850 9920
rect 50982 9868 50988 9920
rect 51040 9868 51046 9920
rect 51077 9911 51135 9917
rect 51077 9877 51089 9911
rect 51123 9908 51135 9911
rect 51258 9908 51264 9920
rect 51123 9880 51264 9908
rect 51123 9877 51135 9880
rect 51077 9871 51135 9877
rect 51258 9868 51264 9880
rect 51316 9868 51322 9920
rect 51442 9868 51448 9920
rect 51500 9908 51506 9920
rect 52288 9908 52316 9939
rect 52914 9936 52920 9988
rect 52972 9936 52978 9988
rect 54202 9936 54208 9988
rect 54260 9976 54266 9988
rect 54481 9979 54539 9985
rect 54481 9976 54493 9979
rect 54260 9948 54493 9976
rect 54260 9936 54266 9948
rect 54481 9945 54493 9948
rect 54527 9945 54539 9979
rect 54481 9939 54539 9945
rect 51500 9880 52316 9908
rect 52549 9911 52607 9917
rect 51500 9868 51506 9880
rect 52549 9877 52561 9911
rect 52595 9908 52607 9911
rect 53006 9908 53012 9920
rect 52595 9880 53012 9908
rect 52595 9877 52607 9880
rect 52549 9871 52607 9877
rect 53006 9868 53012 9880
rect 53064 9868 53070 9920
rect 54386 9868 54392 9920
rect 54444 9908 54450 9920
rect 54956 9908 54984 10016
rect 55033 10013 55045 10016
rect 55079 10013 55091 10047
rect 55033 10007 55091 10013
rect 55582 9936 55588 9988
rect 55640 9936 55646 9988
rect 55784 9948 56074 9976
rect 55784 9920 55812 9948
rect 54444 9880 54984 9908
rect 54444 9868 54450 9880
rect 55766 9868 55772 9920
rect 55824 9908 55830 9920
rect 57149 9911 57207 9917
rect 57149 9908 57161 9911
rect 55824 9880 57161 9908
rect 55824 9868 55830 9880
rect 57149 9877 57161 9880
rect 57195 9877 57207 9911
rect 57149 9871 57207 9877
rect 1104 9818 78844 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 66314 9818
rect 66366 9766 66378 9818
rect 66430 9766 66442 9818
rect 66494 9766 66506 9818
rect 66558 9766 66570 9818
rect 66622 9766 78844 9818
rect 1104 9744 78844 9766
rect 26878 9664 26884 9716
rect 26936 9704 26942 9716
rect 27341 9707 27399 9713
rect 27341 9704 27353 9707
rect 26936 9676 27353 9704
rect 26936 9664 26942 9676
rect 27341 9673 27353 9676
rect 27387 9673 27399 9707
rect 27341 9667 27399 9673
rect 31202 9664 31208 9716
rect 31260 9704 31266 9716
rect 31389 9707 31447 9713
rect 31389 9704 31401 9707
rect 31260 9676 31401 9704
rect 31260 9664 31266 9676
rect 31389 9673 31401 9676
rect 31435 9673 31447 9707
rect 31389 9667 31447 9673
rect 33980 9676 34836 9704
rect 28353 9639 28411 9645
rect 28353 9605 28365 9639
rect 28399 9636 28411 9639
rect 28442 9636 28448 9648
rect 28399 9608 28448 9636
rect 28399 9605 28411 9608
rect 28353 9599 28411 9605
rect 28442 9596 28448 9608
rect 28500 9596 28506 9648
rect 28810 9596 28816 9648
rect 28868 9596 28874 9648
rect 32398 9636 32404 9648
rect 31588 9608 32404 9636
rect 26510 9528 26516 9580
rect 26568 9568 26574 9580
rect 28077 9571 28135 9577
rect 28077 9568 28089 9571
rect 26568 9540 28089 9568
rect 26568 9528 26574 9540
rect 28077 9537 28089 9540
rect 28123 9537 28135 9571
rect 28077 9531 28135 9537
rect 27982 9460 27988 9512
rect 28040 9460 28046 9512
rect 28092 9364 28120 9531
rect 31018 9528 31024 9580
rect 31076 9568 31082 9580
rect 31588 9577 31616 9608
rect 32398 9596 32404 9608
rect 32456 9636 32462 9648
rect 33980 9636 34008 9676
rect 34698 9636 34704 9648
rect 32456 9608 34008 9636
rect 32456 9596 32462 9608
rect 31573 9571 31631 9577
rect 31573 9568 31585 9571
rect 31076 9540 31585 9568
rect 31076 9528 31082 9540
rect 31573 9537 31585 9540
rect 31619 9537 31631 9571
rect 31573 9531 31631 9537
rect 31665 9571 31723 9577
rect 31665 9537 31677 9571
rect 31711 9568 31723 9571
rect 31846 9568 31852 9580
rect 31711 9540 31852 9568
rect 31711 9537 31723 9540
rect 31665 9531 31723 9537
rect 31846 9528 31852 9540
rect 31904 9528 31910 9580
rect 33980 9577 34008 9608
rect 34072 9608 34704 9636
rect 34072 9577 34100 9608
rect 34698 9596 34704 9608
rect 34756 9596 34762 9648
rect 34808 9636 34836 9676
rect 35636 9676 35848 9704
rect 35636 9636 35664 9676
rect 34808 9608 35664 9636
rect 35710 9596 35716 9648
rect 35768 9596 35774 9648
rect 35820 9636 35848 9676
rect 40218 9664 40224 9716
rect 40276 9704 40282 9716
rect 40773 9707 40831 9713
rect 40773 9704 40785 9707
rect 40276 9676 40785 9704
rect 40276 9664 40282 9676
rect 40773 9673 40785 9676
rect 40819 9673 40831 9707
rect 45278 9704 45284 9716
rect 40773 9667 40831 9673
rect 43824 9676 45284 9704
rect 38194 9636 38200 9648
rect 35820 9608 38200 9636
rect 38194 9596 38200 9608
rect 38252 9596 38258 9648
rect 38930 9596 38936 9648
rect 38988 9596 38994 9648
rect 40034 9596 40040 9648
rect 40092 9636 40098 9648
rect 40589 9639 40647 9645
rect 40589 9636 40601 9639
rect 40092 9608 40601 9636
rect 40092 9596 40098 9608
rect 31941 9571 31999 9577
rect 31941 9537 31953 9571
rect 31987 9568 31999 9571
rect 32677 9571 32735 9577
rect 32677 9568 32689 9571
rect 31987 9540 32689 9568
rect 31987 9537 31999 9540
rect 31941 9531 31999 9537
rect 32677 9537 32689 9540
rect 32723 9537 32735 9571
rect 32677 9531 32735 9537
rect 33965 9571 34023 9577
rect 33965 9537 33977 9571
rect 34011 9537 34023 9571
rect 33965 9531 34023 9537
rect 34057 9571 34115 9577
rect 34057 9537 34069 9571
rect 34103 9537 34115 9571
rect 34057 9531 34115 9537
rect 34330 9528 34336 9580
rect 34388 9568 34394 9580
rect 34790 9568 34796 9580
rect 34388 9540 34796 9568
rect 34388 9528 34394 9540
rect 34790 9528 34796 9540
rect 34848 9528 34854 9580
rect 34977 9571 35035 9577
rect 34977 9537 34989 9571
rect 35023 9537 35035 9571
rect 34977 9531 35035 9537
rect 35161 9571 35219 9577
rect 35161 9537 35173 9571
rect 35207 9537 35219 9571
rect 35161 9531 35219 9537
rect 28810 9460 28816 9512
rect 28868 9500 28874 9512
rect 29917 9503 29975 9509
rect 29917 9500 29929 9503
rect 28868 9472 29929 9500
rect 28868 9460 28874 9472
rect 29917 9469 29929 9472
rect 29963 9500 29975 9503
rect 29963 9472 31754 9500
rect 29963 9469 29975 9472
rect 29917 9463 29975 9469
rect 31726 9444 31754 9472
rect 33042 9460 33048 9512
rect 33100 9500 33106 9512
rect 33321 9503 33379 9509
rect 33321 9500 33333 9503
rect 33100 9472 33333 9500
rect 33100 9460 33106 9472
rect 33321 9469 33333 9472
rect 33367 9500 33379 9503
rect 33410 9500 33416 9512
rect 33367 9472 33416 9500
rect 33367 9469 33379 9472
rect 33321 9463 33379 9469
rect 33410 9460 33416 9472
rect 33468 9460 33474 9512
rect 34238 9460 34244 9512
rect 34296 9460 34302 9512
rect 34606 9460 34612 9512
rect 34664 9500 34670 9512
rect 34992 9500 35020 9531
rect 34664 9472 35020 9500
rect 35176 9500 35204 9531
rect 35250 9528 35256 9580
rect 35308 9528 35314 9580
rect 35345 9571 35403 9577
rect 35345 9537 35357 9571
rect 35391 9568 35403 9571
rect 35728 9568 35756 9596
rect 35391 9540 35756 9568
rect 35391 9537 35403 9540
rect 35345 9531 35403 9537
rect 37642 9528 37648 9580
rect 37700 9528 37706 9580
rect 40512 9577 40540 9608
rect 40589 9605 40601 9608
rect 40635 9605 40647 9639
rect 40589 9599 40647 9605
rect 42705 9639 42763 9645
rect 42705 9605 42717 9639
rect 42751 9636 42763 9639
rect 42751 9608 43576 9636
rect 42751 9605 42763 9608
rect 42705 9599 42763 9605
rect 43548 9580 43576 9608
rect 40497 9571 40555 9577
rect 40497 9537 40509 9571
rect 40543 9568 40555 9571
rect 40543 9540 40577 9568
rect 40543 9537 40555 9540
rect 40497 9531 40555 9537
rect 40678 9528 40684 9580
rect 40736 9568 40742 9580
rect 40957 9571 41015 9577
rect 40957 9568 40969 9571
rect 40736 9540 40969 9568
rect 40736 9528 40742 9540
rect 40957 9537 40969 9540
rect 41003 9537 41015 9571
rect 40957 9531 41015 9537
rect 41049 9571 41107 9577
rect 41049 9537 41061 9571
rect 41095 9537 41107 9571
rect 41049 9531 41107 9537
rect 41325 9571 41383 9577
rect 41325 9537 41337 9571
rect 41371 9568 41383 9571
rect 41509 9571 41567 9577
rect 41509 9568 41521 9571
rect 41371 9540 41521 9568
rect 41371 9537 41383 9540
rect 41325 9531 41383 9537
rect 41509 9537 41521 9540
rect 41555 9537 41567 9571
rect 41509 9531 41567 9537
rect 35894 9500 35900 9512
rect 35176 9472 35900 9500
rect 34664 9460 34670 9472
rect 35894 9460 35900 9472
rect 35952 9460 35958 9512
rect 36630 9460 36636 9512
rect 36688 9500 36694 9512
rect 37274 9500 37280 9512
rect 36688 9472 37280 9500
rect 36688 9460 36694 9472
rect 37274 9460 37280 9472
rect 37332 9460 37338 9512
rect 37918 9460 37924 9512
rect 37976 9460 37982 9512
rect 40037 9503 40095 9509
rect 40037 9500 40049 9503
rect 39408 9472 40049 9500
rect 30926 9432 30932 9444
rect 29748 9404 30932 9432
rect 29748 9364 29776 9404
rect 30926 9392 30932 9404
rect 30984 9392 30990 9444
rect 31726 9404 31760 9444
rect 31754 9392 31760 9404
rect 31812 9432 31818 9444
rect 32674 9432 32680 9444
rect 31812 9404 32680 9432
rect 31812 9392 31818 9404
rect 32674 9392 32680 9404
rect 32732 9392 32738 9444
rect 33778 9392 33784 9444
rect 33836 9392 33842 9444
rect 28092 9336 29776 9364
rect 29822 9324 29828 9376
rect 29880 9324 29886 9376
rect 31849 9367 31907 9373
rect 31849 9333 31861 9367
rect 31895 9364 31907 9367
rect 33226 9364 33232 9376
rect 31895 9336 33232 9364
rect 31895 9333 31907 9336
rect 31849 9327 31907 9333
rect 33226 9324 33232 9336
rect 33284 9324 33290 9376
rect 34256 9373 34284 9460
rect 36170 9392 36176 9444
rect 36228 9432 36234 9444
rect 37458 9432 37464 9444
rect 36228 9404 37464 9432
rect 36228 9392 36234 9404
rect 37458 9392 37464 9404
rect 37516 9392 37522 9444
rect 34241 9367 34299 9373
rect 34241 9333 34253 9367
rect 34287 9333 34299 9367
rect 34241 9327 34299 9333
rect 35434 9324 35440 9376
rect 35492 9364 35498 9376
rect 35529 9367 35587 9373
rect 35529 9364 35541 9367
rect 35492 9336 35541 9364
rect 35492 9324 35498 9336
rect 35529 9333 35541 9336
rect 35575 9333 35587 9367
rect 35529 9327 35587 9333
rect 35894 9324 35900 9376
rect 35952 9324 35958 9376
rect 36262 9324 36268 9376
rect 36320 9364 36326 9376
rect 38378 9364 38384 9376
rect 36320 9336 38384 9364
rect 36320 9324 36326 9336
rect 38378 9324 38384 9336
rect 38436 9324 38442 9376
rect 39298 9324 39304 9376
rect 39356 9364 39362 9376
rect 39408 9373 39436 9472
rect 40037 9469 40049 9472
rect 40083 9469 40095 9503
rect 40037 9463 40095 9469
rect 41064 9432 41092 9531
rect 42334 9528 42340 9580
rect 42392 9568 42398 9580
rect 42613 9571 42671 9577
rect 42613 9568 42625 9571
rect 42392 9540 42625 9568
rect 42392 9528 42398 9540
rect 42613 9537 42625 9540
rect 42659 9537 42671 9571
rect 42613 9531 42671 9537
rect 42794 9528 42800 9580
rect 42852 9528 42858 9580
rect 43254 9577 43260 9580
rect 42981 9571 43039 9577
rect 42981 9537 42993 9571
rect 43027 9537 43039 9571
rect 43252 9568 43260 9577
rect 43215 9540 43260 9568
rect 42981 9531 43039 9537
rect 43252 9531 43260 9540
rect 41690 9460 41696 9512
rect 41748 9500 41754 9512
rect 42153 9503 42211 9509
rect 42153 9500 42165 9503
rect 41748 9472 42165 9500
rect 41748 9460 41754 9472
rect 42153 9469 42165 9472
rect 42199 9500 42211 9503
rect 42702 9500 42708 9512
rect 42199 9472 42708 9500
rect 42199 9469 42211 9472
rect 42153 9463 42211 9469
rect 42702 9460 42708 9472
rect 42760 9460 42766 9512
rect 42996 9500 43024 9531
rect 43254 9528 43260 9531
rect 43312 9528 43318 9580
rect 43349 9571 43407 9577
rect 43349 9537 43361 9571
rect 43395 9537 43407 9571
rect 43349 9531 43407 9537
rect 43441 9571 43499 9577
rect 43441 9537 43453 9571
rect 43487 9537 43499 9571
rect 43441 9531 43499 9537
rect 43364 9500 43392 9531
rect 42996 9472 43392 9500
rect 43456 9500 43484 9531
rect 43530 9528 43536 9580
rect 43588 9577 43594 9580
rect 43588 9571 43627 9577
rect 43615 9537 43627 9571
rect 43588 9531 43627 9537
rect 43717 9571 43775 9577
rect 43717 9537 43729 9571
rect 43763 9568 43775 9571
rect 43824 9568 43852 9676
rect 45278 9664 45284 9676
rect 45336 9664 45342 9716
rect 45554 9664 45560 9716
rect 45612 9704 45618 9716
rect 45649 9707 45707 9713
rect 45649 9704 45661 9707
rect 45612 9676 45661 9704
rect 45612 9664 45618 9676
rect 45649 9673 45661 9676
rect 45695 9673 45707 9707
rect 45649 9667 45707 9673
rect 46106 9664 46112 9716
rect 46164 9704 46170 9716
rect 49789 9707 49847 9713
rect 49789 9704 49801 9707
rect 46164 9676 49801 9704
rect 46164 9664 46170 9676
rect 49789 9673 49801 9676
rect 49835 9704 49847 9707
rect 49970 9704 49976 9716
rect 49835 9676 49976 9704
rect 49835 9673 49847 9676
rect 49789 9667 49847 9673
rect 49970 9664 49976 9676
rect 50028 9664 50034 9716
rect 50157 9707 50215 9713
rect 50157 9673 50169 9707
rect 50203 9704 50215 9707
rect 50338 9704 50344 9716
rect 50203 9676 50344 9704
rect 50203 9673 50215 9676
rect 50157 9667 50215 9673
rect 50338 9664 50344 9676
rect 50396 9664 50402 9716
rect 50706 9704 50712 9716
rect 50540 9676 50712 9704
rect 43901 9639 43959 9645
rect 43901 9605 43913 9639
rect 43947 9636 43959 9639
rect 48682 9636 48688 9648
rect 43947 9608 48688 9636
rect 43947 9605 43959 9608
rect 43901 9599 43959 9605
rect 43763 9540 43852 9568
rect 43763 9537 43775 9540
rect 43717 9531 43775 9537
rect 43588 9528 43594 9531
rect 43916 9500 43944 9599
rect 48682 9596 48688 9608
rect 48740 9596 48746 9648
rect 48961 9639 49019 9645
rect 48961 9605 48973 9639
rect 49007 9636 49019 9639
rect 49142 9636 49148 9648
rect 49007 9608 49148 9636
rect 49007 9605 49019 9608
rect 48961 9599 49019 9605
rect 49142 9596 49148 9608
rect 49200 9596 49206 9648
rect 49252 9608 49648 9636
rect 45833 9571 45891 9577
rect 45833 9537 45845 9571
rect 45879 9537 45891 9571
rect 45833 9531 45891 9537
rect 43456 9472 43944 9500
rect 45848 9500 45876 9531
rect 45922 9528 45928 9580
rect 45980 9528 45986 9580
rect 46201 9571 46259 9577
rect 46201 9537 46213 9571
rect 46247 9568 46259 9571
rect 47118 9568 47124 9580
rect 46247 9540 47124 9568
rect 46247 9537 46259 9540
rect 46201 9531 46259 9537
rect 47118 9528 47124 9540
rect 47176 9528 47182 9580
rect 49252 9577 49280 9608
rect 48869 9571 48927 9577
rect 48869 9537 48881 9571
rect 48915 9537 48927 9571
rect 48869 9531 48927 9537
rect 49053 9571 49111 9577
rect 49053 9537 49065 9571
rect 49099 9537 49111 9571
rect 49053 9531 49111 9537
rect 49237 9571 49295 9577
rect 49237 9537 49249 9571
rect 49283 9537 49295 9571
rect 49237 9531 49295 9537
rect 49329 9571 49387 9577
rect 49329 9537 49341 9571
rect 49375 9568 49387 9571
rect 49510 9568 49516 9580
rect 49375 9540 49516 9568
rect 49375 9537 49387 9540
rect 49329 9531 49387 9537
rect 47210 9500 47216 9512
rect 45848 9472 47216 9500
rect 42429 9435 42487 9441
rect 42429 9432 42441 9435
rect 41064 9404 42441 9432
rect 42429 9401 42441 9404
rect 42475 9401 42487 9435
rect 42429 9395 42487 9401
rect 39393 9367 39451 9373
rect 39393 9364 39405 9367
rect 39356 9336 39405 9364
rect 39356 9324 39362 9336
rect 39393 9333 39405 9336
rect 39439 9333 39451 9367
rect 39393 9327 39451 9333
rect 39482 9324 39488 9376
rect 39540 9324 39546 9376
rect 40310 9324 40316 9376
rect 40368 9364 40374 9376
rect 41233 9367 41291 9373
rect 41233 9364 41245 9367
rect 40368 9336 41245 9364
rect 40368 9324 40374 9336
rect 41233 9333 41245 9336
rect 41279 9333 41291 9367
rect 41233 9327 41291 9333
rect 41966 9324 41972 9376
rect 42024 9364 42030 9376
rect 42996 9364 43024 9472
rect 47210 9460 47216 9472
rect 47268 9460 47274 9512
rect 48884 9432 48912 9531
rect 49068 9500 49096 9531
rect 49510 9528 49516 9540
rect 49568 9528 49574 9580
rect 49620 9568 49648 9608
rect 49694 9596 49700 9648
rect 49752 9636 49758 9648
rect 50246 9636 50252 9648
rect 49752 9608 50252 9636
rect 49752 9596 49758 9608
rect 50246 9596 50252 9608
rect 50304 9636 50310 9648
rect 50540 9645 50568 9676
rect 50706 9664 50712 9676
rect 50764 9664 50770 9716
rect 51166 9704 51172 9716
rect 51092 9676 51172 9704
rect 51092 9645 51120 9676
rect 51166 9664 51172 9676
rect 51224 9664 51230 9716
rect 51353 9707 51411 9713
rect 51353 9673 51365 9707
rect 51399 9704 51411 9707
rect 51718 9704 51724 9716
rect 51399 9676 51724 9704
rect 51399 9673 51411 9676
rect 51353 9667 51411 9673
rect 51718 9664 51724 9676
rect 51776 9664 51782 9716
rect 51905 9707 51963 9713
rect 51905 9673 51917 9707
rect 51951 9704 51963 9707
rect 51994 9704 52000 9716
rect 51951 9676 52000 9704
rect 51951 9673 51963 9676
rect 51905 9667 51963 9673
rect 51994 9664 52000 9676
rect 52052 9664 52058 9716
rect 52825 9707 52883 9713
rect 52825 9673 52837 9707
rect 52871 9704 52883 9707
rect 52914 9704 52920 9716
rect 52871 9676 52920 9704
rect 52871 9673 52883 9676
rect 52825 9667 52883 9673
rect 52914 9664 52920 9676
rect 52972 9664 52978 9716
rect 54938 9664 54944 9716
rect 54996 9704 55002 9716
rect 54996 9676 55168 9704
rect 54996 9664 55002 9676
rect 55140 9674 55168 9676
rect 55490 9674 55496 9686
rect 50433 9639 50491 9645
rect 50433 9636 50445 9639
rect 50304 9608 50445 9636
rect 50304 9596 50310 9608
rect 50433 9605 50445 9608
rect 50479 9605 50491 9639
rect 50433 9599 50491 9605
rect 50525 9639 50583 9645
rect 50525 9605 50537 9639
rect 50571 9605 50583 9639
rect 50985 9639 51043 9645
rect 50985 9636 50997 9639
rect 50525 9599 50583 9605
rect 50632 9608 50997 9636
rect 49620 9540 50292 9568
rect 50062 9500 50068 9512
rect 49068 9472 50068 9500
rect 50062 9460 50068 9472
rect 50120 9460 50126 9512
rect 50264 9500 50292 9540
rect 50338 9528 50344 9580
rect 50396 9528 50402 9580
rect 50430 9500 50436 9512
rect 50264 9472 50436 9500
rect 50430 9460 50436 9472
rect 50488 9460 50494 9512
rect 49513 9435 49571 9441
rect 49513 9432 49525 9435
rect 48884 9404 49525 9432
rect 49513 9401 49525 9404
rect 49559 9432 49571 9435
rect 49970 9432 49976 9444
rect 49559 9404 49976 9432
rect 49559 9401 49571 9404
rect 49513 9395 49571 9401
rect 49970 9392 49976 9404
rect 50028 9432 50034 9444
rect 50028 9404 50292 9432
rect 50028 9392 50034 9404
rect 42024 9336 43024 9364
rect 43073 9367 43131 9373
rect 42024 9324 42030 9336
rect 43073 9333 43085 9367
rect 43119 9364 43131 9367
rect 43714 9364 43720 9376
rect 43119 9336 43720 9364
rect 43119 9333 43131 9336
rect 43073 9327 43131 9333
rect 43714 9324 43720 9336
rect 43772 9324 43778 9376
rect 46109 9367 46167 9373
rect 46109 9333 46121 9367
rect 46155 9364 46167 9367
rect 46842 9364 46848 9376
rect 46155 9336 46848 9364
rect 46155 9333 46167 9336
rect 46109 9327 46167 9333
rect 46842 9324 46848 9336
rect 46900 9324 46906 9376
rect 48685 9367 48743 9373
rect 48685 9333 48697 9367
rect 48731 9364 48743 9367
rect 48866 9364 48872 9376
rect 48731 9336 48872 9364
rect 48731 9333 48743 9336
rect 48685 9327 48743 9333
rect 48866 9324 48872 9336
rect 48924 9324 48930 9376
rect 49881 9367 49939 9373
rect 49881 9333 49893 9367
rect 49927 9364 49939 9367
rect 50154 9364 50160 9376
rect 49927 9336 50160 9364
rect 49927 9333 49939 9336
rect 49881 9327 49939 9333
rect 50154 9324 50160 9336
rect 50212 9324 50218 9376
rect 50264 9364 50292 9404
rect 50338 9392 50344 9444
rect 50396 9432 50402 9444
rect 50632 9432 50660 9608
rect 50985 9605 50997 9608
rect 51031 9605 51043 9639
rect 50985 9599 51043 9605
rect 51077 9639 51135 9645
rect 51077 9605 51089 9639
rect 51123 9605 51135 9639
rect 51626 9636 51632 9648
rect 51077 9599 51135 9605
rect 51184 9608 51632 9636
rect 50709 9571 50767 9577
rect 50709 9537 50721 9571
rect 50755 9537 50767 9571
rect 50709 9531 50767 9537
rect 50801 9571 50859 9577
rect 50801 9537 50813 9571
rect 50847 9568 50859 9571
rect 50890 9568 50896 9580
rect 50847 9540 50896 9568
rect 50847 9537 50859 9540
rect 50801 9531 50859 9537
rect 50396 9404 50660 9432
rect 50724 9500 50752 9531
rect 50890 9528 50896 9540
rect 50948 9528 50954 9580
rect 51184 9577 51212 9608
rect 51626 9596 51632 9608
rect 51684 9596 51690 9648
rect 55140 9646 55496 9674
rect 55490 9634 55496 9646
rect 55548 9634 55554 9686
rect 55582 9664 55588 9716
rect 55640 9704 55646 9716
rect 55677 9707 55735 9713
rect 55677 9704 55689 9707
rect 55640 9676 55689 9704
rect 55640 9664 55646 9676
rect 55677 9673 55689 9676
rect 55723 9673 55735 9707
rect 55677 9667 55735 9673
rect 51169 9571 51227 9577
rect 51169 9537 51181 9571
rect 51215 9537 51227 9571
rect 51169 9531 51227 9537
rect 51350 9528 51356 9580
rect 51408 9568 51414 9580
rect 51445 9571 51503 9577
rect 51445 9568 51457 9571
rect 51408 9540 51457 9568
rect 51408 9528 51414 9540
rect 51445 9537 51457 9540
rect 51491 9537 51503 9571
rect 51445 9531 51503 9537
rect 53006 9528 53012 9580
rect 53064 9528 53070 9580
rect 53285 9571 53343 9577
rect 53285 9537 53297 9571
rect 53331 9568 53343 9571
rect 54202 9568 54208 9580
rect 53331 9540 54208 9568
rect 53331 9537 53343 9540
rect 53285 9531 53343 9537
rect 54202 9528 54208 9540
rect 54260 9528 54266 9580
rect 54478 9528 54484 9580
rect 54536 9528 54542 9580
rect 54662 9528 54668 9580
rect 54720 9528 54726 9580
rect 54757 9571 54815 9577
rect 54757 9537 54769 9571
rect 54803 9537 54815 9571
rect 54757 9531 54815 9537
rect 54849 9571 54907 9577
rect 54849 9537 54861 9571
rect 54895 9568 54907 9571
rect 54938 9568 54944 9580
rect 54895 9540 54944 9568
rect 54895 9537 54907 9540
rect 54849 9531 54907 9537
rect 54386 9500 54392 9512
rect 50724 9472 54392 9500
rect 50724 9432 50752 9472
rect 54386 9460 54392 9472
rect 54444 9500 54450 9512
rect 54772 9500 54800 9531
rect 54938 9528 54944 9540
rect 54996 9528 55002 9580
rect 55171 9571 55229 9577
rect 55171 9537 55183 9571
rect 55217 9537 55229 9571
rect 55171 9531 55229 9537
rect 54444 9472 54800 9500
rect 55186 9500 55214 9531
rect 55306 9528 55312 9580
rect 55364 9568 55370 9580
rect 55401 9571 55459 9577
rect 55401 9568 55413 9571
rect 55364 9540 55413 9568
rect 55364 9528 55370 9540
rect 55401 9537 55413 9540
rect 55447 9537 55459 9571
rect 55401 9531 55459 9537
rect 55490 9528 55496 9580
rect 55548 9528 55554 9580
rect 56594 9528 56600 9580
rect 56652 9528 56658 9580
rect 55186 9472 56088 9500
rect 54444 9460 54450 9472
rect 50798 9432 50804 9444
rect 50724 9404 50804 9432
rect 50396 9392 50402 9404
rect 50798 9392 50804 9404
rect 50856 9392 50862 9444
rect 51166 9392 51172 9444
rect 51224 9432 51230 9444
rect 51442 9432 51448 9444
rect 51224 9404 51448 9432
rect 51224 9392 51230 9404
rect 51442 9392 51448 9404
rect 51500 9392 51506 9444
rect 52362 9432 52368 9444
rect 51736 9404 52368 9432
rect 51736 9364 51764 9404
rect 52362 9392 52368 9404
rect 52420 9392 52426 9444
rect 56060 9441 56088 9472
rect 56045 9435 56103 9441
rect 56045 9401 56057 9435
rect 56091 9401 56103 9435
rect 56045 9395 56103 9401
rect 50264 9336 51764 9364
rect 51902 9324 51908 9376
rect 51960 9364 51966 9376
rect 53190 9364 53196 9376
rect 51960 9336 53196 9364
rect 51960 9324 51966 9336
rect 53190 9324 53196 9336
rect 53248 9324 53254 9376
rect 55030 9324 55036 9376
rect 55088 9324 55094 9376
rect 55217 9367 55275 9373
rect 55217 9333 55229 9367
rect 55263 9364 55275 9367
rect 55490 9364 55496 9376
rect 55263 9336 55496 9364
rect 55263 9333 55275 9336
rect 55217 9327 55275 9333
rect 55490 9324 55496 9336
rect 55548 9324 55554 9376
rect 1104 9274 78844 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 78844 9274
rect 1104 9200 78844 9222
rect 28258 9120 28264 9172
rect 28316 9120 28322 9172
rect 31294 9120 31300 9172
rect 31352 9160 31358 9172
rect 31478 9160 31484 9172
rect 31352 9132 31484 9160
rect 31352 9120 31358 9132
rect 31478 9120 31484 9132
rect 31536 9120 31542 9172
rect 31846 9120 31852 9172
rect 31904 9120 31910 9172
rect 34517 9163 34575 9169
rect 34517 9160 34529 9163
rect 32876 9132 34529 9160
rect 32876 9092 32904 9132
rect 34517 9129 34529 9132
rect 34563 9129 34575 9163
rect 34517 9123 34575 9129
rect 31404 9064 32904 9092
rect 26510 8984 26516 9036
rect 26568 8984 26574 9036
rect 26789 9027 26847 9033
rect 26789 8993 26801 9027
rect 26835 9024 26847 9027
rect 27154 9024 27160 9036
rect 26835 8996 27160 9024
rect 26835 8993 26847 8996
rect 26789 8987 26847 8993
rect 27154 8984 27160 8996
rect 27212 8984 27218 9036
rect 30745 8959 30803 8965
rect 30745 8925 30757 8959
rect 30791 8956 30803 8959
rect 31113 8959 31171 8965
rect 31113 8956 31125 8959
rect 30791 8928 31125 8956
rect 30791 8925 30803 8928
rect 30745 8919 30803 8925
rect 31113 8925 31125 8928
rect 31159 8925 31171 8959
rect 31113 8919 31171 8925
rect 31128 8888 31156 8919
rect 31202 8916 31208 8968
rect 31260 8956 31266 8968
rect 31297 8959 31355 8965
rect 31297 8956 31309 8959
rect 31260 8928 31309 8956
rect 31260 8916 31266 8928
rect 31297 8925 31309 8928
rect 31343 8956 31355 8959
rect 31404 8956 31432 9064
rect 32769 9027 32827 9033
rect 32769 8993 32781 9027
rect 32815 9024 32827 9027
rect 33594 9024 33600 9036
rect 32815 8996 33600 9024
rect 32815 8993 32827 8996
rect 32769 8987 32827 8993
rect 33594 8984 33600 8996
rect 33652 8984 33658 9036
rect 34532 9024 34560 9123
rect 37918 9120 37924 9172
rect 37976 9160 37982 9172
rect 38197 9163 38255 9169
rect 38197 9160 38209 9163
rect 37976 9132 38209 9160
rect 37976 9120 37982 9132
rect 38197 9129 38209 9132
rect 38243 9129 38255 9163
rect 38197 9123 38255 9129
rect 38378 9120 38384 9172
rect 38436 9160 38442 9172
rect 42610 9160 42616 9172
rect 38436 9132 42616 9160
rect 38436 9120 38442 9132
rect 42610 9120 42616 9132
rect 42668 9120 42674 9172
rect 42886 9120 42892 9172
rect 42944 9160 42950 9172
rect 43254 9160 43260 9172
rect 42944 9132 43260 9160
rect 42944 9120 42950 9132
rect 43254 9120 43260 9132
rect 43312 9120 43318 9172
rect 49237 9163 49295 9169
rect 49237 9129 49249 9163
rect 49283 9160 49295 9163
rect 49510 9160 49516 9172
rect 49283 9132 49516 9160
rect 49283 9129 49295 9132
rect 49237 9123 49295 9129
rect 49510 9120 49516 9132
rect 49568 9120 49574 9172
rect 49694 9120 49700 9172
rect 49752 9120 49758 9172
rect 49878 9120 49884 9172
rect 49936 9160 49942 9172
rect 50617 9163 50675 9169
rect 50617 9160 50629 9163
rect 49936 9132 50629 9160
rect 49936 9120 49942 9132
rect 50617 9129 50629 9132
rect 50663 9129 50675 9163
rect 50617 9123 50675 9129
rect 50890 9120 50896 9172
rect 50948 9160 50954 9172
rect 51261 9163 51319 9169
rect 51261 9160 51273 9163
rect 50948 9132 51273 9160
rect 50948 9120 50954 9132
rect 51261 9129 51273 9132
rect 51307 9129 51319 9163
rect 51261 9123 51319 9129
rect 55030 9120 55036 9172
rect 55088 9160 55094 9172
rect 55306 9160 55312 9172
rect 55088 9132 55312 9160
rect 55088 9120 55094 9132
rect 55306 9120 55312 9132
rect 55364 9120 55370 9172
rect 35986 9052 35992 9104
rect 36044 9052 36050 9104
rect 36998 9092 37004 9104
rect 36280 9064 37004 9092
rect 35158 9024 35164 9036
rect 34532 8996 35164 9024
rect 35158 8984 35164 8996
rect 35216 9024 35222 9036
rect 35253 9027 35311 9033
rect 35253 9024 35265 9027
rect 35216 8996 35265 9024
rect 35216 8984 35222 8996
rect 35253 8993 35265 8996
rect 35299 8993 35311 9027
rect 35253 8987 35311 8993
rect 31343 8928 31432 8956
rect 31343 8925 31355 8928
rect 31297 8919 31355 8925
rect 31478 8916 31484 8968
rect 31536 8916 31542 8968
rect 31662 8916 31668 8968
rect 31720 8916 31726 8968
rect 32214 8965 32220 8968
rect 32033 8959 32091 8965
rect 32033 8925 32045 8959
rect 32079 8925 32091 8959
rect 32033 8919 32091 8925
rect 32181 8959 32220 8965
rect 32181 8925 32193 8959
rect 32181 8919 32220 8925
rect 31386 8888 31392 8900
rect 22066 8860 27278 8888
rect 31128 8860 31392 8888
rect 22066 8832 22094 8860
rect 22002 8780 22008 8832
rect 22060 8792 22094 8832
rect 27172 8820 27200 8860
rect 31386 8848 31392 8860
rect 31444 8848 31450 8900
rect 31570 8848 31576 8900
rect 31628 8848 31634 8900
rect 28353 8823 28411 8829
rect 28353 8820 28365 8823
rect 27172 8792 28365 8820
rect 22060 8780 22066 8792
rect 28353 8789 28365 8792
rect 28399 8820 28411 8823
rect 28810 8820 28816 8832
rect 28399 8792 28816 8820
rect 28399 8789 28411 8792
rect 28353 8783 28411 8789
rect 28810 8780 28816 8792
rect 28868 8780 28874 8832
rect 30929 8823 30987 8829
rect 30929 8789 30941 8823
rect 30975 8820 30987 8823
rect 31478 8820 31484 8832
rect 30975 8792 31484 8820
rect 30975 8789 30987 8792
rect 30929 8783 30987 8789
rect 31478 8780 31484 8792
rect 31536 8780 31542 8832
rect 32048 8820 32076 8919
rect 32214 8916 32220 8919
rect 32272 8916 32278 8968
rect 32398 8916 32404 8968
rect 32456 8916 32462 8968
rect 32537 8959 32595 8965
rect 32537 8925 32549 8959
rect 32583 8956 32595 8959
rect 32583 8928 32812 8956
rect 32583 8925 32595 8928
rect 32537 8919 32595 8925
rect 32784 8900 32812 8928
rect 35894 8916 35900 8968
rect 35952 8916 35958 8968
rect 36004 8965 36032 9052
rect 36280 8965 36308 9064
rect 36998 9052 37004 9064
rect 37056 9052 37062 9104
rect 37274 9052 37280 9104
rect 37332 9052 37338 9104
rect 38562 9052 38568 9104
rect 38620 9092 38626 9104
rect 38657 9095 38715 9101
rect 38657 9092 38669 9095
rect 38620 9064 38669 9092
rect 38620 9052 38626 9064
rect 38657 9061 38669 9064
rect 38703 9092 38715 9095
rect 40310 9092 40316 9104
rect 38703 9064 40316 9092
rect 38703 9061 38715 9064
rect 38657 9055 38715 9061
rect 40310 9052 40316 9064
rect 40368 9052 40374 9104
rect 43625 9095 43683 9101
rect 43625 9092 43637 9095
rect 40420 9064 43637 9092
rect 36814 8984 36820 9036
rect 36872 8984 36878 9036
rect 37369 9027 37427 9033
rect 37369 8993 37381 9027
rect 37415 8993 37427 9027
rect 37369 8987 37427 8993
rect 35990 8959 36048 8965
rect 35990 8925 36002 8959
rect 36036 8925 36048 8959
rect 35990 8919 36048 8925
rect 36265 8959 36323 8965
rect 36265 8925 36277 8959
rect 36311 8925 36323 8959
rect 36265 8919 36323 8925
rect 36354 8916 36360 8968
rect 36412 8965 36418 8968
rect 36412 8956 36420 8965
rect 36412 8928 36457 8956
rect 36412 8919 36420 8928
rect 36412 8916 36418 8919
rect 36630 8916 36636 8968
rect 36688 8916 36694 8968
rect 36726 8959 36784 8965
rect 36726 8925 36738 8959
rect 36772 8925 36784 8959
rect 36832 8956 36860 8984
rect 37098 8959 37156 8965
rect 37098 8956 37110 8959
rect 36832 8928 37110 8956
rect 36726 8919 36784 8925
rect 37098 8925 37110 8928
rect 37144 8956 37156 8959
rect 37384 8956 37412 8987
rect 37458 8984 37464 9036
rect 37516 9024 37522 9036
rect 38010 9024 38016 9036
rect 37516 8996 38016 9024
rect 37516 8984 37522 8996
rect 38010 8984 38016 8996
rect 38068 9024 38074 9036
rect 40420 9024 40448 9064
rect 43625 9061 43637 9064
rect 43671 9061 43683 9095
rect 43625 9055 43683 9061
rect 38068 8996 40448 9024
rect 38068 8984 38074 8996
rect 42610 8984 42616 9036
rect 42668 9024 42674 9036
rect 43441 9027 43499 9033
rect 43441 9024 43453 9027
rect 42668 8996 43453 9024
rect 42668 8984 42674 8996
rect 43441 8993 43453 8996
rect 43487 8993 43499 9027
rect 43441 8987 43499 8993
rect 37144 8928 37412 8956
rect 37553 8959 37611 8965
rect 37144 8925 37156 8928
rect 37098 8919 37156 8925
rect 37553 8925 37565 8959
rect 37599 8956 37611 8959
rect 38286 8956 38292 8968
rect 37599 8928 38292 8956
rect 37599 8925 37611 8928
rect 37553 8919 37611 8925
rect 32309 8891 32367 8897
rect 32309 8857 32321 8891
rect 32355 8857 32367 8891
rect 32309 8851 32367 8857
rect 32214 8820 32220 8832
rect 32048 8792 32220 8820
rect 32214 8780 32220 8792
rect 32272 8780 32278 8832
rect 32324 8820 32352 8851
rect 32766 8848 32772 8900
rect 32824 8848 32830 8900
rect 33042 8848 33048 8900
rect 33100 8848 33106 8900
rect 34422 8888 34428 8900
rect 34270 8860 34428 8888
rect 32582 8820 32588 8832
rect 32324 8792 32588 8820
rect 32582 8780 32588 8792
rect 32640 8780 32646 8832
rect 32674 8780 32680 8832
rect 32732 8780 32738 8832
rect 33962 8780 33968 8832
rect 34020 8820 34026 8832
rect 34348 8820 34376 8860
rect 34422 8848 34428 8860
rect 34480 8848 34486 8900
rect 36170 8848 36176 8900
rect 36228 8848 36234 8900
rect 34020 8792 34376 8820
rect 34020 8780 34026 8792
rect 34698 8780 34704 8832
rect 34756 8780 34762 8832
rect 36538 8780 36544 8832
rect 36596 8780 36602 8832
rect 36630 8780 36636 8832
rect 36688 8820 36694 8832
rect 36740 8820 36768 8919
rect 36909 8891 36967 8897
rect 36909 8857 36921 8891
rect 36955 8857 36967 8891
rect 36909 8851 36967 8857
rect 37001 8891 37059 8897
rect 37001 8857 37013 8891
rect 37047 8888 37059 8891
rect 37642 8888 37648 8900
rect 37047 8860 37648 8888
rect 37047 8857 37059 8860
rect 37001 8851 37059 8857
rect 36688 8792 36768 8820
rect 36924 8820 36952 8851
rect 37642 8848 37648 8860
rect 37700 8848 37706 8900
rect 37752 8820 37780 8928
rect 38286 8916 38292 8928
rect 38344 8916 38350 8968
rect 38378 8916 38384 8968
rect 38436 8916 38442 8968
rect 38470 8916 38476 8968
rect 38528 8916 38534 8968
rect 38749 8959 38807 8965
rect 38749 8925 38761 8959
rect 38795 8956 38807 8959
rect 39482 8956 39488 8968
rect 38795 8928 39488 8956
rect 38795 8925 38807 8928
rect 38749 8919 38807 8925
rect 39482 8916 39488 8928
rect 39540 8916 39546 8968
rect 41966 8916 41972 8968
rect 42024 8916 42030 8968
rect 42058 8916 42064 8968
rect 42116 8916 42122 8968
rect 38304 8888 38332 8916
rect 41690 8888 41696 8900
rect 38304 8860 41696 8888
rect 41690 8848 41696 8860
rect 41748 8848 41754 8900
rect 43456 8888 43484 8987
rect 43640 8956 43668 9055
rect 46290 9052 46296 9104
rect 46348 9092 46354 9104
rect 50338 9092 50344 9104
rect 46348 9064 50344 9092
rect 46348 9052 46354 9064
rect 50338 9052 50344 9064
rect 50396 9092 50402 9104
rect 50433 9095 50491 9101
rect 50433 9092 50445 9095
rect 50396 9064 50445 9092
rect 50396 9052 50402 9064
rect 50433 9061 50445 9064
rect 50479 9061 50491 9095
rect 50433 9055 50491 9061
rect 50706 9052 50712 9104
rect 50764 9052 50770 9104
rect 51074 9052 51080 9104
rect 51132 9092 51138 9104
rect 51132 9064 51580 9092
rect 51132 9052 51138 9064
rect 44174 8984 44180 9036
rect 44232 9024 44238 9036
rect 49602 9024 49608 9036
rect 44232 8996 49608 9024
rect 44232 8984 44238 8996
rect 49602 8984 49608 8996
rect 49660 8984 49666 9036
rect 49694 8984 49700 9036
rect 49752 9024 49758 9036
rect 49789 9027 49847 9033
rect 49789 9024 49801 9027
rect 49752 8996 49801 9024
rect 49752 8984 49758 8996
rect 49789 8993 49801 8996
rect 49835 9024 49847 9027
rect 50724 9024 50752 9052
rect 49835 8996 50752 9024
rect 49835 8993 49847 8996
rect 49789 8987 49847 8993
rect 50982 8984 50988 9036
rect 51040 9024 51046 9036
rect 51353 9027 51411 9033
rect 51353 9024 51365 9027
rect 51040 8996 51365 9024
rect 51040 8984 51046 8996
rect 51353 8993 51365 8996
rect 51399 8993 51411 9027
rect 51353 8987 51411 8993
rect 43947 8959 44005 8965
rect 43947 8956 43959 8959
rect 43640 8928 43959 8956
rect 43947 8925 43959 8928
rect 43993 8925 44005 8959
rect 43947 8919 44005 8925
rect 44082 8916 44088 8968
rect 44140 8916 44146 8968
rect 44358 8916 44364 8968
rect 44416 8916 44422 8968
rect 44450 8916 44456 8968
rect 44508 8916 44514 8968
rect 45462 8916 45468 8968
rect 45520 8956 45526 8968
rect 49050 8956 49056 8968
rect 45520 8928 49056 8956
rect 45520 8916 45526 8928
rect 49050 8916 49056 8928
rect 49108 8956 49114 8968
rect 50801 8959 50859 8965
rect 50801 8956 50813 8959
rect 49108 8928 50813 8956
rect 49108 8916 49114 8928
rect 50801 8925 50813 8928
rect 50847 8956 50859 8959
rect 51074 8956 51080 8968
rect 50847 8928 51080 8956
rect 50847 8925 50859 8928
rect 50801 8919 50859 8925
rect 51074 8916 51080 8928
rect 51132 8916 51138 8968
rect 51169 8959 51227 8965
rect 51169 8925 51181 8959
rect 51215 8925 51227 8959
rect 51169 8919 51227 8925
rect 44177 8891 44235 8897
rect 44177 8888 44189 8891
rect 43456 8860 44189 8888
rect 44177 8857 44189 8860
rect 44223 8857 44235 8891
rect 44177 8851 44235 8857
rect 44910 8848 44916 8900
rect 44968 8888 44974 8900
rect 45373 8891 45431 8897
rect 45373 8888 45385 8891
rect 44968 8860 45385 8888
rect 44968 8848 44974 8860
rect 45373 8857 45385 8860
rect 45419 8888 45431 8891
rect 49694 8888 49700 8900
rect 45419 8860 49700 8888
rect 45419 8857 45431 8860
rect 45373 8851 45431 8857
rect 49694 8848 49700 8860
rect 49752 8848 49758 8900
rect 50338 8848 50344 8900
rect 50396 8888 50402 8900
rect 50893 8891 50951 8897
rect 50893 8888 50905 8891
rect 50396 8860 50905 8888
rect 50396 8848 50402 8860
rect 50893 8857 50905 8860
rect 50939 8857 50951 8891
rect 50893 8851 50951 8857
rect 50982 8848 50988 8900
rect 51040 8848 51046 8900
rect 51184 8888 51212 8919
rect 51258 8916 51264 8968
rect 51316 8916 51322 8968
rect 51552 8965 51580 9064
rect 51537 8959 51595 8965
rect 51537 8925 51549 8959
rect 51583 8925 51595 8959
rect 51537 8919 51595 8925
rect 51626 8888 51632 8900
rect 51184 8860 51632 8888
rect 51626 8848 51632 8860
rect 51684 8848 51690 8900
rect 36924 8792 37780 8820
rect 36688 8780 36694 8792
rect 38378 8780 38384 8832
rect 38436 8820 38442 8832
rect 38838 8820 38844 8832
rect 38436 8792 38844 8820
rect 38436 8780 38442 8792
rect 38838 8780 38844 8792
rect 38896 8820 38902 8832
rect 40678 8820 40684 8832
rect 38896 8792 40684 8820
rect 38896 8780 38902 8792
rect 40678 8780 40684 8792
rect 40736 8780 40742 8832
rect 40862 8780 40868 8832
rect 40920 8820 40926 8832
rect 41325 8823 41383 8829
rect 41325 8820 41337 8823
rect 40920 8792 41337 8820
rect 40920 8780 40926 8792
rect 41325 8789 41337 8792
rect 41371 8789 41383 8823
rect 41325 8783 41383 8789
rect 41782 8780 41788 8832
rect 41840 8820 41846 8832
rect 42245 8823 42303 8829
rect 42245 8820 42257 8823
rect 41840 8792 42257 8820
rect 41840 8780 41846 8792
rect 42245 8789 42257 8792
rect 42291 8820 42303 8823
rect 42334 8820 42340 8832
rect 42291 8792 42340 8820
rect 42291 8789 42303 8792
rect 42245 8783 42303 8789
rect 42334 8780 42340 8792
rect 42392 8780 42398 8832
rect 43806 8780 43812 8832
rect 43864 8780 43870 8832
rect 46842 8780 46848 8832
rect 46900 8820 46906 8832
rect 48958 8820 48964 8832
rect 46900 8792 48964 8820
rect 46900 8780 46906 8792
rect 48958 8780 48964 8792
rect 49016 8780 49022 8832
rect 50154 8780 50160 8832
rect 50212 8780 50218 8832
rect 51350 8780 51356 8832
rect 51408 8820 51414 8832
rect 51721 8823 51779 8829
rect 51721 8820 51733 8823
rect 51408 8792 51733 8820
rect 51408 8780 51414 8792
rect 51721 8789 51733 8792
rect 51767 8789 51779 8823
rect 51721 8783 51779 8789
rect 1104 8730 78844 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 66314 8730
rect 66366 8678 66378 8730
rect 66430 8678 66442 8730
rect 66494 8678 66506 8730
rect 66558 8678 66570 8730
rect 66622 8678 78844 8730
rect 1104 8656 78844 8678
rect 31573 8619 31631 8625
rect 31573 8616 31585 8619
rect 31128 8588 31585 8616
rect 29454 8548 29460 8560
rect 28920 8520 29460 8548
rect 28920 8489 28948 8520
rect 29454 8508 29460 8520
rect 29512 8508 29518 8560
rect 31128 8548 31156 8588
rect 31573 8585 31585 8588
rect 31619 8616 31631 8619
rect 31754 8616 31760 8628
rect 31619 8588 31760 8616
rect 31619 8585 31631 8588
rect 31573 8579 31631 8585
rect 31754 8576 31760 8588
rect 31812 8576 31818 8628
rect 32861 8619 32919 8625
rect 32861 8585 32873 8619
rect 32907 8616 32919 8619
rect 33042 8616 33048 8628
rect 32907 8588 33048 8616
rect 32907 8585 32919 8588
rect 32861 8579 32919 8585
rect 33042 8576 33048 8588
rect 33100 8576 33106 8628
rect 35342 8576 35348 8628
rect 35400 8576 35406 8628
rect 35434 8576 35440 8628
rect 35492 8576 35498 8628
rect 35526 8576 35532 8628
rect 35584 8616 35590 8628
rect 36449 8619 36507 8625
rect 35584 8588 35940 8616
rect 35584 8576 35590 8588
rect 30406 8520 31156 8548
rect 31205 8551 31263 8557
rect 31205 8517 31217 8551
rect 31251 8548 31263 8551
rect 31294 8548 31300 8560
rect 31251 8520 31300 8548
rect 31251 8517 31263 8520
rect 31205 8511 31263 8517
rect 31294 8508 31300 8520
rect 31352 8548 31358 8560
rect 32122 8548 32128 8560
rect 31352 8520 32128 8548
rect 31352 8508 31358 8520
rect 32122 8508 32128 8520
rect 32180 8548 32186 8560
rect 32582 8548 32588 8560
rect 32180 8520 32588 8548
rect 32180 8508 32186 8520
rect 32582 8508 32588 8520
rect 32640 8508 32646 8560
rect 32766 8508 32772 8560
rect 32824 8548 32830 8560
rect 35360 8548 35388 8576
rect 32824 8520 35388 8548
rect 35452 8548 35480 8576
rect 35452 8520 35848 8548
rect 32824 8508 32830 8520
rect 31018 8489 31024 8492
rect 28905 8483 28963 8489
rect 28905 8449 28917 8483
rect 28951 8449 28963 8483
rect 31016 8480 31024 8489
rect 30979 8452 31024 8480
rect 28905 8443 28963 8449
rect 31016 8443 31024 8452
rect 31018 8440 31024 8443
rect 31076 8440 31082 8492
rect 31110 8440 31116 8492
rect 31168 8440 31174 8492
rect 31386 8440 31392 8492
rect 31444 8440 31450 8492
rect 31478 8440 31484 8492
rect 31536 8440 31542 8492
rect 32674 8440 32680 8492
rect 32732 8480 32738 8492
rect 33045 8483 33103 8489
rect 33045 8480 33057 8483
rect 32732 8452 33057 8480
rect 32732 8440 32738 8452
rect 33045 8449 33057 8452
rect 33091 8449 33103 8483
rect 33045 8443 33103 8449
rect 33321 8483 33379 8489
rect 33321 8449 33333 8483
rect 33367 8480 33379 8483
rect 34698 8480 34704 8492
rect 33367 8452 34704 8480
rect 33367 8449 33379 8452
rect 33321 8443 33379 8449
rect 34698 8440 34704 8452
rect 34756 8440 34762 8492
rect 35069 8483 35127 8489
rect 35069 8449 35081 8483
rect 35115 8449 35127 8483
rect 35069 8443 35127 8449
rect 29178 8372 29184 8424
rect 29236 8372 29242 8424
rect 31496 8412 31524 8440
rect 32214 8412 32220 8424
rect 31496 8384 32220 8412
rect 32214 8372 32220 8384
rect 32272 8412 32278 8424
rect 32950 8412 32956 8424
rect 32272 8384 32956 8412
rect 32272 8372 32278 8384
rect 32950 8372 32956 8384
rect 33008 8372 33014 8424
rect 33226 8372 33232 8424
rect 33284 8412 33290 8424
rect 33686 8412 33692 8424
rect 33284 8384 33692 8412
rect 33284 8372 33290 8384
rect 33686 8372 33692 8384
rect 33744 8412 33750 8424
rect 33870 8412 33876 8424
rect 33744 8384 33876 8412
rect 33744 8372 33750 8384
rect 33870 8372 33876 8384
rect 33928 8372 33934 8424
rect 30653 8347 30711 8353
rect 30653 8313 30665 8347
rect 30699 8344 30711 8347
rect 31110 8344 31116 8356
rect 30699 8316 31116 8344
rect 30699 8313 30711 8316
rect 30653 8307 30711 8313
rect 31110 8304 31116 8316
rect 31168 8304 31174 8356
rect 31386 8304 31392 8356
rect 31444 8344 31450 8356
rect 32766 8344 32772 8356
rect 31444 8316 32772 8344
rect 31444 8304 31450 8316
rect 32766 8304 32772 8316
rect 32824 8304 32830 8356
rect 35084 8344 35112 8443
rect 35158 8440 35164 8492
rect 35216 8480 35222 8492
rect 35345 8483 35403 8489
rect 35216 8452 35261 8480
rect 35216 8440 35222 8452
rect 35345 8449 35357 8483
rect 35391 8449 35403 8483
rect 35345 8443 35403 8449
rect 35360 8412 35388 8443
rect 35434 8440 35440 8492
rect 35492 8440 35498 8492
rect 35575 8483 35633 8489
rect 35575 8449 35587 8483
rect 35621 8480 35633 8483
rect 35710 8480 35716 8492
rect 35621 8452 35716 8480
rect 35621 8449 35633 8452
rect 35575 8443 35633 8449
rect 35710 8440 35716 8452
rect 35768 8440 35774 8492
rect 35820 8489 35848 8520
rect 35912 8489 35940 8588
rect 36449 8585 36461 8619
rect 36495 8585 36507 8619
rect 36449 8579 36507 8585
rect 35805 8483 35863 8489
rect 35805 8449 35817 8483
rect 35851 8449 35863 8483
rect 35805 8443 35863 8449
rect 35898 8483 35956 8489
rect 35898 8449 35910 8483
rect 35944 8449 35956 8483
rect 35898 8443 35956 8449
rect 36081 8483 36139 8489
rect 36081 8449 36093 8483
rect 36127 8449 36139 8483
rect 36081 8443 36139 8449
rect 36096 8412 36124 8443
rect 36170 8440 36176 8492
rect 36228 8440 36234 8492
rect 36262 8440 36268 8492
rect 36320 8489 36326 8492
rect 36320 8480 36328 8489
rect 36464 8480 36492 8579
rect 36538 8576 36544 8628
rect 36596 8616 36602 8628
rect 37550 8616 37556 8628
rect 36596 8588 37556 8616
rect 36596 8576 36602 8588
rect 37550 8576 37556 8588
rect 37608 8576 37614 8628
rect 38470 8576 38476 8628
rect 38528 8616 38534 8628
rect 38749 8619 38807 8625
rect 38749 8616 38761 8619
rect 38528 8588 38761 8616
rect 38528 8576 38534 8588
rect 38749 8585 38761 8588
rect 38795 8585 38807 8619
rect 42794 8616 42800 8628
rect 38749 8579 38807 8585
rect 41156 8588 42800 8616
rect 36722 8508 36728 8560
rect 36780 8508 36786 8560
rect 37093 8551 37151 8557
rect 37093 8517 37105 8551
rect 37139 8548 37151 8551
rect 37182 8548 37188 8560
rect 37139 8520 37188 8548
rect 37139 8517 37151 8520
rect 37093 8511 37151 8517
rect 37182 8508 37188 8520
rect 37240 8508 37246 8560
rect 37274 8508 37280 8560
rect 37332 8508 37338 8560
rect 38102 8508 38108 8560
rect 38160 8548 38166 8560
rect 38381 8551 38439 8557
rect 38381 8548 38393 8551
rect 38160 8520 38393 8548
rect 38160 8508 38166 8520
rect 38381 8517 38393 8520
rect 38427 8548 38439 8551
rect 41156 8548 41184 8588
rect 41340 8557 41368 8588
rect 42794 8576 42800 8588
rect 42852 8576 42858 8628
rect 43162 8576 43168 8628
rect 43220 8616 43226 8628
rect 43441 8619 43499 8625
rect 43441 8616 43453 8619
rect 43220 8588 43453 8616
rect 43220 8576 43226 8588
rect 43441 8585 43453 8588
rect 43487 8585 43499 8619
rect 43441 8579 43499 8585
rect 43530 8576 43536 8628
rect 43588 8616 43594 8628
rect 45462 8616 45468 8628
rect 43588 8588 44312 8616
rect 43588 8576 43594 8588
rect 38427 8520 41184 8548
rect 41233 8551 41291 8557
rect 38427 8517 38439 8520
rect 38381 8511 38439 8517
rect 41233 8517 41245 8551
rect 41279 8517 41291 8551
rect 41233 8511 41291 8517
rect 41325 8551 41383 8557
rect 41325 8517 41337 8551
rect 41371 8517 41383 8551
rect 41325 8511 41383 8517
rect 37461 8483 37519 8489
rect 37461 8480 37473 8483
rect 36320 8452 36365 8480
rect 36464 8452 37473 8480
rect 36320 8443 36328 8452
rect 37461 8449 37473 8452
rect 37507 8449 37519 8483
rect 37461 8443 37519 8449
rect 36320 8440 36326 8443
rect 37550 8440 37556 8492
rect 37608 8440 37614 8492
rect 37642 8440 37648 8492
rect 37700 8480 37706 8492
rect 38197 8483 38255 8489
rect 38197 8480 38209 8483
rect 37700 8452 38209 8480
rect 37700 8440 37706 8452
rect 38197 8449 38209 8452
rect 38243 8449 38255 8483
rect 38197 8443 38255 8449
rect 38473 8483 38531 8489
rect 38473 8449 38485 8483
rect 38519 8449 38531 8483
rect 38473 8443 38531 8449
rect 38565 8483 38623 8489
rect 38565 8449 38577 8483
rect 38611 8449 38623 8483
rect 38565 8443 38623 8449
rect 40589 8483 40647 8489
rect 40589 8449 40601 8483
rect 40635 8480 40647 8483
rect 41136 8483 41194 8489
rect 40635 8452 41000 8480
rect 40635 8449 40647 8452
rect 40589 8443 40647 8449
rect 37182 8412 37188 8424
rect 35360 8384 35664 8412
rect 36096 8384 37188 8412
rect 35434 8344 35440 8356
rect 35084 8316 35440 8344
rect 35434 8304 35440 8316
rect 35492 8304 35498 8356
rect 30374 8236 30380 8288
rect 30432 8276 30438 8288
rect 30837 8279 30895 8285
rect 30837 8276 30849 8279
rect 30432 8248 30849 8276
rect 30432 8236 30438 8248
rect 30837 8245 30849 8248
rect 30883 8245 30895 8279
rect 35636 8276 35664 8384
rect 37182 8372 37188 8384
rect 37240 8372 37246 8424
rect 37274 8372 37280 8424
rect 37332 8412 37338 8424
rect 38488 8412 38516 8443
rect 37332 8384 38516 8412
rect 37332 8372 37338 8384
rect 35713 8347 35771 8353
rect 35713 8313 35725 8347
rect 35759 8344 35771 8347
rect 36817 8347 36875 8353
rect 35759 8316 36768 8344
rect 35759 8313 35771 8316
rect 35713 8307 35771 8313
rect 36078 8276 36084 8288
rect 35636 8248 36084 8276
rect 30837 8239 30895 8245
rect 36078 8236 36084 8248
rect 36136 8236 36142 8288
rect 36740 8276 36768 8316
rect 36817 8313 36829 8347
rect 36863 8344 36875 8347
rect 37458 8344 37464 8356
rect 36863 8316 37464 8344
rect 36863 8313 36875 8316
rect 36817 8307 36875 8313
rect 37458 8304 37464 8316
rect 37516 8304 37522 8356
rect 37737 8347 37795 8353
rect 37737 8313 37749 8347
rect 37783 8344 37795 8347
rect 38010 8344 38016 8356
rect 37783 8316 38016 8344
rect 37783 8313 37795 8316
rect 37737 8307 37795 8313
rect 38010 8304 38016 8316
rect 38068 8304 38074 8356
rect 38580 8344 38608 8443
rect 40310 8372 40316 8424
rect 40368 8412 40374 8424
rect 40773 8415 40831 8421
rect 40773 8412 40785 8415
rect 40368 8384 40785 8412
rect 40368 8372 40374 8384
rect 40773 8381 40785 8384
rect 40819 8381 40831 8415
rect 40773 8375 40831 8381
rect 40862 8372 40868 8424
rect 40920 8372 40926 8424
rect 38488 8316 38608 8344
rect 37277 8279 37335 8285
rect 37277 8276 37289 8279
rect 36740 8248 37289 8276
rect 37277 8245 37289 8248
rect 37323 8245 37335 8279
rect 37277 8239 37335 8245
rect 37366 8236 37372 8288
rect 37424 8276 37430 8288
rect 38286 8276 38292 8288
rect 37424 8248 38292 8276
rect 37424 8236 37430 8248
rect 38286 8236 38292 8248
rect 38344 8276 38350 8288
rect 38488 8276 38516 8316
rect 39206 8304 39212 8356
rect 39264 8344 39270 8356
rect 40972 8353 41000 8452
rect 41136 8449 41148 8483
rect 41182 8449 41194 8483
rect 41248 8480 41276 8511
rect 41414 8508 41420 8560
rect 41472 8548 41478 8560
rect 41472 8520 41644 8548
rect 41472 8508 41478 8520
rect 41506 8480 41512 8492
rect 41248 8452 41414 8480
rect 41467 8452 41512 8480
rect 41136 8443 41194 8449
rect 40957 8347 41015 8353
rect 39264 8316 40540 8344
rect 39264 8304 39270 8316
rect 39224 8276 39252 8304
rect 38344 8248 39252 8276
rect 38344 8236 38350 8248
rect 40126 8236 40132 8288
rect 40184 8276 40190 8288
rect 40405 8279 40463 8285
rect 40405 8276 40417 8279
rect 40184 8248 40417 8276
rect 40184 8236 40190 8248
rect 40405 8245 40417 8248
rect 40451 8245 40463 8279
rect 40512 8276 40540 8316
rect 40957 8313 40969 8347
rect 41003 8313 41015 8347
rect 40957 8307 41015 8313
rect 41151 8276 41179 8443
rect 41386 8412 41414 8452
rect 41506 8440 41512 8452
rect 41564 8440 41570 8492
rect 41616 8489 41644 8520
rect 41690 8508 41696 8560
rect 41748 8548 41754 8560
rect 41748 8520 43116 8548
rect 41748 8508 41754 8520
rect 41601 8483 41659 8489
rect 41601 8449 41613 8483
rect 41647 8449 41659 8483
rect 41601 8443 41659 8449
rect 42334 8440 42340 8492
rect 42392 8480 42398 8492
rect 42429 8483 42487 8489
rect 42429 8480 42441 8483
rect 42392 8452 42441 8480
rect 42392 8440 42398 8452
rect 42429 8449 42441 8452
rect 42475 8449 42487 8483
rect 42429 8443 42487 8449
rect 42610 8440 42616 8492
rect 42668 8440 42674 8492
rect 42702 8440 42708 8492
rect 42760 8440 42766 8492
rect 42886 8440 42892 8492
rect 42944 8440 42950 8492
rect 42978 8440 42984 8492
rect 43036 8440 43042 8492
rect 43088 8489 43116 8520
rect 43714 8508 43720 8560
rect 43772 8548 43778 8560
rect 44284 8557 44312 8588
rect 44376 8588 45468 8616
rect 43901 8551 43959 8557
rect 43901 8548 43913 8551
rect 43772 8520 43913 8548
rect 43772 8508 43778 8520
rect 43901 8517 43913 8520
rect 43947 8517 43959 8551
rect 43901 8511 43959 8517
rect 44269 8551 44327 8557
rect 44269 8517 44281 8551
rect 44315 8517 44327 8551
rect 44269 8511 44327 8517
rect 43078 8483 43136 8489
rect 43078 8449 43090 8483
rect 43124 8480 43136 8483
rect 43346 8480 43352 8492
rect 43124 8452 43352 8480
rect 43124 8449 43136 8452
rect 43078 8443 43136 8449
rect 43346 8440 43352 8452
rect 43404 8440 43410 8492
rect 43625 8483 43683 8489
rect 43625 8449 43637 8483
rect 43671 8480 43683 8483
rect 43806 8480 43812 8492
rect 43671 8452 43812 8480
rect 43671 8449 43683 8452
rect 43625 8443 43683 8449
rect 43806 8440 43812 8452
rect 43864 8440 43870 8492
rect 43993 8483 44051 8489
rect 43993 8449 44005 8483
rect 44039 8449 44051 8483
rect 43993 8443 44051 8449
rect 42720 8412 42748 8440
rect 41386 8384 42748 8412
rect 43714 8372 43720 8424
rect 43772 8372 43778 8424
rect 44008 8412 44036 8443
rect 44174 8440 44180 8492
rect 44232 8440 44238 8492
rect 44376 8489 44404 8588
rect 45462 8576 45468 8588
rect 45520 8576 45526 8628
rect 45649 8619 45707 8625
rect 45649 8585 45661 8619
rect 45695 8585 45707 8619
rect 48774 8616 48780 8628
rect 45649 8579 45707 8585
rect 45848 8588 48780 8616
rect 45005 8551 45063 8557
rect 44569 8520 44864 8548
rect 44361 8483 44419 8489
rect 44361 8449 44373 8483
rect 44407 8449 44419 8483
rect 44361 8443 44419 8449
rect 44569 8412 44597 8520
rect 44637 8483 44695 8489
rect 44637 8449 44649 8483
rect 44683 8449 44695 8483
rect 44637 8443 44695 8449
rect 44008 8384 44597 8412
rect 43257 8347 43315 8353
rect 43257 8313 43269 8347
rect 43303 8344 43315 8347
rect 43303 8316 43668 8344
rect 43303 8313 43315 8316
rect 43257 8307 43315 8313
rect 40512 8248 41179 8276
rect 40405 8239 40463 8245
rect 42058 8236 42064 8288
rect 42116 8276 42122 8288
rect 42702 8276 42708 8288
rect 42116 8248 42708 8276
rect 42116 8236 42122 8248
rect 42702 8236 42708 8248
rect 42760 8236 42766 8288
rect 43640 8285 43668 8316
rect 43625 8279 43683 8285
rect 43625 8245 43637 8279
rect 43671 8245 43683 8279
rect 43625 8239 43683 8245
rect 44545 8279 44603 8285
rect 44545 8245 44557 8279
rect 44591 8276 44603 8279
rect 44652 8276 44680 8443
rect 44726 8440 44732 8492
rect 44784 8440 44790 8492
rect 44836 8412 44864 8520
rect 45005 8517 45017 8551
rect 45051 8548 45063 8551
rect 45370 8548 45376 8560
rect 45051 8520 45376 8548
rect 45051 8517 45063 8520
rect 45005 8511 45063 8517
rect 45370 8508 45376 8520
rect 45428 8548 45434 8560
rect 45664 8548 45692 8579
rect 45428 8520 45692 8548
rect 45428 8508 45434 8520
rect 44910 8440 44916 8492
rect 44968 8440 44974 8492
rect 45094 8440 45100 8492
rect 45152 8489 45158 8492
rect 45152 8480 45160 8489
rect 45848 8480 45876 8588
rect 48774 8576 48780 8588
rect 48832 8576 48838 8628
rect 49513 8619 49571 8625
rect 49513 8585 49525 8619
rect 49559 8616 49571 8619
rect 50522 8616 50528 8628
rect 49559 8588 50528 8616
rect 49559 8585 49571 8588
rect 49513 8579 49571 8585
rect 50522 8576 50528 8588
rect 50580 8576 50586 8628
rect 50798 8576 50804 8628
rect 50856 8576 50862 8628
rect 50890 8576 50896 8628
rect 50948 8616 50954 8628
rect 50985 8619 51043 8625
rect 50985 8616 50997 8619
rect 50948 8588 50997 8616
rect 50948 8576 50954 8588
rect 50985 8585 50997 8588
rect 51031 8585 51043 8619
rect 50985 8579 51043 8585
rect 51166 8576 51172 8628
rect 51224 8576 51230 8628
rect 46566 8508 46572 8560
rect 46624 8508 46630 8560
rect 47210 8508 47216 8560
rect 47268 8548 47274 8560
rect 50540 8548 50568 8576
rect 50617 8551 50675 8557
rect 50617 8548 50629 8551
rect 47268 8520 48820 8548
rect 50540 8520 50629 8548
rect 47268 8508 47274 8520
rect 48792 8489 48820 8520
rect 50617 8517 50629 8520
rect 50663 8517 50675 8551
rect 50617 8511 50675 8517
rect 50706 8508 50712 8560
rect 50764 8508 50770 8560
rect 50816 8548 50844 8576
rect 50816 8520 51028 8548
rect 45152 8452 45876 8480
rect 48777 8483 48835 8489
rect 45152 8443 45160 8452
rect 48777 8449 48789 8483
rect 48823 8449 48835 8483
rect 48777 8443 48835 8449
rect 45152 8440 45158 8443
rect 48866 8440 48872 8492
rect 48924 8440 48930 8492
rect 49145 8483 49203 8489
rect 49145 8449 49157 8483
rect 49191 8480 49203 8483
rect 49605 8483 49663 8489
rect 49605 8480 49617 8483
rect 49191 8452 49617 8480
rect 49191 8449 49203 8452
rect 49145 8443 49203 8449
rect 49605 8449 49617 8452
rect 49651 8449 49663 8483
rect 49605 8443 49663 8449
rect 49786 8440 49792 8492
rect 49844 8480 49850 8492
rect 50522 8489 50528 8492
rect 50341 8483 50399 8489
rect 50341 8480 50353 8483
rect 49844 8452 50353 8480
rect 49844 8440 49850 8452
rect 50341 8449 50353 8452
rect 50387 8449 50399 8483
rect 50341 8443 50399 8449
rect 50489 8483 50528 8489
rect 50489 8449 50501 8483
rect 50489 8443 50528 8449
rect 50522 8440 50528 8443
rect 50580 8440 50586 8492
rect 50806 8483 50864 8489
rect 50806 8449 50818 8483
rect 50852 8449 50864 8483
rect 51000 8480 51028 8520
rect 51074 8508 51080 8560
rect 51132 8548 51138 8560
rect 51537 8551 51595 8557
rect 51537 8548 51549 8551
rect 51132 8520 51549 8548
rect 51132 8508 51138 8520
rect 51537 8517 51549 8520
rect 51583 8548 51595 8551
rect 52178 8548 52184 8560
rect 51583 8520 52184 8548
rect 51583 8517 51595 8520
rect 51537 8511 51595 8517
rect 52178 8508 52184 8520
rect 52236 8508 52242 8560
rect 51000 8452 51212 8480
rect 50806 8443 50864 8449
rect 45646 8412 45652 8424
rect 44836 8384 45652 8412
rect 45646 8372 45652 8384
rect 45704 8372 45710 8424
rect 47118 8372 47124 8424
rect 47176 8372 47182 8424
rect 47397 8415 47455 8421
rect 47397 8381 47409 8415
rect 47443 8412 47455 8415
rect 48038 8412 48044 8424
rect 47443 8384 48044 8412
rect 47443 8381 47455 8384
rect 47397 8375 47455 8381
rect 44591 8248 44680 8276
rect 44591 8245 44603 8248
rect 44545 8239 44603 8245
rect 45278 8236 45284 8288
rect 45336 8236 45342 8288
rect 46934 8236 46940 8288
rect 46992 8276 46998 8288
rect 47412 8276 47440 8375
rect 48038 8372 48044 8384
rect 48096 8372 48102 8424
rect 48958 8372 48964 8424
rect 49016 8412 49022 8424
rect 49053 8415 49111 8421
rect 49053 8412 49065 8415
rect 49016 8384 49065 8412
rect 49016 8372 49022 8384
rect 49053 8381 49065 8384
rect 49099 8381 49111 8415
rect 49053 8375 49111 8381
rect 50246 8372 50252 8424
rect 50304 8372 50310 8424
rect 50614 8372 50620 8424
rect 50672 8412 50678 8424
rect 50821 8412 50849 8443
rect 50672 8384 50849 8412
rect 51184 8412 51212 8452
rect 51258 8440 51264 8492
rect 51316 8440 51322 8492
rect 51354 8483 51412 8489
rect 51354 8449 51366 8483
rect 51400 8449 51412 8483
rect 51354 8443 51412 8449
rect 51369 8412 51397 8443
rect 51626 8440 51632 8492
rect 51684 8440 51690 8492
rect 51718 8440 51724 8492
rect 51776 8489 51782 8492
rect 51776 8480 51784 8489
rect 51776 8452 51821 8480
rect 51776 8443 51784 8452
rect 51776 8440 51782 8443
rect 53466 8440 53472 8492
rect 53524 8440 53530 8492
rect 54846 8480 54852 8492
rect 53668 8452 54852 8480
rect 51184 8384 51397 8412
rect 51644 8412 51672 8440
rect 53668 8412 53696 8452
rect 54846 8440 54852 8452
rect 54904 8480 54910 8492
rect 54941 8483 54999 8489
rect 54941 8480 54953 8483
rect 54904 8452 54953 8480
rect 54904 8440 54910 8452
rect 54941 8449 54953 8452
rect 54987 8449 54999 8483
rect 54941 8443 54999 8449
rect 78030 8440 78036 8492
rect 78088 8440 78094 8492
rect 51644 8384 53696 8412
rect 53745 8415 53803 8421
rect 50672 8372 50678 8384
rect 53745 8381 53757 8415
rect 53791 8412 53803 8415
rect 54389 8415 54447 8421
rect 54389 8412 54401 8415
rect 53791 8384 54401 8412
rect 53791 8381 53803 8384
rect 53745 8375 53803 8381
rect 54389 8381 54401 8384
rect 54435 8381 54447 8415
rect 54389 8375 54447 8381
rect 51258 8304 51264 8356
rect 51316 8344 51322 8356
rect 51994 8344 52000 8356
rect 51316 8316 52000 8344
rect 51316 8304 51322 8316
rect 51994 8304 52000 8316
rect 52052 8304 52058 8356
rect 52914 8304 52920 8356
rect 52972 8344 52978 8356
rect 53009 8347 53067 8353
rect 53009 8344 53021 8347
rect 52972 8316 53021 8344
rect 52972 8304 52978 8316
rect 53009 8313 53021 8316
rect 53055 8313 53067 8347
rect 53009 8307 53067 8313
rect 53558 8304 53564 8356
rect 53616 8344 53622 8356
rect 53653 8347 53711 8353
rect 53653 8344 53665 8347
rect 53616 8316 53665 8344
rect 53616 8304 53622 8316
rect 53653 8313 53665 8316
rect 53699 8313 53711 8347
rect 53653 8307 53711 8313
rect 78214 8304 78220 8356
rect 78272 8304 78278 8356
rect 46992 8248 47440 8276
rect 46992 8236 46998 8248
rect 48498 8236 48504 8288
rect 48556 8276 48562 8288
rect 48593 8279 48651 8285
rect 48593 8276 48605 8279
rect 48556 8248 48605 8276
rect 48556 8236 48562 8248
rect 48593 8245 48605 8248
rect 48639 8245 48651 8279
rect 48593 8239 48651 8245
rect 50062 8236 50068 8288
rect 50120 8276 50126 8288
rect 50890 8276 50896 8288
rect 50120 8248 50896 8276
rect 50120 8236 50126 8248
rect 50890 8236 50896 8248
rect 50948 8236 50954 8288
rect 51718 8236 51724 8288
rect 51776 8276 51782 8288
rect 51905 8279 51963 8285
rect 51905 8276 51917 8279
rect 51776 8248 51917 8276
rect 51776 8236 51782 8248
rect 51905 8245 51917 8248
rect 51951 8245 51963 8279
rect 51905 8239 51963 8245
rect 53282 8236 53288 8288
rect 53340 8236 53346 8288
rect 1104 8186 78844 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 78844 8186
rect 1104 8112 78844 8134
rect 29178 8032 29184 8084
rect 29236 8072 29242 8084
rect 30193 8075 30251 8081
rect 30193 8072 30205 8075
rect 29236 8044 30205 8072
rect 29236 8032 29242 8044
rect 30193 8041 30205 8044
rect 30239 8041 30251 8075
rect 30193 8035 30251 8041
rect 35434 8032 35440 8084
rect 35492 8032 35498 8084
rect 35621 8075 35679 8081
rect 35621 8041 35633 8075
rect 35667 8072 35679 8075
rect 41601 8075 41659 8081
rect 35667 8044 41414 8072
rect 35667 8041 35679 8044
rect 35621 8035 35679 8041
rect 31110 7896 31116 7948
rect 31168 7936 31174 7948
rect 31389 7939 31447 7945
rect 31389 7936 31401 7939
rect 31168 7908 31401 7936
rect 31168 7896 31174 7908
rect 31389 7905 31401 7908
rect 31435 7936 31447 7939
rect 32306 7936 32312 7948
rect 31435 7908 32312 7936
rect 31435 7905 31447 7908
rect 31389 7899 31447 7905
rect 30374 7828 30380 7880
rect 30432 7828 30438 7880
rect 30558 7828 30564 7880
rect 30616 7828 30622 7880
rect 30653 7871 30711 7877
rect 30653 7837 30665 7871
rect 30699 7868 30711 7871
rect 30745 7871 30803 7877
rect 30745 7868 30757 7871
rect 30699 7840 30757 7868
rect 30699 7837 30711 7840
rect 30653 7831 30711 7837
rect 30745 7837 30757 7840
rect 30791 7837 30803 7871
rect 30745 7831 30803 7837
rect 31018 7828 31024 7880
rect 31076 7868 31082 7880
rect 31478 7868 31484 7880
rect 31076 7840 31484 7868
rect 31076 7828 31082 7840
rect 31478 7828 31484 7840
rect 31536 7868 31542 7880
rect 31662 7868 31668 7880
rect 31536 7840 31668 7868
rect 31536 7828 31542 7840
rect 31662 7828 31668 7840
rect 31720 7828 31726 7880
rect 31757 7871 31815 7877
rect 31757 7837 31769 7871
rect 31803 7868 31815 7871
rect 31956 7868 31984 7908
rect 32306 7896 32312 7908
rect 32364 7896 32370 7948
rect 31803 7840 31984 7868
rect 31803 7837 31815 7840
rect 31757 7831 31815 7837
rect 32030 7828 32036 7880
rect 32088 7828 32094 7880
rect 34422 7828 34428 7880
rect 34480 7868 34486 7880
rect 34885 7871 34943 7877
rect 34885 7868 34897 7871
rect 34480 7840 34897 7868
rect 34480 7828 34486 7840
rect 34885 7837 34897 7840
rect 34931 7837 34943 7871
rect 35253 7871 35311 7877
rect 34885 7831 34943 7837
rect 34992 7840 35204 7868
rect 31849 7803 31907 7809
rect 31849 7769 31861 7803
rect 31895 7800 31907 7803
rect 32582 7800 32588 7812
rect 31895 7772 32588 7800
rect 31895 7769 31907 7772
rect 31849 7763 31907 7769
rect 31018 7692 31024 7744
rect 31076 7732 31082 7744
rect 31481 7735 31539 7741
rect 31481 7732 31493 7735
rect 31076 7704 31493 7732
rect 31076 7692 31082 7704
rect 31481 7701 31493 7704
rect 31527 7701 31539 7735
rect 31481 7695 31539 7701
rect 31754 7692 31760 7744
rect 31812 7732 31818 7744
rect 31864 7732 31892 7763
rect 32582 7760 32588 7772
rect 32640 7760 32646 7812
rect 34698 7760 34704 7812
rect 34756 7800 34762 7812
rect 34992 7800 35020 7840
rect 35176 7809 35204 7840
rect 35253 7837 35265 7871
rect 35299 7868 35311 7871
rect 35636 7868 35664 8035
rect 36078 7964 36084 8016
rect 36136 7964 36142 8016
rect 36262 7964 36268 8016
rect 36320 8004 36326 8016
rect 36541 8007 36599 8013
rect 36541 8004 36553 8007
rect 36320 7976 36553 8004
rect 36320 7964 36326 7976
rect 36541 7973 36553 7976
rect 36587 7973 36599 8007
rect 41386 8004 41414 8044
rect 41601 8041 41613 8075
rect 41647 8072 41659 8075
rect 41966 8072 41972 8084
rect 41647 8044 41972 8072
rect 41647 8041 41659 8044
rect 41601 8035 41659 8041
rect 41966 8032 41972 8044
rect 42024 8032 42030 8084
rect 42610 8032 42616 8084
rect 42668 8032 42674 8084
rect 42797 8075 42855 8081
rect 42797 8041 42809 8075
rect 42843 8072 42855 8075
rect 43070 8072 43076 8084
rect 42843 8044 43076 8072
rect 42843 8041 42855 8044
rect 42797 8035 42855 8041
rect 41874 8004 41880 8016
rect 36541 7967 36599 7973
rect 37200 7976 39160 8004
rect 41386 7976 41880 8004
rect 35894 7896 35900 7948
rect 35952 7936 35958 7948
rect 37200 7936 37228 7976
rect 35952 7908 37228 7936
rect 35952 7896 35958 7908
rect 37274 7896 37280 7948
rect 37332 7936 37338 7948
rect 37642 7936 37648 7948
rect 37332 7908 37648 7936
rect 37332 7896 37338 7908
rect 37642 7896 37648 7908
rect 37700 7896 37706 7948
rect 38470 7896 38476 7948
rect 38528 7896 38534 7948
rect 35299 7840 35664 7868
rect 38289 7871 38347 7877
rect 35299 7837 35311 7840
rect 35253 7831 35311 7837
rect 38289 7837 38301 7871
rect 38335 7868 38347 7871
rect 38381 7871 38439 7877
rect 38381 7868 38393 7871
rect 38335 7840 38393 7868
rect 38335 7837 38347 7840
rect 38289 7831 38347 7837
rect 38381 7837 38393 7840
rect 38427 7837 38439 7871
rect 38381 7831 38439 7837
rect 38657 7871 38715 7877
rect 38657 7837 38669 7871
rect 38703 7837 38715 7871
rect 38657 7831 38715 7837
rect 38749 7871 38807 7877
rect 38749 7837 38761 7871
rect 38795 7868 38807 7871
rect 38838 7868 38844 7880
rect 38795 7840 38844 7868
rect 38795 7837 38807 7840
rect 38749 7831 38807 7837
rect 34756 7772 35020 7800
rect 35069 7803 35127 7809
rect 34756 7760 34762 7772
rect 35069 7769 35081 7803
rect 35115 7769 35127 7803
rect 35069 7763 35127 7769
rect 35161 7803 35219 7809
rect 35161 7769 35173 7803
rect 35207 7769 35219 7803
rect 38672 7800 38700 7831
rect 38838 7828 38844 7840
rect 38896 7828 38902 7880
rect 39025 7803 39083 7809
rect 39025 7800 39037 7803
rect 38672 7772 39037 7800
rect 35161 7763 35219 7769
rect 39025 7769 39037 7772
rect 39071 7769 39083 7803
rect 39025 7763 39083 7769
rect 31812 7704 31892 7732
rect 35084 7732 35112 7763
rect 36265 7735 36323 7741
rect 36265 7732 36277 7735
rect 35084 7704 36277 7732
rect 31812 7692 31818 7704
rect 36265 7701 36277 7704
rect 36311 7732 36323 7735
rect 38654 7732 38660 7744
rect 36311 7704 38660 7732
rect 36311 7701 36323 7704
rect 36265 7695 36323 7701
rect 38654 7692 38660 7704
rect 38712 7692 38718 7744
rect 38746 7692 38752 7744
rect 38804 7732 38810 7744
rect 38933 7735 38991 7741
rect 38933 7732 38945 7735
rect 38804 7704 38945 7732
rect 38804 7692 38810 7704
rect 38933 7701 38945 7704
rect 38979 7701 38991 7735
rect 39132 7732 39160 7976
rect 41874 7964 41880 7976
rect 41932 7964 41938 8016
rect 39850 7896 39856 7948
rect 39908 7896 39914 7948
rect 40126 7896 40132 7948
rect 40184 7896 40190 7948
rect 41892 7936 41920 7964
rect 42889 7939 42947 7945
rect 42889 7936 42901 7939
rect 41892 7908 42901 7936
rect 39206 7828 39212 7880
rect 39264 7828 39270 7880
rect 39298 7828 39304 7880
rect 39356 7828 39362 7880
rect 41230 7828 41236 7880
rect 41288 7828 41294 7880
rect 41874 7828 41880 7880
rect 41932 7868 41938 7880
rect 42260 7877 42288 7908
rect 42889 7905 42901 7908
rect 42935 7905 42947 7939
rect 42889 7899 42947 7905
rect 42061 7871 42119 7877
rect 42061 7868 42073 7871
rect 41932 7840 42073 7868
rect 41932 7828 41938 7840
rect 42061 7837 42073 7840
rect 42107 7837 42119 7871
rect 42061 7831 42119 7837
rect 42245 7871 42303 7877
rect 42245 7837 42257 7871
rect 42291 7837 42303 7871
rect 42245 7831 42303 7837
rect 42429 7871 42487 7877
rect 42429 7837 42441 7871
rect 42475 7868 42487 7871
rect 42996 7868 43024 8044
rect 43070 8032 43076 8044
rect 43128 8032 43134 8084
rect 43346 8032 43352 8084
rect 43404 8032 43410 8084
rect 44545 8075 44603 8081
rect 44545 8041 44557 8075
rect 44591 8072 44603 8075
rect 45094 8072 45100 8084
rect 44591 8044 45100 8072
rect 44591 8041 44603 8044
rect 44545 8035 44603 8041
rect 45094 8032 45100 8044
rect 45152 8032 45158 8084
rect 45922 8032 45928 8084
rect 45980 8032 45986 8084
rect 47118 8032 47124 8084
rect 47176 8072 47182 8084
rect 47305 8075 47363 8081
rect 47305 8072 47317 8075
rect 47176 8044 47317 8072
rect 47176 8032 47182 8044
rect 47305 8041 47317 8044
rect 47351 8041 47363 8075
rect 47305 8035 47363 8041
rect 49970 8032 49976 8084
rect 50028 8072 50034 8084
rect 50246 8072 50252 8084
rect 50028 8044 50252 8072
rect 50028 8032 50034 8044
rect 50246 8032 50252 8044
rect 50304 8032 50310 8084
rect 50798 8032 50804 8084
rect 50856 8072 50862 8084
rect 51258 8072 51264 8084
rect 50856 8044 51264 8072
rect 50856 8032 50862 8044
rect 51258 8032 51264 8044
rect 51316 8032 51322 8084
rect 51442 8032 51448 8084
rect 51500 8072 51506 8084
rect 52178 8072 52184 8084
rect 51500 8044 52184 8072
rect 51500 8032 51506 8044
rect 52178 8032 52184 8044
rect 52236 8072 52242 8084
rect 52917 8075 52975 8081
rect 52917 8072 52929 8075
rect 52236 8044 52929 8072
rect 52236 8032 52242 8044
rect 52917 8041 52929 8044
rect 52963 8041 52975 8075
rect 52917 8035 52975 8041
rect 54846 8032 54852 8084
rect 54904 8072 54910 8084
rect 54904 8044 55904 8072
rect 54904 8032 54910 8044
rect 44174 7964 44180 8016
rect 44232 8004 44238 8016
rect 45005 8007 45063 8013
rect 45005 8004 45017 8007
rect 44232 7976 45017 8004
rect 44232 7964 44238 7976
rect 45005 7973 45017 7976
rect 45051 7973 45063 8007
rect 45005 7967 45063 7973
rect 55033 8007 55091 8013
rect 55033 7973 55045 8007
rect 55079 8004 55091 8007
rect 55766 8004 55772 8016
rect 55079 7976 55772 8004
rect 55079 7973 55091 7976
rect 55033 7967 55091 7973
rect 55766 7964 55772 7976
rect 55824 7964 55830 8016
rect 46017 7939 46075 7945
rect 46017 7936 46029 7939
rect 45388 7908 46029 7936
rect 45388 7880 45416 7908
rect 46017 7905 46029 7908
rect 46063 7905 46075 7939
rect 46017 7899 46075 7905
rect 46842 7896 46848 7948
rect 46900 7896 46906 7948
rect 48038 7896 48044 7948
rect 48096 7936 48102 7948
rect 48225 7939 48283 7945
rect 48225 7936 48237 7939
rect 48096 7908 48237 7936
rect 48096 7896 48102 7908
rect 48225 7905 48237 7908
rect 48271 7905 48283 7939
rect 48225 7899 48283 7905
rect 48498 7896 48504 7948
rect 48556 7896 48562 7948
rect 50249 7939 50307 7945
rect 50249 7905 50261 7939
rect 50295 7936 50307 7939
rect 50614 7936 50620 7948
rect 50295 7908 50620 7936
rect 50295 7905 50307 7908
rect 50249 7899 50307 7905
rect 50614 7896 50620 7908
rect 50672 7896 50678 7948
rect 51169 7939 51227 7945
rect 51169 7905 51181 7939
rect 51215 7936 51227 7939
rect 51810 7936 51816 7948
rect 51215 7908 51816 7936
rect 51215 7905 51227 7908
rect 51169 7899 51227 7905
rect 51810 7896 51816 7908
rect 51868 7896 51874 7948
rect 53101 7939 53159 7945
rect 53101 7905 53113 7939
rect 53147 7936 53159 7939
rect 53374 7936 53380 7948
rect 53147 7908 53380 7936
rect 53147 7905 53159 7908
rect 53101 7899 53159 7905
rect 53374 7896 53380 7908
rect 53432 7896 53438 7948
rect 54018 7896 54024 7948
rect 54076 7936 54082 7948
rect 54662 7936 54668 7948
rect 54076 7908 54668 7936
rect 54076 7896 54082 7908
rect 54662 7896 54668 7908
rect 54720 7936 54726 7948
rect 54720 7908 55720 7936
rect 54720 7896 54726 7908
rect 42475 7840 43024 7868
rect 42475 7837 42487 7840
rect 42429 7831 42487 7837
rect 42334 7760 42340 7812
rect 42392 7760 42398 7812
rect 42444 7732 42472 7831
rect 45370 7828 45376 7880
rect 45428 7828 45434 7880
rect 45646 7828 45652 7880
rect 45704 7828 45710 7880
rect 45738 7828 45744 7880
rect 45796 7828 45802 7880
rect 46661 7871 46719 7877
rect 46661 7837 46673 7871
rect 46707 7868 46719 7871
rect 46753 7871 46811 7877
rect 46753 7868 46765 7871
rect 46707 7840 46765 7868
rect 46707 7837 46719 7840
rect 46661 7831 46719 7837
rect 46753 7837 46765 7840
rect 46799 7837 46811 7871
rect 46753 7831 46811 7837
rect 47029 7871 47087 7877
rect 47029 7837 47041 7871
rect 47075 7837 47087 7871
rect 47029 7831 47087 7837
rect 42610 7760 42616 7812
rect 42668 7800 42674 7812
rect 45557 7803 45615 7809
rect 45557 7800 45569 7803
rect 42668 7772 45569 7800
rect 42668 7760 42674 7772
rect 45557 7769 45569 7772
rect 45603 7800 45615 7803
rect 45830 7800 45836 7812
rect 45603 7772 45836 7800
rect 45603 7769 45615 7772
rect 45557 7763 45615 7769
rect 45830 7760 45836 7772
rect 45888 7760 45894 7812
rect 47044 7800 47072 7831
rect 47118 7828 47124 7880
rect 47176 7828 47182 7880
rect 47581 7871 47639 7877
rect 47581 7837 47593 7871
rect 47627 7837 47639 7871
rect 47581 7831 47639 7837
rect 47397 7803 47455 7809
rect 47397 7800 47409 7803
rect 47044 7772 47409 7800
rect 47397 7769 47409 7772
rect 47443 7769 47455 7803
rect 47397 7763 47455 7769
rect 39132 7704 42472 7732
rect 38933 7695 38991 7701
rect 42702 7692 42708 7744
rect 42760 7732 42766 7744
rect 47596 7732 47624 7831
rect 47670 7828 47676 7880
rect 47728 7828 47734 7880
rect 54938 7868 54944 7880
rect 54680 7840 54944 7868
rect 48222 7760 48228 7812
rect 48280 7800 48286 7812
rect 51445 7803 51503 7809
rect 48280 7772 48990 7800
rect 48280 7760 48286 7772
rect 42760 7704 47624 7732
rect 48884 7732 48912 7772
rect 51445 7769 51457 7803
rect 51491 7800 51503 7803
rect 51534 7800 51540 7812
rect 51491 7772 51540 7800
rect 51491 7769 51503 7772
rect 51445 7763 51503 7769
rect 51534 7760 51540 7772
rect 51592 7760 51598 7812
rect 52670 7772 52776 7800
rect 50341 7735 50399 7741
rect 50341 7732 50353 7735
rect 48884 7704 50353 7732
rect 42760 7692 42766 7704
rect 50341 7701 50353 7704
rect 50387 7732 50399 7735
rect 52748 7732 52776 7772
rect 53282 7760 53288 7812
rect 53340 7800 53346 7812
rect 53377 7803 53435 7809
rect 53377 7800 53389 7803
rect 53340 7772 53389 7800
rect 53340 7760 53346 7772
rect 53377 7769 53389 7772
rect 53423 7769 53435 7803
rect 53377 7763 53435 7769
rect 53576 7772 53866 7800
rect 52914 7732 52920 7744
rect 50387 7704 52920 7732
rect 50387 7701 50399 7704
rect 50341 7695 50399 7701
rect 52914 7692 52920 7704
rect 52972 7732 52978 7744
rect 53576 7732 53604 7772
rect 52972 7704 53604 7732
rect 52972 7692 52978 7704
rect 53650 7692 53656 7744
rect 53708 7732 53714 7744
rect 54680 7732 54708 7840
rect 54938 7828 54944 7840
rect 54996 7868 55002 7880
rect 55692 7877 55720 7908
rect 55876 7877 55904 8044
rect 78030 8032 78036 8084
rect 78088 8032 78094 8084
rect 77757 8007 77815 8013
rect 77757 7973 77769 8007
rect 77803 7973 77815 8007
rect 77757 7967 77815 7973
rect 77772 7936 77800 7967
rect 77772 7908 78260 7936
rect 78232 7877 78260 7908
rect 55493 7871 55551 7877
rect 55493 7868 55505 7871
rect 54996 7840 55505 7868
rect 54996 7828 55002 7840
rect 55493 7837 55505 7840
rect 55539 7837 55551 7871
rect 55493 7831 55551 7837
rect 55677 7871 55735 7877
rect 55677 7837 55689 7871
rect 55723 7837 55735 7871
rect 55677 7831 55735 7837
rect 55861 7871 55919 7877
rect 55861 7837 55873 7871
rect 55907 7837 55919 7871
rect 55861 7831 55919 7837
rect 77573 7871 77631 7877
rect 77573 7837 77585 7871
rect 77619 7868 77631 7871
rect 77849 7871 77907 7877
rect 77849 7868 77861 7871
rect 77619 7840 77861 7868
rect 77619 7837 77631 7840
rect 77573 7831 77631 7837
rect 77849 7837 77861 7840
rect 77895 7837 77907 7871
rect 77849 7831 77907 7837
rect 78217 7871 78275 7877
rect 78217 7837 78229 7871
rect 78263 7837 78275 7871
rect 78217 7831 78275 7837
rect 55582 7760 55588 7812
rect 55640 7760 55646 7812
rect 53708 7704 54708 7732
rect 53708 7692 53714 7704
rect 55030 7692 55036 7744
rect 55088 7732 55094 7744
rect 55309 7735 55367 7741
rect 55309 7732 55321 7735
rect 55088 7704 55321 7732
rect 55088 7692 55094 7704
rect 55309 7701 55321 7704
rect 55355 7701 55367 7735
rect 55309 7695 55367 7701
rect 77297 7735 77355 7741
rect 77297 7701 77309 7735
rect 77343 7732 77355 7735
rect 77389 7735 77447 7741
rect 77389 7732 77401 7735
rect 77343 7704 77401 7732
rect 77343 7701 77355 7704
rect 77297 7695 77355 7701
rect 77389 7701 77401 7704
rect 77435 7732 77447 7735
rect 77588 7732 77616 7831
rect 77662 7732 77668 7744
rect 77435 7704 77668 7732
rect 77435 7701 77447 7704
rect 77389 7695 77447 7701
rect 77662 7692 77668 7704
rect 77720 7692 77726 7744
rect 78398 7692 78404 7744
rect 78456 7692 78462 7744
rect 1104 7642 78844 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 66314 7642
rect 66366 7590 66378 7642
rect 66430 7590 66442 7642
rect 66494 7590 66506 7642
rect 66558 7590 66570 7642
rect 66622 7590 78844 7642
rect 1104 7568 78844 7590
rect 31757 7531 31815 7537
rect 31757 7497 31769 7531
rect 31803 7528 31815 7531
rect 31846 7528 31852 7540
rect 31803 7500 31852 7528
rect 31803 7497 31815 7500
rect 31757 7491 31815 7497
rect 31846 7488 31852 7500
rect 31904 7488 31910 7540
rect 37274 7488 37280 7540
rect 37332 7488 37338 7540
rect 38654 7488 38660 7540
rect 38712 7528 38718 7540
rect 40770 7528 40776 7540
rect 38712 7500 40776 7528
rect 38712 7488 38718 7500
rect 40770 7488 40776 7500
rect 40828 7488 40834 7540
rect 42518 7488 42524 7540
rect 42576 7528 42582 7540
rect 43257 7531 43315 7537
rect 43257 7528 43269 7531
rect 42576 7500 43269 7528
rect 42576 7488 42582 7500
rect 43257 7497 43269 7500
rect 43303 7528 43315 7531
rect 43993 7531 44051 7537
rect 43303 7500 43852 7528
rect 43303 7497 43315 7500
rect 43257 7491 43315 7497
rect 37366 7420 37372 7472
rect 37424 7460 37430 7472
rect 37424 7432 37582 7460
rect 37424 7420 37430 7432
rect 41966 7420 41972 7472
rect 42024 7460 42030 7472
rect 42705 7463 42763 7469
rect 42705 7460 42717 7463
rect 42024 7432 42717 7460
rect 42024 7420 42030 7432
rect 42705 7429 42717 7432
rect 42751 7429 42763 7463
rect 42705 7423 42763 7429
rect 42812 7432 43576 7460
rect 30926 7352 30932 7404
rect 30984 7352 30990 7404
rect 31018 7352 31024 7404
rect 31076 7352 31082 7404
rect 31297 7395 31355 7401
rect 31297 7361 31309 7395
rect 31343 7392 31355 7395
rect 32125 7395 32183 7401
rect 32125 7392 32137 7395
rect 31343 7364 32137 7392
rect 31343 7361 31355 7364
rect 31297 7355 31355 7361
rect 32125 7361 32137 7364
rect 32171 7361 32183 7395
rect 32125 7355 32183 7361
rect 32766 7352 32772 7404
rect 32824 7352 32830 7404
rect 33686 7392 33692 7404
rect 32876 7364 33692 7392
rect 30558 7284 30564 7336
rect 30616 7324 30622 7336
rect 31205 7327 31263 7333
rect 31205 7324 31217 7327
rect 30616 7296 31217 7324
rect 30616 7284 30622 7296
rect 31205 7293 31217 7296
rect 31251 7324 31263 7327
rect 32876 7324 32904 7364
rect 33686 7352 33692 7364
rect 33744 7352 33750 7404
rect 33870 7352 33876 7404
rect 33928 7352 33934 7404
rect 39025 7395 39083 7401
rect 39025 7361 39037 7395
rect 39071 7392 39083 7395
rect 39850 7392 39856 7404
rect 39071 7364 39856 7392
rect 39071 7361 39083 7364
rect 39025 7355 39083 7361
rect 39850 7352 39856 7364
rect 39908 7352 39914 7404
rect 40770 7352 40776 7404
rect 40828 7392 40834 7404
rect 41506 7392 41512 7404
rect 40828 7364 41512 7392
rect 40828 7352 40834 7364
rect 41506 7352 41512 7364
rect 41564 7352 41570 7404
rect 41690 7352 41696 7404
rect 41748 7392 41754 7404
rect 42334 7392 42340 7404
rect 41748 7364 42340 7392
rect 41748 7352 41754 7364
rect 42334 7352 42340 7364
rect 42392 7392 42398 7404
rect 42429 7395 42487 7401
rect 42429 7392 42441 7395
rect 42392 7364 42441 7392
rect 42392 7352 42398 7364
rect 42429 7361 42441 7364
rect 42475 7361 42487 7395
rect 42429 7355 42487 7361
rect 42610 7352 42616 7404
rect 42668 7352 42674 7404
rect 42812 7401 42840 7432
rect 42797 7395 42855 7401
rect 42797 7361 42809 7395
rect 42843 7361 42855 7395
rect 42797 7355 42855 7361
rect 43441 7395 43499 7401
rect 43441 7361 43453 7395
rect 43487 7361 43499 7395
rect 43441 7355 43499 7361
rect 31251 7296 32904 7324
rect 32953 7327 33011 7333
rect 31251 7293 31263 7296
rect 31205 7287 31263 7293
rect 32953 7293 32965 7327
rect 32999 7324 33011 7327
rect 33042 7324 33048 7336
rect 32999 7296 33048 7324
rect 32999 7293 33011 7296
rect 32953 7287 33011 7293
rect 33042 7284 33048 7296
rect 33100 7284 33106 7336
rect 33505 7327 33563 7333
rect 33505 7293 33517 7327
rect 33551 7324 33563 7327
rect 33597 7327 33655 7333
rect 33597 7324 33609 7327
rect 33551 7296 33609 7324
rect 33551 7293 33563 7296
rect 33505 7287 33563 7293
rect 33597 7293 33609 7296
rect 33643 7293 33655 7327
rect 33597 7287 33655 7293
rect 38746 7284 38752 7336
rect 38804 7284 38810 7336
rect 41524 7256 41552 7352
rect 41782 7284 41788 7336
rect 41840 7324 41846 7336
rect 42812 7324 42840 7355
rect 41840 7296 42840 7324
rect 41840 7284 41846 7296
rect 43346 7256 43352 7268
rect 41524 7228 43352 7256
rect 43346 7216 43352 7228
rect 43404 7216 43410 7268
rect 30742 7148 30748 7200
rect 30800 7148 30806 7200
rect 34054 7148 34060 7200
rect 34112 7148 34118 7200
rect 38746 7148 38752 7200
rect 38804 7188 38810 7200
rect 41414 7188 41420 7200
rect 38804 7160 41420 7188
rect 38804 7148 38810 7160
rect 41414 7148 41420 7160
rect 41472 7148 41478 7200
rect 42981 7191 43039 7197
rect 42981 7157 42993 7191
rect 43027 7188 43039 7191
rect 43070 7188 43076 7200
rect 43027 7160 43076 7188
rect 43027 7157 43039 7160
rect 42981 7151 43039 7157
rect 43070 7148 43076 7160
rect 43128 7148 43134 7200
rect 43456 7188 43484 7355
rect 43548 7256 43576 7432
rect 43625 7395 43683 7401
rect 43625 7361 43637 7395
rect 43671 7361 43683 7395
rect 43625 7355 43683 7361
rect 43640 7324 43668 7355
rect 43714 7352 43720 7404
rect 43772 7352 43778 7404
rect 43824 7401 43852 7500
rect 43993 7497 44005 7531
rect 44039 7528 44051 7531
rect 44450 7528 44456 7540
rect 44039 7500 44456 7528
rect 44039 7497 44051 7500
rect 43993 7491 44051 7497
rect 44450 7488 44456 7500
rect 44508 7488 44514 7540
rect 46474 7488 46480 7540
rect 46532 7528 46538 7540
rect 47670 7528 47676 7540
rect 46532 7500 47676 7528
rect 46532 7488 46538 7500
rect 47670 7488 47676 7500
rect 47728 7488 47734 7540
rect 51534 7488 51540 7540
rect 51592 7488 51598 7540
rect 53466 7488 53472 7540
rect 53524 7488 53530 7540
rect 53742 7488 53748 7540
rect 53800 7528 53806 7540
rect 54202 7528 54208 7540
rect 53800 7500 54208 7528
rect 53800 7488 53806 7500
rect 54202 7488 54208 7500
rect 54260 7528 54266 7540
rect 55030 7528 55036 7540
rect 54260 7500 54432 7528
rect 54260 7488 54266 7500
rect 49970 7420 49976 7472
rect 50028 7420 50034 7472
rect 50062 7420 50068 7472
rect 50120 7420 50126 7472
rect 53300 7432 53972 7460
rect 43809 7395 43867 7401
rect 43809 7361 43821 7395
rect 43855 7361 43867 7395
rect 43809 7355 43867 7361
rect 44177 7395 44235 7401
rect 44177 7361 44189 7395
rect 44223 7392 44235 7395
rect 44634 7392 44640 7404
rect 44223 7364 44640 7392
rect 44223 7361 44235 7364
rect 44177 7355 44235 7361
rect 44192 7324 44220 7355
rect 44634 7352 44640 7364
rect 44692 7352 44698 7404
rect 49878 7352 49884 7404
rect 49936 7352 49942 7404
rect 50249 7395 50307 7401
rect 50249 7361 50261 7395
rect 50295 7392 50307 7395
rect 50338 7392 50344 7404
rect 50295 7364 50344 7392
rect 50295 7361 50307 7364
rect 50249 7355 50307 7361
rect 50338 7352 50344 7364
rect 50396 7392 50402 7404
rect 51166 7392 51172 7404
rect 50396 7364 51172 7392
rect 50396 7352 50402 7364
rect 51166 7352 51172 7364
rect 51224 7352 51230 7404
rect 51718 7352 51724 7404
rect 51776 7352 51782 7404
rect 52178 7352 52184 7404
rect 52236 7392 52242 7404
rect 53300 7401 53328 7432
rect 53650 7401 53656 7404
rect 53285 7395 53343 7401
rect 53285 7392 53297 7395
rect 52236 7364 53297 7392
rect 52236 7352 52242 7364
rect 53285 7361 53297 7364
rect 53331 7361 53343 7395
rect 53648 7392 53656 7401
rect 53611 7364 53656 7392
rect 53285 7355 53343 7361
rect 53648 7355 53656 7364
rect 53650 7352 53656 7355
rect 53708 7352 53714 7404
rect 53742 7352 53748 7404
rect 53800 7352 53806 7404
rect 53834 7352 53840 7404
rect 53892 7352 53898 7404
rect 53944 7401 53972 7432
rect 53944 7395 54023 7401
rect 53944 7364 53977 7395
rect 53965 7361 53977 7364
rect 54011 7361 54023 7395
rect 53965 7355 54023 7361
rect 54110 7352 54116 7404
rect 54168 7352 54174 7404
rect 54404 7401 54432 7500
rect 54680 7500 55036 7528
rect 54680 7401 54708 7500
rect 55030 7488 55036 7500
rect 55088 7488 55094 7540
rect 54941 7463 54999 7469
rect 54941 7429 54953 7463
rect 54987 7460 54999 7463
rect 55309 7463 55367 7469
rect 55309 7460 55321 7463
rect 54987 7432 55321 7460
rect 54987 7429 54999 7432
rect 54941 7423 54999 7429
rect 55309 7429 55321 7432
rect 55355 7429 55367 7463
rect 55309 7423 55367 7429
rect 55766 7420 55772 7472
rect 55824 7420 55830 7472
rect 54389 7395 54447 7401
rect 54389 7361 54401 7395
rect 54435 7361 54447 7395
rect 54389 7355 54447 7361
rect 54665 7395 54723 7401
rect 54665 7361 54677 7395
rect 54711 7361 54723 7395
rect 54665 7355 54723 7361
rect 54754 7352 54760 7404
rect 54812 7352 54818 7404
rect 77662 7352 77668 7404
rect 77720 7392 77726 7404
rect 77757 7395 77815 7401
rect 77757 7392 77769 7395
rect 77720 7364 77769 7392
rect 77720 7352 77726 7364
rect 77757 7361 77769 7364
rect 77803 7361 77815 7395
rect 78033 7395 78091 7401
rect 78033 7392 78045 7395
rect 77757 7355 77815 7361
rect 77956 7364 78045 7392
rect 43640 7296 44220 7324
rect 51997 7327 52055 7333
rect 51997 7293 52009 7327
rect 52043 7324 52055 7327
rect 52733 7327 52791 7333
rect 52733 7324 52745 7327
rect 52043 7296 52745 7324
rect 52043 7293 52055 7296
rect 51997 7287 52055 7293
rect 52733 7293 52745 7296
rect 52779 7293 52791 7327
rect 53760 7324 53788 7352
rect 55033 7327 55091 7333
rect 55033 7324 55045 7327
rect 52733 7287 52791 7293
rect 53300 7296 53788 7324
rect 53852 7296 55045 7324
rect 45738 7256 45744 7268
rect 43548 7228 45744 7256
rect 45738 7216 45744 7228
rect 45796 7216 45802 7268
rect 50522 7216 50528 7268
rect 50580 7256 50586 7268
rect 53300 7256 53328 7296
rect 50580 7228 53328 7256
rect 50580 7216 50586 7228
rect 53374 7216 53380 7268
rect 53432 7256 53438 7268
rect 53852 7256 53880 7296
rect 55033 7293 55045 7296
rect 55079 7293 55091 7327
rect 56781 7327 56839 7333
rect 56781 7324 56793 7327
rect 55033 7287 55091 7293
rect 55140 7296 56793 7324
rect 53432 7228 53880 7256
rect 53432 7216 53438 7228
rect 54202 7216 54208 7268
rect 54260 7256 54266 7268
rect 55140 7256 55168 7296
rect 56781 7293 56793 7296
rect 56827 7293 56839 7327
rect 56781 7287 56839 7293
rect 77956 7265 77984 7364
rect 78033 7361 78045 7364
rect 78079 7361 78091 7395
rect 78033 7355 78091 7361
rect 54260 7228 55168 7256
rect 77941 7259 77999 7265
rect 54260 7216 54266 7228
rect 77941 7225 77953 7259
rect 77987 7225 77999 7259
rect 77941 7219 77999 7225
rect 44818 7188 44824 7200
rect 43456 7160 44824 7188
rect 44818 7148 44824 7160
rect 44876 7148 44882 7200
rect 49694 7148 49700 7200
rect 49752 7148 49758 7200
rect 51905 7191 51963 7197
rect 51905 7157 51917 7191
rect 51951 7188 51963 7191
rect 52546 7188 52552 7200
rect 51951 7160 52552 7188
rect 51951 7157 51963 7160
rect 51905 7151 51963 7157
rect 52546 7148 52552 7160
rect 52604 7188 52610 7200
rect 53558 7188 53564 7200
rect 52604 7160 53564 7188
rect 52604 7148 52610 7160
rect 53558 7148 53564 7160
rect 53616 7188 53622 7200
rect 54481 7191 54539 7197
rect 54481 7188 54493 7191
rect 53616 7160 54493 7188
rect 53616 7148 53622 7160
rect 54481 7157 54493 7160
rect 54527 7157 54539 7191
rect 54481 7151 54539 7157
rect 55766 7148 55772 7200
rect 55824 7188 55830 7200
rect 56873 7191 56931 7197
rect 56873 7188 56885 7191
rect 55824 7160 56885 7188
rect 55824 7148 55830 7160
rect 56873 7157 56885 7160
rect 56919 7157 56931 7191
rect 56873 7151 56931 7157
rect 77662 7148 77668 7200
rect 77720 7148 77726 7200
rect 78214 7148 78220 7200
rect 78272 7148 78278 7200
rect 1104 7098 78844 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 78844 7098
rect 1104 7024 78844 7046
rect 30088 6987 30146 6993
rect 30088 6953 30100 6987
rect 30134 6984 30146 6987
rect 30742 6984 30748 6996
rect 30134 6956 30748 6984
rect 30134 6953 30146 6956
rect 30088 6947 30146 6953
rect 30742 6944 30748 6956
rect 30800 6944 30806 6996
rect 31754 6944 31760 6996
rect 31812 6984 31818 6996
rect 32217 6987 32275 6993
rect 32217 6984 32229 6987
rect 31812 6956 32229 6984
rect 31812 6944 31818 6956
rect 32217 6953 32229 6956
rect 32263 6984 32275 6987
rect 33410 6984 33416 6996
rect 32263 6956 33416 6984
rect 32263 6953 32275 6956
rect 32217 6947 32275 6953
rect 33410 6944 33416 6956
rect 33468 6944 33474 6996
rect 34054 6944 34060 6996
rect 34112 6993 34118 6996
rect 34112 6987 34127 6993
rect 34115 6953 34127 6987
rect 34112 6947 34127 6953
rect 34112 6944 34118 6947
rect 44266 6944 44272 6996
rect 44324 6984 44330 6996
rect 46198 6984 46204 6996
rect 44324 6956 46204 6984
rect 44324 6944 44330 6956
rect 46198 6944 46204 6956
rect 46256 6944 46262 6996
rect 46290 6944 46296 6996
rect 46348 6984 46354 6996
rect 46842 6984 46848 6996
rect 46348 6956 46848 6984
rect 46348 6944 46354 6956
rect 46842 6944 46848 6956
rect 46900 6984 46906 6996
rect 47213 6987 47271 6993
rect 47213 6984 47225 6987
rect 46900 6956 47225 6984
rect 46900 6944 46906 6956
rect 47213 6953 47225 6956
rect 47259 6953 47271 6987
rect 47213 6947 47271 6953
rect 50798 6944 50804 6996
rect 50856 6984 50862 6996
rect 53285 6987 53343 6993
rect 53285 6984 53297 6987
rect 50856 6956 53297 6984
rect 50856 6944 50862 6956
rect 53285 6953 53297 6956
rect 53331 6984 53343 6987
rect 54110 6984 54116 6996
rect 53331 6956 54116 6984
rect 53331 6953 53343 6956
rect 53285 6947 53343 6953
rect 54110 6944 54116 6956
rect 54168 6944 54174 6996
rect 37366 6916 37372 6928
rect 37108 6888 37372 6916
rect 29454 6808 29460 6860
rect 29512 6848 29518 6860
rect 29825 6851 29883 6857
rect 29825 6848 29837 6851
rect 29512 6820 29837 6848
rect 29512 6808 29518 6820
rect 29825 6817 29837 6820
rect 29871 6817 29883 6851
rect 29825 6811 29883 6817
rect 31386 6808 31392 6860
rect 31444 6848 31450 6860
rect 31573 6851 31631 6857
rect 31573 6848 31585 6851
rect 31444 6820 31585 6848
rect 31444 6808 31450 6820
rect 31573 6817 31585 6820
rect 31619 6817 31631 6851
rect 31573 6811 31631 6817
rect 32493 6851 32551 6857
rect 32493 6817 32505 6851
rect 32539 6848 32551 6851
rect 33318 6848 33324 6860
rect 32539 6820 33324 6848
rect 32539 6817 32551 6820
rect 32493 6811 32551 6817
rect 31662 6740 31668 6792
rect 31720 6740 31726 6792
rect 31846 6740 31852 6792
rect 31904 6740 31910 6792
rect 32033 6783 32091 6789
rect 32033 6749 32045 6783
rect 32079 6780 32091 6783
rect 32508 6780 32536 6811
rect 33318 6808 33324 6820
rect 33376 6808 33382 6860
rect 33686 6808 33692 6860
rect 33744 6848 33750 6860
rect 35437 6851 35495 6857
rect 35437 6848 35449 6851
rect 33744 6820 35449 6848
rect 33744 6808 33750 6820
rect 35437 6817 35449 6820
rect 35483 6817 35495 6851
rect 37108 6848 37136 6888
rect 37366 6876 37372 6888
rect 37424 6876 37430 6928
rect 38286 6876 38292 6928
rect 38344 6916 38350 6928
rect 41049 6919 41107 6925
rect 38344 6888 39804 6916
rect 38344 6876 38350 6888
rect 35437 6811 35495 6817
rect 36556 6820 37136 6848
rect 32079 6752 32536 6780
rect 34333 6783 34391 6789
rect 32079 6749 32091 6752
rect 32033 6743 32091 6749
rect 34333 6749 34345 6783
rect 34379 6780 34391 6783
rect 34790 6780 34796 6792
rect 34379 6752 34796 6780
rect 34379 6749 34391 6752
rect 34333 6743 34391 6749
rect 31864 6712 31892 6740
rect 31326 6684 31892 6712
rect 31849 6647 31907 6653
rect 31849 6613 31861 6647
rect 31895 6644 31907 6647
rect 32048 6644 32076 6743
rect 34790 6740 34796 6752
rect 34848 6740 34854 6792
rect 35253 6783 35311 6789
rect 35253 6749 35265 6783
rect 35299 6780 35311 6783
rect 35342 6780 35348 6792
rect 35299 6752 35348 6780
rect 35299 6749 35311 6752
rect 35253 6743 35311 6749
rect 35342 6740 35348 6752
rect 35400 6740 35406 6792
rect 35529 6783 35587 6789
rect 35529 6749 35541 6783
rect 35575 6780 35587 6783
rect 36081 6783 36139 6789
rect 36081 6780 36093 6783
rect 35575 6752 36093 6780
rect 35575 6749 35587 6752
rect 35529 6743 35587 6749
rect 36081 6749 36093 6752
rect 36127 6749 36139 6783
rect 36081 6743 36139 6749
rect 33594 6672 33600 6724
rect 33652 6712 33658 6724
rect 33962 6712 33968 6724
rect 33652 6684 33968 6712
rect 33652 6672 33658 6684
rect 33962 6672 33968 6684
rect 34020 6712 34026 6724
rect 35158 6712 35164 6724
rect 34020 6684 35164 6712
rect 34020 6672 34026 6684
rect 35158 6672 35164 6684
rect 35216 6712 35222 6724
rect 36556 6712 36584 6820
rect 37182 6808 37188 6860
rect 37240 6848 37246 6860
rect 37240 6820 37412 6848
rect 37240 6808 37246 6820
rect 36630 6740 36636 6792
rect 36688 6740 36694 6792
rect 37384 6789 37412 6820
rect 38102 6808 38108 6860
rect 38160 6848 38166 6860
rect 39298 6848 39304 6860
rect 38160 6820 38516 6848
rect 38160 6808 38166 6820
rect 37001 6783 37059 6789
rect 37001 6749 37013 6783
rect 37047 6780 37059 6783
rect 37369 6783 37427 6789
rect 37047 6752 37320 6780
rect 37047 6749 37059 6752
rect 37001 6743 37059 6749
rect 35216 6684 36584 6712
rect 36648 6712 36676 6740
rect 37093 6715 37151 6721
rect 37093 6712 37105 6715
rect 36648 6684 37105 6712
rect 35216 6672 35222 6684
rect 37093 6681 37105 6684
rect 37139 6681 37151 6715
rect 37093 6675 37151 6681
rect 37185 6715 37243 6721
rect 37185 6681 37197 6715
rect 37231 6681 37243 6715
rect 37292 6712 37320 6752
rect 37369 6749 37381 6783
rect 37415 6749 37427 6783
rect 37369 6743 37427 6749
rect 37458 6740 37464 6792
rect 37516 6780 37522 6792
rect 38286 6789 38292 6792
rect 38284 6780 38292 6789
rect 37516 6752 38292 6780
rect 37516 6740 37522 6752
rect 38284 6743 38292 6752
rect 38286 6740 38292 6743
rect 38344 6740 38350 6792
rect 38488 6789 38516 6820
rect 38672 6820 39304 6848
rect 38672 6789 38700 6820
rect 39298 6808 39304 6820
rect 39356 6808 39362 6860
rect 39776 6848 39804 6888
rect 41049 6885 41061 6919
rect 41095 6916 41107 6919
rect 41138 6916 41144 6928
rect 41095 6888 41144 6916
rect 41095 6885 41107 6888
rect 41049 6879 41107 6885
rect 41138 6876 41144 6888
rect 41196 6876 41202 6928
rect 44634 6876 44640 6928
rect 44692 6916 44698 6928
rect 45646 6916 45652 6928
rect 44692 6888 45652 6916
rect 44692 6876 44698 6888
rect 45646 6876 45652 6888
rect 45704 6916 45710 6928
rect 45704 6888 47164 6916
rect 45704 6876 45710 6888
rect 39776 6820 40908 6848
rect 38473 6783 38531 6789
rect 38473 6749 38485 6783
rect 38519 6749 38531 6783
rect 38473 6743 38531 6749
rect 38656 6783 38714 6789
rect 38656 6749 38668 6783
rect 38702 6749 38714 6783
rect 38656 6743 38714 6749
rect 37553 6715 37611 6721
rect 37553 6712 37565 6715
rect 37292 6684 37565 6712
rect 37185 6675 37243 6681
rect 37553 6681 37565 6684
rect 37599 6712 37611 6715
rect 37599 6684 38332 6712
rect 37599 6681 37611 6684
rect 37553 6675 37611 6681
rect 31895 6616 32076 6644
rect 32585 6647 32643 6653
rect 31895 6613 31907 6616
rect 31849 6607 31907 6613
rect 32585 6613 32597 6647
rect 32631 6644 32643 6647
rect 33042 6644 33048 6656
rect 32631 6616 33048 6644
rect 32631 6613 32643 6616
rect 32585 6607 32643 6613
rect 33042 6604 33048 6616
rect 33100 6604 33106 6656
rect 33318 6604 33324 6656
rect 33376 6644 33382 6656
rect 34238 6644 34244 6656
rect 33376 6616 34244 6644
rect 33376 6604 33382 6616
rect 34238 6604 34244 6616
rect 34296 6604 34302 6656
rect 35066 6604 35072 6656
rect 35124 6604 35130 6656
rect 35986 6604 35992 6656
rect 36044 6644 36050 6656
rect 36817 6647 36875 6653
rect 36817 6644 36829 6647
rect 36044 6616 36829 6644
rect 36044 6604 36050 6616
rect 36817 6613 36829 6616
rect 36863 6613 36875 6647
rect 36817 6607 36875 6613
rect 36906 6604 36912 6656
rect 36964 6644 36970 6656
rect 37200 6644 37228 6675
rect 37645 6647 37703 6653
rect 37645 6644 37657 6647
rect 36964 6616 37657 6644
rect 36964 6604 36970 6616
rect 37645 6613 37657 6616
rect 37691 6613 37703 6647
rect 37645 6607 37703 6613
rect 38102 6604 38108 6656
rect 38160 6604 38166 6656
rect 38304 6644 38332 6684
rect 38378 6672 38384 6724
rect 38436 6672 38442 6724
rect 38488 6712 38516 6743
rect 38746 6740 38752 6792
rect 38804 6740 38810 6792
rect 40494 6740 40500 6792
rect 40552 6740 40558 6792
rect 40880 6789 40908 6820
rect 41506 6808 41512 6860
rect 41564 6848 41570 6860
rect 41969 6851 42027 6857
rect 41969 6848 41981 6851
rect 41564 6820 41981 6848
rect 41564 6808 41570 6820
rect 41969 6817 41981 6820
rect 42015 6817 42027 6851
rect 42426 6848 42432 6860
rect 41969 6811 42027 6817
rect 42260 6820 42432 6848
rect 40865 6783 40923 6789
rect 40865 6749 40877 6783
rect 40911 6749 40923 6783
rect 40865 6743 40923 6749
rect 40954 6740 40960 6792
rect 41012 6780 41018 6792
rect 42260 6789 42288 6820
rect 42426 6808 42432 6820
rect 42484 6848 42490 6860
rect 42521 6851 42579 6857
rect 42521 6848 42533 6851
rect 42484 6820 42533 6848
rect 42484 6808 42490 6820
rect 42521 6817 42533 6820
rect 42567 6817 42579 6851
rect 42521 6811 42579 6817
rect 43346 6808 43352 6860
rect 43404 6848 43410 6860
rect 44729 6851 44787 6857
rect 44729 6848 44741 6851
rect 43404 6820 44741 6848
rect 43404 6808 43410 6820
rect 44729 6817 44741 6820
rect 44775 6817 44787 6851
rect 44729 6811 44787 6817
rect 45002 6808 45008 6860
rect 45060 6808 45066 6860
rect 45830 6808 45836 6860
rect 45888 6848 45894 6860
rect 46658 6848 46664 6860
rect 45888 6820 46664 6848
rect 45888 6808 45894 6820
rect 46658 6808 46664 6820
rect 46716 6808 46722 6860
rect 41233 6783 41291 6789
rect 41233 6780 41245 6783
rect 41012 6752 41245 6780
rect 41012 6740 41018 6752
rect 41233 6749 41245 6752
rect 41279 6749 41291 6783
rect 41233 6743 41291 6749
rect 41785 6783 41843 6789
rect 41785 6749 41797 6783
rect 41831 6780 41843 6783
rect 41877 6783 41935 6789
rect 41877 6780 41889 6783
rect 41831 6752 41889 6780
rect 41831 6749 41843 6752
rect 41785 6743 41843 6749
rect 41877 6749 41889 6752
rect 41923 6749 41935 6783
rect 41877 6743 41935 6749
rect 42153 6783 42211 6789
rect 42153 6749 42165 6783
rect 42199 6749 42211 6783
rect 42153 6743 42211 6749
rect 42245 6783 42303 6789
rect 42245 6749 42257 6783
rect 42291 6749 42303 6783
rect 42245 6743 42303 6749
rect 40678 6712 40684 6724
rect 38488 6684 40684 6712
rect 40678 6672 40684 6684
rect 40736 6672 40742 6724
rect 40770 6672 40776 6724
rect 40828 6672 40834 6724
rect 41138 6672 41144 6724
rect 41196 6712 41202 6724
rect 42168 6712 42196 6743
rect 42794 6740 42800 6792
rect 42852 6780 42858 6792
rect 42981 6783 43039 6789
rect 42981 6780 42993 6783
rect 42852 6752 42993 6780
rect 42852 6740 42858 6752
rect 42981 6749 42993 6752
rect 43027 6749 43039 6783
rect 42981 6743 43039 6749
rect 46198 6740 46204 6792
rect 46256 6780 46262 6792
rect 46385 6783 46443 6789
rect 46385 6780 46397 6783
rect 46256 6752 46397 6780
rect 46256 6740 46262 6752
rect 46385 6749 46397 6752
rect 46431 6749 46443 6783
rect 46385 6743 46443 6749
rect 46474 6740 46480 6792
rect 46532 6740 46538 6792
rect 47136 6789 47164 6888
rect 49878 6876 49884 6928
rect 49936 6916 49942 6928
rect 49936 6888 51074 6916
rect 49936 6876 49942 6888
rect 51046 6860 51074 6888
rect 49786 6808 49792 6860
rect 49844 6808 49850 6860
rect 50982 6808 50988 6860
rect 51040 6848 51074 6860
rect 51626 6848 51632 6860
rect 51040 6820 51632 6848
rect 51040 6808 51046 6820
rect 51626 6808 51632 6820
rect 51684 6808 51690 6860
rect 46850 6783 46908 6789
rect 46850 6749 46862 6783
rect 46896 6749 46908 6783
rect 46850 6743 46908 6749
rect 47121 6783 47179 6789
rect 47121 6749 47133 6783
rect 47167 6780 47179 6783
rect 47302 6780 47308 6792
rect 47167 6752 47308 6780
rect 47167 6749 47179 6752
rect 47121 6743 47179 6749
rect 41196 6684 42196 6712
rect 41196 6672 41202 6684
rect 43254 6672 43260 6724
rect 43312 6672 43318 6724
rect 44266 6672 44272 6724
rect 44324 6672 44330 6724
rect 45554 6672 45560 6724
rect 45612 6712 45618 6724
rect 45738 6712 45744 6724
rect 45612 6684 45744 6712
rect 45612 6672 45618 6684
rect 45738 6672 45744 6684
rect 45796 6712 45802 6724
rect 45796 6684 46612 6712
rect 45796 6672 45802 6684
rect 41506 6644 41512 6656
rect 38304 6616 41512 6644
rect 41506 6604 41512 6616
rect 41564 6604 41570 6656
rect 41598 6604 41604 6656
rect 41656 6644 41662 6656
rect 42429 6647 42487 6653
rect 42429 6644 42441 6647
rect 41656 6616 42441 6644
rect 41656 6604 41662 6616
rect 42429 6613 42441 6616
rect 42475 6613 42487 6647
rect 42429 6607 42487 6613
rect 44910 6604 44916 6656
rect 44968 6644 44974 6656
rect 45830 6644 45836 6656
rect 44968 6616 45836 6644
rect 44968 6604 44974 6616
rect 45830 6604 45836 6616
rect 45888 6604 45894 6656
rect 46584 6644 46612 6684
rect 46658 6672 46664 6724
rect 46716 6672 46722 6724
rect 46750 6672 46756 6724
rect 46808 6672 46814 6724
rect 46860 6644 46888 6743
rect 47302 6740 47308 6752
rect 47360 6740 47366 6792
rect 47397 6783 47455 6789
rect 47397 6749 47409 6783
rect 47443 6749 47455 6783
rect 47397 6743 47455 6749
rect 49513 6783 49571 6789
rect 49513 6749 49525 6783
rect 49559 6749 49571 6783
rect 49513 6743 49571 6749
rect 49605 6783 49663 6789
rect 49605 6749 49617 6783
rect 49651 6780 49663 6783
rect 49694 6780 49700 6792
rect 49651 6752 49700 6780
rect 49651 6749 49663 6752
rect 49605 6743 49663 6749
rect 47412 6712 47440 6743
rect 47044 6684 47440 6712
rect 49528 6712 49556 6743
rect 49694 6740 49700 6752
rect 49752 6740 49758 6792
rect 49881 6783 49939 6789
rect 49881 6749 49893 6783
rect 49927 6780 49939 6783
rect 50430 6780 50436 6792
rect 49927 6752 50436 6780
rect 49927 6749 49939 6752
rect 49881 6743 49939 6749
rect 50430 6740 50436 6752
rect 50488 6740 50494 6792
rect 77757 6783 77815 6789
rect 77757 6749 77769 6783
rect 77803 6780 77815 6783
rect 77846 6780 77852 6792
rect 77803 6752 77852 6780
rect 77803 6749 77815 6752
rect 77757 6743 77815 6749
rect 77846 6740 77852 6752
rect 77904 6740 77910 6792
rect 51902 6712 51908 6724
rect 49528 6684 51908 6712
rect 47044 6653 47072 6684
rect 51902 6672 51908 6684
rect 51960 6672 51966 6724
rect 46584 6616 46888 6644
rect 47029 6647 47087 6653
rect 47029 6613 47041 6647
rect 47075 6613 47087 6647
rect 47029 6607 47087 6613
rect 47581 6647 47639 6653
rect 47581 6613 47593 6647
rect 47627 6644 47639 6647
rect 49050 6644 49056 6656
rect 47627 6616 49056 6644
rect 47627 6613 47639 6616
rect 47581 6607 47639 6613
rect 49050 6604 49056 6616
rect 49108 6604 49114 6656
rect 49329 6647 49387 6653
rect 49329 6613 49341 6647
rect 49375 6644 49387 6647
rect 49694 6644 49700 6656
rect 49375 6616 49700 6644
rect 49375 6613 49387 6616
rect 49329 6607 49387 6613
rect 49694 6604 49700 6616
rect 49752 6604 49758 6656
rect 78030 6604 78036 6656
rect 78088 6604 78094 6656
rect 1104 6554 78844 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 66314 6554
rect 66366 6502 66378 6554
rect 66430 6502 66442 6554
rect 66494 6502 66506 6554
rect 66558 6502 66570 6554
rect 66622 6502 78844 6554
rect 1104 6480 78844 6502
rect 30098 6400 30104 6452
rect 30156 6400 30162 6452
rect 31478 6400 31484 6452
rect 31536 6440 31542 6452
rect 33502 6440 33508 6452
rect 31536 6412 33508 6440
rect 31536 6400 31542 6412
rect 33502 6400 33508 6412
rect 33560 6400 33566 6452
rect 33689 6443 33747 6449
rect 33689 6409 33701 6443
rect 33735 6440 33747 6443
rect 33870 6440 33876 6452
rect 33735 6412 33876 6440
rect 33735 6409 33747 6412
rect 33689 6403 33747 6409
rect 33870 6400 33876 6412
rect 33928 6400 33934 6452
rect 36541 6443 36599 6449
rect 36541 6440 36553 6443
rect 34992 6412 36553 6440
rect 30116 6372 30144 6400
rect 30285 6375 30343 6381
rect 30285 6372 30297 6375
rect 30116 6344 30297 6372
rect 30285 6341 30297 6344
rect 30331 6341 30343 6375
rect 30285 6335 30343 6341
rect 31386 6332 31392 6384
rect 31444 6372 31450 6384
rect 31573 6375 31631 6381
rect 31573 6372 31585 6375
rect 31444 6344 31585 6372
rect 31444 6332 31450 6344
rect 31573 6341 31585 6344
rect 31619 6341 31631 6375
rect 31573 6335 31631 6341
rect 31665 6375 31723 6381
rect 31665 6341 31677 6375
rect 31711 6372 31723 6375
rect 31754 6372 31760 6384
rect 31711 6344 31760 6372
rect 31711 6341 31723 6344
rect 31665 6335 31723 6341
rect 31754 6332 31760 6344
rect 31812 6332 31818 6384
rect 33413 6375 33471 6381
rect 33413 6372 33425 6375
rect 31864 6344 33425 6372
rect 31478 6264 31484 6316
rect 31536 6264 31542 6316
rect 31864 6313 31892 6344
rect 33413 6341 33425 6344
rect 33459 6372 33471 6375
rect 34992 6372 35020 6412
rect 36541 6409 36553 6412
rect 36587 6440 36599 6443
rect 36630 6440 36636 6452
rect 36587 6412 36636 6440
rect 36587 6409 36599 6412
rect 36541 6403 36599 6409
rect 36630 6400 36636 6412
rect 36688 6400 36694 6452
rect 40129 6443 40187 6449
rect 40129 6409 40141 6443
rect 40175 6440 40187 6443
rect 40954 6440 40960 6452
rect 40175 6412 40960 6440
rect 40175 6409 40187 6412
rect 40129 6403 40187 6409
rect 40954 6400 40960 6412
rect 41012 6440 41018 6452
rect 41690 6440 41696 6452
rect 41012 6412 41696 6440
rect 41012 6400 41018 6412
rect 41690 6400 41696 6412
rect 41748 6400 41754 6452
rect 42426 6400 42432 6452
rect 42484 6440 42490 6452
rect 42797 6443 42855 6449
rect 42797 6440 42809 6443
rect 42484 6412 42809 6440
rect 42484 6400 42490 6412
rect 42797 6409 42809 6412
rect 42843 6409 42855 6443
rect 42797 6403 42855 6409
rect 42981 6443 43039 6449
rect 42981 6409 42993 6443
rect 43027 6440 43039 6443
rect 43254 6440 43260 6452
rect 43027 6412 43260 6440
rect 43027 6409 43039 6412
rect 42981 6403 43039 6409
rect 33459 6344 35020 6372
rect 33459 6341 33471 6344
rect 33413 6335 33471 6341
rect 35066 6332 35072 6384
rect 35124 6332 35130 6384
rect 35158 6332 35164 6384
rect 35216 6372 35222 6384
rect 38746 6372 38752 6384
rect 35216 6344 35558 6372
rect 36740 6344 38752 6372
rect 35216 6332 35222 6344
rect 31849 6307 31907 6313
rect 31849 6273 31861 6307
rect 31895 6273 31907 6307
rect 31849 6267 31907 6273
rect 32950 6264 32956 6316
rect 33008 6304 33014 6316
rect 33045 6307 33103 6313
rect 33045 6304 33057 6307
rect 33008 6276 33057 6304
rect 33008 6264 33014 6276
rect 33045 6273 33057 6276
rect 33091 6273 33103 6307
rect 33045 6267 33103 6273
rect 33193 6307 33251 6313
rect 33193 6273 33205 6307
rect 33239 6304 33251 6307
rect 33239 6273 33272 6304
rect 33193 6267 33272 6273
rect 29454 6196 29460 6248
rect 29512 6236 29518 6248
rect 31021 6239 31079 6245
rect 31021 6236 31033 6239
rect 29512 6208 31033 6236
rect 29512 6196 29518 6208
rect 31021 6205 31033 6208
rect 31067 6205 31079 6239
rect 33244 6236 33272 6267
rect 33318 6264 33324 6316
rect 33376 6264 33382 6316
rect 33502 6264 33508 6316
rect 33560 6313 33566 6316
rect 33560 6304 33568 6313
rect 33560 6276 33605 6304
rect 33560 6267 33568 6276
rect 33560 6264 33566 6267
rect 34790 6264 34796 6316
rect 34848 6264 34854 6316
rect 36630 6264 36636 6316
rect 36688 6304 36694 6316
rect 36740 6304 36768 6344
rect 38746 6332 38752 6344
rect 38804 6332 38810 6384
rect 41138 6332 41144 6384
rect 41196 6332 41202 6384
rect 41598 6332 41604 6384
rect 41656 6332 41662 6384
rect 36688 6276 36768 6304
rect 36688 6264 36694 6276
rect 38102 6264 38108 6316
rect 38160 6304 38166 6316
rect 38473 6307 38531 6313
rect 38473 6304 38485 6307
rect 38160 6276 38485 6304
rect 38160 6264 38166 6276
rect 38473 6273 38485 6276
rect 38519 6273 38531 6307
rect 42812 6304 42840 6403
rect 43254 6400 43260 6412
rect 43312 6400 43318 6452
rect 44174 6400 44180 6452
rect 44232 6440 44238 6452
rect 44269 6443 44327 6449
rect 44269 6440 44281 6443
rect 44232 6412 44281 6440
rect 44232 6400 44238 6412
rect 44269 6409 44281 6412
rect 44315 6440 44327 6443
rect 44450 6440 44456 6452
rect 44315 6412 44456 6440
rect 44315 6409 44327 6412
rect 44269 6403 44327 6409
rect 44450 6400 44456 6412
rect 44508 6400 44514 6452
rect 44910 6440 44916 6452
rect 44744 6412 44916 6440
rect 43070 6332 43076 6384
rect 43128 6372 43134 6384
rect 44744 6381 44772 6412
rect 44910 6400 44916 6412
rect 44968 6400 44974 6452
rect 45002 6400 45008 6452
rect 45060 6400 45066 6452
rect 45097 6443 45155 6449
rect 45097 6409 45109 6443
rect 45143 6440 45155 6443
rect 45143 6412 46520 6440
rect 45143 6409 45155 6412
rect 45097 6403 45155 6409
rect 44729 6375 44787 6381
rect 43128 6344 43300 6372
rect 43128 6332 43134 6344
rect 43272 6313 43300 6344
rect 44729 6341 44741 6375
rect 44775 6341 44787 6375
rect 44729 6335 44787 6341
rect 44818 6332 44824 6384
rect 44876 6332 44882 6384
rect 45020 6372 45048 6400
rect 45189 6375 45247 6381
rect 45189 6372 45201 6375
rect 45020 6344 45201 6372
rect 45189 6341 45201 6344
rect 45235 6341 45247 6375
rect 45189 6335 45247 6341
rect 43165 6307 43223 6313
rect 43165 6304 43177 6307
rect 42812 6276 43177 6304
rect 38473 6267 38531 6273
rect 43165 6273 43177 6276
rect 43211 6273 43223 6307
rect 43165 6267 43223 6273
rect 43257 6307 43315 6313
rect 43257 6273 43269 6307
rect 43303 6273 43315 6307
rect 43257 6267 43315 6273
rect 43346 6264 43352 6316
rect 43404 6304 43410 6316
rect 43533 6307 43591 6313
rect 43533 6304 43545 6307
rect 43404 6276 43545 6304
rect 43404 6264 43410 6276
rect 43533 6273 43545 6276
rect 43579 6273 43591 6307
rect 43533 6267 43591 6273
rect 44450 6264 44456 6316
rect 44508 6264 44514 6316
rect 44634 6313 44640 6316
rect 44601 6307 44640 6313
rect 44601 6273 44613 6307
rect 44601 6267 44640 6273
rect 44634 6264 44640 6267
rect 44692 6264 44698 6316
rect 44959 6307 45017 6313
rect 44959 6273 44971 6307
rect 45005 6304 45017 6307
rect 45554 6304 45560 6316
rect 45005 6276 45560 6304
rect 45005 6273 45017 6276
rect 44959 6267 45017 6273
rect 45554 6264 45560 6276
rect 45612 6264 45618 6316
rect 46492 6313 46520 6412
rect 47302 6400 47308 6452
rect 47360 6440 47366 6452
rect 47581 6443 47639 6449
rect 47581 6440 47593 6443
rect 47360 6412 47593 6440
rect 47360 6400 47366 6412
rect 47581 6409 47593 6412
rect 47627 6409 47639 6443
rect 47581 6403 47639 6409
rect 47780 6412 49832 6440
rect 47780 6384 47808 6412
rect 46566 6332 46572 6384
rect 46624 6372 46630 6384
rect 47762 6372 47768 6384
rect 46624 6344 47768 6372
rect 46624 6332 46630 6344
rect 47762 6332 47768 6344
rect 47820 6372 47826 6384
rect 47820 6344 47886 6372
rect 47820 6332 47826 6344
rect 49050 6332 49056 6384
rect 49108 6332 49114 6384
rect 49694 6332 49700 6384
rect 49752 6332 49758 6384
rect 49804 6372 49832 6412
rect 50430 6400 50436 6452
rect 50488 6440 50494 6452
rect 51169 6443 51227 6449
rect 51169 6440 51181 6443
rect 50488 6412 51181 6440
rect 50488 6400 50494 6412
rect 51169 6409 51181 6412
rect 51215 6409 51227 6443
rect 51169 6403 51227 6409
rect 54941 6443 54999 6449
rect 54941 6409 54953 6443
rect 54987 6440 54999 6443
rect 55122 6440 55128 6452
rect 54987 6412 55128 6440
rect 54987 6409 54999 6412
rect 54941 6403 54999 6409
rect 55122 6400 55128 6412
rect 55180 6400 55186 6452
rect 49970 6372 49976 6384
rect 49804 6344 49976 6372
rect 49970 6332 49976 6344
rect 50028 6372 50034 6384
rect 50028 6344 50186 6372
rect 50028 6332 50034 6344
rect 46477 6307 46535 6313
rect 46477 6273 46489 6307
rect 46523 6273 46535 6307
rect 46477 6267 46535 6273
rect 51626 6264 51632 6316
rect 51684 6304 51690 6316
rect 53650 6304 53656 6316
rect 51684 6276 53656 6304
rect 51684 6264 51690 6276
rect 53650 6264 53656 6276
rect 53708 6304 53714 6316
rect 53745 6307 53803 6313
rect 53745 6304 53757 6307
rect 53708 6276 53757 6304
rect 53708 6264 53714 6276
rect 53745 6273 53757 6276
rect 53791 6273 53803 6307
rect 53745 6267 53803 6273
rect 53837 6307 53895 6313
rect 53837 6273 53849 6307
rect 53883 6273 53895 6307
rect 53837 6267 53895 6273
rect 53929 6307 53987 6313
rect 53929 6273 53941 6307
rect 53975 6304 53987 6307
rect 54018 6304 54024 6316
rect 53975 6276 54024 6304
rect 53975 6273 53987 6276
rect 53929 6267 53987 6273
rect 34422 6236 34428 6248
rect 33244 6208 34428 6236
rect 31021 6199 31079 6205
rect 34422 6196 34428 6208
rect 34480 6196 34486 6248
rect 31202 6060 31208 6112
rect 31260 6100 31266 6112
rect 31297 6103 31355 6109
rect 31297 6100 31309 6103
rect 31260 6072 31309 6100
rect 31260 6060 31266 6072
rect 31297 6069 31309 6072
rect 31343 6069 31355 6103
rect 31297 6063 31355 6069
rect 32950 6060 32956 6112
rect 33008 6100 33014 6112
rect 34146 6100 34152 6112
rect 33008 6072 34152 6100
rect 33008 6060 33014 6072
rect 34146 6060 34152 6072
rect 34204 6060 34210 6112
rect 34808 6100 34836 6264
rect 36906 6196 36912 6248
rect 36964 6236 36970 6248
rect 38194 6236 38200 6248
rect 36964 6208 38200 6236
rect 36964 6196 36970 6208
rect 38194 6196 38200 6208
rect 38252 6196 38258 6248
rect 38749 6239 38807 6245
rect 38749 6205 38761 6239
rect 38795 6236 38807 6239
rect 39209 6239 39267 6245
rect 39209 6236 39221 6239
rect 38795 6208 39221 6236
rect 38795 6205 38807 6208
rect 38749 6199 38807 6205
rect 39209 6205 39221 6208
rect 39255 6205 39267 6239
rect 39209 6199 39267 6205
rect 39758 6196 39764 6248
rect 39816 6196 39822 6248
rect 41046 6236 41052 6248
rect 40604 6208 41052 6236
rect 37550 6128 37556 6180
rect 37608 6168 37614 6180
rect 38470 6168 38476 6180
rect 37608 6140 38476 6168
rect 37608 6128 37614 6140
rect 38470 6128 38476 6140
rect 38528 6168 38534 6180
rect 38657 6171 38715 6177
rect 38657 6168 38669 6171
rect 38528 6140 38669 6168
rect 38528 6128 38534 6140
rect 38657 6137 38669 6140
rect 38703 6168 38715 6171
rect 40604 6168 40632 6208
rect 41046 6196 41052 6208
rect 41104 6196 41110 6248
rect 41138 6196 41144 6248
rect 41196 6236 41202 6248
rect 41877 6239 41935 6245
rect 41196 6208 41828 6236
rect 41196 6196 41202 6208
rect 38703 6140 40632 6168
rect 41800 6168 41828 6208
rect 41877 6205 41889 6239
rect 41923 6236 41935 6239
rect 42794 6236 42800 6248
rect 41923 6208 42800 6236
rect 41923 6205 41935 6208
rect 41877 6199 41935 6205
rect 42794 6196 42800 6208
rect 42852 6196 42858 6248
rect 45094 6196 45100 6248
rect 45152 6236 45158 6248
rect 45925 6239 45983 6245
rect 45925 6236 45937 6239
rect 45152 6208 45937 6236
rect 45152 6196 45158 6208
rect 45925 6205 45937 6208
rect 45971 6205 45983 6239
rect 45925 6199 45983 6205
rect 42242 6168 42248 6180
rect 41800 6140 42248 6168
rect 38703 6137 38715 6140
rect 38657 6131 38715 6137
rect 42242 6128 42248 6140
rect 42300 6128 42306 6180
rect 45940 6168 45968 6199
rect 46106 6196 46112 6248
rect 46164 6236 46170 6248
rect 46201 6239 46259 6245
rect 46201 6236 46213 6239
rect 46164 6208 46213 6236
rect 46164 6196 46170 6208
rect 46201 6205 46213 6208
rect 46247 6236 46259 6239
rect 46750 6236 46756 6248
rect 46247 6208 46756 6236
rect 46247 6205 46259 6208
rect 46201 6199 46259 6205
rect 46750 6196 46756 6208
rect 46808 6196 46814 6248
rect 48038 6236 48044 6248
rect 46860 6208 48044 6236
rect 46860 6168 46888 6208
rect 48038 6196 48044 6208
rect 48096 6236 48102 6248
rect 49329 6239 49387 6245
rect 49329 6236 49341 6239
rect 48096 6208 49341 6236
rect 48096 6196 48102 6208
rect 49329 6205 49341 6208
rect 49375 6236 49387 6239
rect 49421 6239 49479 6245
rect 49421 6236 49433 6239
rect 49375 6208 49433 6236
rect 49375 6205 49387 6208
rect 49329 6199 49387 6205
rect 49421 6205 49433 6208
rect 49467 6205 49479 6239
rect 49421 6199 49479 6205
rect 50706 6196 50712 6248
rect 50764 6236 50770 6248
rect 53282 6236 53288 6248
rect 50764 6208 53288 6236
rect 50764 6196 50770 6208
rect 53282 6196 53288 6208
rect 53340 6236 53346 6248
rect 53377 6239 53435 6245
rect 53377 6236 53389 6239
rect 53340 6208 53389 6236
rect 53340 6196 53346 6208
rect 53377 6205 53389 6208
rect 53423 6236 53435 6239
rect 53852 6236 53880 6267
rect 54018 6264 54024 6276
rect 54076 6264 54082 6316
rect 54113 6307 54171 6313
rect 54113 6273 54125 6307
rect 54159 6304 54171 6307
rect 54202 6304 54208 6316
rect 54159 6276 54208 6304
rect 54159 6273 54171 6276
rect 54113 6267 54171 6273
rect 54202 6264 54208 6276
rect 54260 6264 54266 6316
rect 54757 6307 54815 6313
rect 54757 6273 54769 6307
rect 54803 6304 54815 6307
rect 54803 6276 55260 6304
rect 54803 6273 54815 6276
rect 54757 6267 54815 6273
rect 53423 6208 53880 6236
rect 53423 6205 53435 6208
rect 53377 6199 53435 6205
rect 45940 6140 46888 6168
rect 46768 6112 46796 6140
rect 36078 6100 36084 6112
rect 34808 6072 36084 6100
rect 36078 6060 36084 6072
rect 36136 6060 36142 6112
rect 38102 6060 38108 6112
rect 38160 6100 38166 6112
rect 38289 6103 38347 6109
rect 38289 6100 38301 6103
rect 38160 6072 38301 6100
rect 38160 6060 38166 6072
rect 38289 6069 38301 6072
rect 38335 6069 38347 6103
rect 38289 6063 38347 6069
rect 41506 6060 41512 6112
rect 41564 6100 41570 6112
rect 42518 6100 42524 6112
rect 41564 6072 42524 6100
rect 41564 6060 41570 6072
rect 42518 6060 42524 6072
rect 42576 6060 42582 6112
rect 43441 6103 43499 6109
rect 43441 6069 43453 6103
rect 43487 6100 43499 6103
rect 43714 6100 43720 6112
rect 43487 6072 43720 6100
rect 43487 6069 43499 6072
rect 43441 6063 43499 6069
rect 43714 6060 43720 6072
rect 43772 6060 43778 6112
rect 46290 6060 46296 6112
rect 46348 6060 46354 6112
rect 46474 6060 46480 6112
rect 46532 6100 46538 6112
rect 46661 6103 46719 6109
rect 46661 6100 46673 6103
rect 46532 6072 46673 6100
rect 46532 6060 46538 6072
rect 46661 6069 46673 6072
rect 46707 6069 46719 6103
rect 46661 6063 46719 6069
rect 46750 6060 46756 6112
rect 46808 6060 46814 6112
rect 49510 6060 49516 6112
rect 49568 6100 49574 6112
rect 52454 6100 52460 6112
rect 49568 6072 52460 6100
rect 49568 6060 49574 6072
rect 52454 6060 52460 6072
rect 52512 6060 52518 6112
rect 52822 6060 52828 6112
rect 52880 6060 52886 6112
rect 53561 6103 53619 6109
rect 53561 6069 53573 6103
rect 53607 6100 53619 6103
rect 53650 6100 53656 6112
rect 53607 6072 53656 6100
rect 53607 6069 53619 6072
rect 53561 6063 53619 6069
rect 53650 6060 53656 6072
rect 53708 6060 53714 6112
rect 53742 6060 53748 6112
rect 53800 6100 53806 6112
rect 55232 6109 55260 6276
rect 78030 6264 78036 6316
rect 78088 6264 78094 6316
rect 78214 6128 78220 6180
rect 78272 6128 78278 6180
rect 54205 6103 54263 6109
rect 54205 6100 54217 6103
rect 53800 6072 54217 6100
rect 53800 6060 53806 6072
rect 54205 6069 54217 6072
rect 54251 6069 54263 6103
rect 54205 6063 54263 6069
rect 55217 6103 55275 6109
rect 55217 6069 55229 6103
rect 55263 6100 55275 6103
rect 55306 6100 55312 6112
rect 55263 6072 55312 6100
rect 55263 6069 55275 6072
rect 55217 6063 55275 6069
rect 55306 6060 55312 6072
rect 55364 6060 55370 6112
rect 1104 6010 78844 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 78844 6010
rect 1104 5936 78844 5958
rect 31846 5856 31852 5908
rect 31904 5896 31910 5908
rect 32217 5899 32275 5905
rect 32217 5896 32229 5899
rect 31904 5868 32229 5896
rect 31904 5856 31910 5868
rect 32217 5865 32229 5868
rect 32263 5865 32275 5899
rect 32217 5859 32275 5865
rect 34238 5856 34244 5908
rect 34296 5896 34302 5908
rect 34296 5868 35204 5896
rect 34296 5856 34302 5868
rect 32030 5788 32036 5840
rect 32088 5828 32094 5840
rect 32125 5831 32183 5837
rect 32125 5828 32137 5831
rect 32088 5800 32137 5828
rect 32088 5788 32094 5800
rect 32125 5797 32137 5800
rect 32171 5828 32183 5831
rect 35176 5828 35204 5868
rect 35342 5856 35348 5908
rect 35400 5856 35406 5908
rect 36814 5856 36820 5908
rect 36872 5896 36878 5908
rect 39577 5899 39635 5905
rect 39577 5896 39589 5899
rect 36872 5868 39589 5896
rect 36872 5856 36878 5868
rect 39577 5865 39589 5868
rect 39623 5896 39635 5899
rect 39758 5896 39764 5908
rect 39623 5868 39764 5896
rect 39623 5865 39635 5868
rect 39577 5859 39635 5865
rect 39758 5856 39764 5868
rect 39816 5856 39822 5908
rect 44358 5856 44364 5908
rect 44416 5896 44422 5908
rect 45005 5899 45063 5905
rect 45005 5896 45017 5899
rect 44416 5868 45017 5896
rect 44416 5856 44422 5868
rect 45005 5865 45017 5868
rect 45051 5896 45063 5899
rect 46106 5896 46112 5908
rect 45051 5868 46112 5896
rect 45051 5865 45063 5868
rect 45005 5859 45063 5865
rect 46106 5856 46112 5868
rect 46164 5856 46170 5908
rect 49881 5899 49939 5905
rect 49881 5865 49893 5899
rect 49927 5896 49939 5899
rect 50062 5896 50068 5908
rect 49927 5868 50068 5896
rect 49927 5865 49939 5868
rect 49881 5859 49939 5865
rect 50062 5856 50068 5868
rect 50120 5856 50126 5908
rect 50338 5856 50344 5908
rect 50396 5896 50402 5908
rect 50982 5896 50988 5908
rect 50396 5868 50988 5896
rect 50396 5856 50402 5868
rect 50982 5856 50988 5868
rect 51040 5856 51046 5908
rect 53282 5856 53288 5908
rect 53340 5856 53346 5908
rect 35986 5828 35992 5840
rect 32171 5800 35112 5828
rect 35176 5800 35992 5828
rect 32171 5797 32183 5800
rect 32125 5791 32183 5797
rect 29454 5720 29460 5772
rect 29512 5760 29518 5772
rect 30282 5760 30288 5772
rect 29512 5732 30288 5760
rect 29512 5720 29518 5732
rect 30282 5720 30288 5732
rect 30340 5760 30346 5772
rect 30377 5763 30435 5769
rect 30377 5760 30389 5763
rect 30340 5732 30389 5760
rect 30340 5720 30346 5732
rect 30377 5729 30389 5732
rect 30423 5729 30435 5763
rect 30377 5723 30435 5729
rect 33042 5720 33048 5772
rect 33100 5760 33106 5772
rect 33100 5732 34836 5760
rect 33100 5720 33106 5732
rect 31754 5652 31760 5704
rect 31812 5652 31818 5704
rect 33502 5652 33508 5704
rect 33560 5692 33566 5704
rect 33796 5701 33824 5732
rect 34808 5704 34836 5732
rect 33643 5695 33701 5701
rect 33643 5692 33655 5695
rect 33560 5664 33655 5692
rect 33560 5652 33566 5664
rect 33643 5661 33655 5664
rect 33689 5661 33701 5695
rect 33643 5655 33701 5661
rect 33781 5695 33839 5701
rect 33781 5661 33793 5695
rect 33827 5661 33839 5695
rect 34054 5692 34060 5704
rect 34015 5664 34060 5692
rect 33781 5655 33839 5661
rect 34054 5652 34060 5664
rect 34112 5652 34118 5704
rect 34146 5652 34152 5704
rect 34204 5692 34210 5704
rect 34606 5692 34612 5704
rect 34204 5664 34612 5692
rect 34204 5652 34210 5664
rect 34606 5652 34612 5664
rect 34664 5692 34670 5704
rect 34701 5695 34759 5701
rect 34701 5692 34713 5695
rect 34664 5664 34713 5692
rect 34664 5652 34670 5664
rect 34701 5661 34713 5664
rect 34747 5661 34759 5695
rect 34701 5655 34759 5661
rect 34790 5652 34796 5704
rect 34848 5692 34854 5704
rect 34848 5664 34893 5692
rect 34848 5652 34854 5664
rect 30650 5584 30656 5636
rect 30708 5584 30714 5636
rect 33318 5584 33324 5636
rect 33376 5624 33382 5636
rect 33873 5627 33931 5633
rect 33873 5624 33885 5627
rect 33376 5596 33885 5624
rect 33376 5584 33382 5596
rect 33873 5593 33885 5596
rect 33919 5624 33931 5627
rect 34514 5624 34520 5636
rect 33919 5596 34520 5624
rect 33919 5593 33931 5596
rect 33873 5587 33931 5593
rect 34514 5584 34520 5596
rect 34572 5584 34578 5636
rect 34882 5584 34888 5636
rect 34940 5624 34946 5636
rect 35084 5633 35112 5800
rect 35986 5788 35992 5800
rect 36044 5788 36050 5840
rect 36170 5788 36176 5840
rect 36228 5828 36234 5840
rect 37458 5828 37464 5840
rect 36228 5800 37464 5828
rect 36228 5788 36234 5800
rect 37458 5788 37464 5800
rect 37516 5788 37522 5840
rect 41414 5788 41420 5840
rect 41472 5828 41478 5840
rect 51442 5828 51448 5840
rect 41472 5800 42104 5828
rect 41472 5788 41478 5800
rect 36078 5720 36084 5772
rect 36136 5760 36142 5772
rect 37829 5763 37887 5769
rect 37829 5760 37841 5763
rect 36136 5732 37841 5760
rect 36136 5720 36142 5732
rect 37829 5729 37841 5732
rect 37875 5729 37887 5763
rect 37829 5723 37887 5729
rect 38102 5720 38108 5772
rect 38160 5720 38166 5772
rect 41386 5732 41828 5760
rect 35158 5652 35164 5704
rect 35216 5701 35222 5704
rect 35216 5692 35224 5701
rect 35216 5664 35261 5692
rect 35216 5655 35224 5664
rect 35216 5652 35222 5655
rect 36630 5652 36636 5704
rect 36688 5652 36694 5704
rect 36814 5701 36820 5704
rect 36781 5695 36820 5701
rect 36781 5661 36793 5695
rect 36781 5655 36820 5661
rect 36814 5652 36820 5655
rect 36872 5652 36878 5704
rect 36906 5652 36912 5704
rect 36964 5652 36970 5704
rect 37139 5695 37197 5701
rect 37139 5661 37151 5695
rect 37185 5692 37197 5695
rect 37458 5692 37464 5704
rect 37185 5664 37464 5692
rect 37185 5661 37197 5664
rect 37139 5655 37197 5661
rect 37458 5652 37464 5664
rect 37516 5652 37522 5704
rect 40678 5652 40684 5704
rect 40736 5692 40742 5704
rect 41386 5692 41414 5732
rect 40736 5664 41414 5692
rect 41596 5695 41654 5701
rect 40736 5652 40742 5664
rect 41596 5661 41608 5695
rect 41642 5661 41654 5695
rect 41596 5655 41654 5661
rect 34977 5627 35035 5633
rect 34977 5624 34989 5627
rect 34940 5596 34989 5624
rect 34940 5584 34946 5596
rect 34977 5593 34989 5596
rect 35023 5593 35035 5627
rect 34977 5587 35035 5593
rect 35069 5627 35127 5633
rect 35069 5593 35081 5627
rect 35115 5624 35127 5627
rect 35434 5624 35440 5636
rect 35115 5596 35440 5624
rect 35115 5593 35127 5596
rect 35069 5587 35127 5593
rect 35434 5584 35440 5596
rect 35492 5584 35498 5636
rect 33134 5516 33140 5568
rect 33192 5556 33198 5568
rect 33505 5559 33563 5565
rect 33505 5556 33517 5559
rect 33192 5528 33517 5556
rect 33192 5516 33198 5528
rect 33505 5525 33517 5528
rect 33551 5525 33563 5559
rect 33505 5519 33563 5525
rect 34606 5516 34612 5568
rect 34664 5556 34670 5568
rect 36648 5556 36676 5652
rect 37001 5627 37059 5633
rect 37001 5593 37013 5627
rect 37047 5624 37059 5627
rect 37047 5596 37228 5624
rect 37047 5593 37059 5596
rect 37001 5587 37059 5593
rect 37200 5568 37228 5596
rect 37366 5584 37372 5636
rect 37424 5624 37430 5636
rect 41230 5624 41236 5636
rect 37424 5596 37596 5624
rect 39330 5596 41236 5624
rect 37424 5584 37430 5596
rect 34664 5528 36676 5556
rect 34664 5516 34670 5528
rect 37182 5516 37188 5568
rect 37240 5516 37246 5568
rect 37277 5559 37335 5565
rect 37277 5525 37289 5559
rect 37323 5556 37335 5559
rect 37458 5556 37464 5568
rect 37323 5528 37464 5556
rect 37323 5525 37335 5528
rect 37277 5519 37335 5525
rect 37458 5516 37464 5528
rect 37516 5516 37522 5568
rect 37568 5556 37596 5596
rect 41230 5584 41236 5596
rect 41288 5584 41294 5636
rect 41616 5624 41644 5655
rect 41690 5652 41696 5704
rect 41748 5652 41754 5704
rect 41800 5701 41828 5732
rect 41785 5695 41843 5701
rect 41785 5661 41797 5695
rect 41831 5661 41843 5695
rect 41785 5655 41843 5661
rect 41874 5652 41880 5704
rect 41932 5701 41938 5704
rect 42076 5701 42104 5800
rect 50984 5800 51448 5828
rect 46474 5720 46480 5772
rect 46532 5720 46538 5772
rect 46750 5720 46756 5772
rect 46808 5720 46814 5772
rect 50984 5760 51012 5800
rect 51442 5788 51448 5800
rect 51500 5788 51506 5840
rect 78033 5831 78091 5837
rect 78033 5797 78045 5831
rect 78079 5797 78091 5831
rect 78033 5791 78091 5797
rect 49344 5732 50844 5760
rect 41932 5695 41971 5701
rect 41959 5661 41971 5695
rect 41932 5655 41971 5661
rect 42061 5695 42119 5701
rect 42061 5661 42073 5695
rect 42107 5661 42119 5695
rect 42061 5655 42119 5661
rect 41932 5652 41938 5655
rect 46566 5624 46572 5636
rect 41616 5596 41828 5624
rect 46046 5596 46572 5624
rect 41800 5568 41828 5596
rect 46566 5584 46572 5596
rect 46624 5584 46630 5636
rect 41138 5556 41144 5568
rect 37568 5528 41144 5556
rect 41138 5516 41144 5528
rect 41196 5516 41202 5568
rect 41414 5516 41420 5568
rect 41472 5516 41478 5568
rect 41782 5516 41788 5568
rect 41840 5516 41846 5568
rect 46198 5516 46204 5568
rect 46256 5556 46262 5568
rect 49344 5565 49372 5732
rect 50816 5704 50844 5732
rect 50908 5732 51012 5760
rect 50338 5701 50344 5704
rect 49697 5695 49755 5701
rect 49697 5692 49709 5695
rect 49528 5664 49709 5692
rect 49528 5568 49556 5664
rect 49697 5661 49709 5664
rect 49743 5661 49755 5695
rect 50336 5692 50344 5701
rect 50299 5664 50344 5692
rect 49697 5655 49755 5661
rect 50336 5655 50344 5664
rect 50338 5652 50344 5655
rect 50396 5652 50402 5704
rect 50430 5652 50436 5704
rect 50488 5652 50494 5704
rect 50706 5692 50712 5704
rect 50667 5664 50712 5692
rect 50706 5652 50712 5664
rect 50764 5652 50770 5704
rect 50798 5652 50804 5704
rect 50856 5652 50862 5704
rect 50908 5701 50936 5732
rect 51074 5720 51080 5772
rect 51132 5760 51138 5772
rect 54018 5760 54024 5772
rect 51132 5732 51304 5760
rect 51132 5720 51138 5732
rect 50908 5695 50971 5701
rect 50908 5664 50925 5695
rect 50913 5661 50925 5664
rect 50959 5661 50971 5695
rect 50913 5655 50971 5661
rect 51166 5652 51172 5704
rect 51224 5652 51230 5704
rect 51276 5701 51304 5732
rect 51460 5732 54024 5760
rect 51261 5695 51319 5701
rect 51261 5661 51273 5695
rect 51307 5661 51319 5695
rect 51261 5655 51319 5661
rect 50062 5584 50068 5636
rect 50120 5624 50126 5636
rect 50525 5627 50583 5633
rect 50120 5596 50384 5624
rect 50120 5584 50126 5596
rect 49329 5559 49387 5565
rect 49329 5556 49341 5559
rect 46256 5528 49341 5556
rect 46256 5516 46262 5528
rect 49329 5525 49341 5528
rect 49375 5525 49387 5559
rect 49329 5519 49387 5525
rect 49510 5516 49516 5568
rect 49568 5516 49574 5568
rect 49694 5516 49700 5568
rect 49752 5556 49758 5568
rect 50157 5559 50215 5565
rect 50157 5556 50169 5559
rect 49752 5528 50169 5556
rect 49752 5516 49758 5528
rect 50157 5525 50169 5528
rect 50203 5525 50215 5559
rect 50356 5556 50384 5596
rect 50525 5593 50537 5627
rect 50571 5624 50583 5627
rect 51077 5627 51135 5633
rect 51077 5624 51089 5627
rect 50571 5596 51089 5624
rect 50571 5593 50583 5596
rect 50525 5587 50583 5593
rect 51077 5593 51089 5596
rect 51123 5624 51135 5627
rect 51460 5624 51488 5732
rect 54018 5720 54024 5732
rect 54076 5720 54082 5772
rect 55030 5720 55036 5772
rect 55088 5760 55094 5772
rect 55125 5763 55183 5769
rect 55125 5760 55137 5763
rect 55088 5732 55137 5760
rect 55088 5720 55094 5732
rect 55125 5729 55137 5732
rect 55171 5760 55183 5763
rect 55582 5760 55588 5772
rect 55171 5732 55588 5760
rect 55171 5729 55183 5732
rect 55125 5723 55183 5729
rect 55582 5720 55588 5732
rect 55640 5720 55646 5772
rect 51537 5695 51595 5701
rect 51537 5661 51549 5695
rect 51583 5661 51595 5695
rect 51537 5655 51595 5661
rect 51123 5596 51488 5624
rect 51123 5593 51135 5596
rect 51077 5587 51135 5593
rect 50540 5556 50568 5587
rect 50356 5528 50568 5556
rect 50157 5519 50215 5525
rect 51442 5516 51448 5568
rect 51500 5516 51506 5568
rect 51552 5556 51580 5655
rect 52914 5652 52920 5704
rect 52972 5652 52978 5704
rect 53374 5652 53380 5704
rect 53432 5652 53438 5704
rect 77849 5695 77907 5701
rect 77849 5692 77861 5695
rect 77680 5664 77861 5692
rect 51718 5584 51724 5636
rect 51776 5624 51782 5636
rect 51813 5627 51871 5633
rect 51813 5624 51825 5627
rect 51776 5596 51825 5624
rect 51776 5584 51782 5596
rect 51813 5593 51825 5596
rect 51859 5593 51871 5627
rect 51813 5587 51871 5593
rect 52086 5556 52092 5568
rect 51552 5528 52092 5556
rect 52086 5516 52092 5528
rect 52144 5516 52150 5568
rect 52932 5556 52960 5652
rect 53558 5584 53564 5636
rect 53616 5624 53622 5636
rect 53653 5627 53711 5633
rect 53653 5624 53665 5627
rect 53616 5596 53665 5624
rect 53616 5584 53622 5596
rect 53653 5593 53665 5596
rect 53699 5593 53711 5627
rect 53653 5587 53711 5593
rect 54036 5596 54142 5624
rect 53742 5556 53748 5568
rect 52932 5528 53748 5556
rect 53742 5516 53748 5528
rect 53800 5556 53806 5568
rect 54036 5556 54064 5596
rect 55398 5584 55404 5636
rect 55456 5624 55462 5636
rect 55861 5627 55919 5633
rect 55861 5624 55873 5627
rect 55456 5596 55873 5624
rect 55456 5584 55462 5596
rect 55861 5593 55873 5596
rect 55907 5593 55919 5627
rect 55861 5587 55919 5593
rect 77680 5568 77708 5664
rect 77849 5661 77861 5664
rect 77895 5661 77907 5695
rect 78048 5692 78076 5791
rect 78217 5695 78275 5701
rect 78217 5692 78229 5695
rect 78048 5664 78229 5692
rect 77849 5655 77907 5661
rect 78217 5661 78229 5664
rect 78263 5661 78275 5695
rect 78217 5655 78275 5661
rect 55493 5559 55551 5565
rect 55493 5556 55505 5559
rect 53800 5528 55505 5556
rect 53800 5516 53806 5528
rect 55493 5525 55505 5528
rect 55539 5556 55551 5559
rect 55766 5556 55772 5568
rect 55539 5528 55772 5556
rect 55539 5525 55551 5528
rect 55493 5519 55551 5525
rect 55766 5516 55772 5528
rect 55824 5556 55830 5568
rect 56137 5559 56195 5565
rect 56137 5556 56149 5559
rect 55824 5528 56149 5556
rect 55824 5516 55830 5528
rect 56137 5525 56149 5528
rect 56183 5525 56195 5559
rect 56137 5519 56195 5525
rect 77662 5516 77668 5568
rect 77720 5516 77726 5568
rect 78398 5516 78404 5568
rect 78456 5516 78462 5568
rect 1104 5466 78844 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 66314 5466
rect 66366 5414 66378 5466
rect 66430 5414 66442 5466
rect 66494 5414 66506 5466
rect 66558 5414 66570 5466
rect 66622 5414 78844 5466
rect 1104 5392 78844 5414
rect 30650 5312 30656 5364
rect 30708 5352 30714 5364
rect 30929 5355 30987 5361
rect 30929 5352 30941 5355
rect 30708 5324 30941 5352
rect 30708 5312 30714 5324
rect 30929 5321 30941 5324
rect 30975 5321 30987 5355
rect 30929 5315 30987 5321
rect 36262 5312 36268 5364
rect 36320 5312 36326 5364
rect 36538 5312 36544 5364
rect 36596 5352 36602 5364
rect 36817 5355 36875 5361
rect 36817 5352 36829 5355
rect 36596 5324 36829 5352
rect 36596 5312 36602 5324
rect 36817 5321 36829 5324
rect 36863 5352 36875 5355
rect 36906 5352 36912 5364
rect 36863 5324 36912 5352
rect 36863 5321 36875 5324
rect 36817 5315 36875 5321
rect 36906 5312 36912 5324
rect 36964 5312 36970 5364
rect 42610 5312 42616 5364
rect 42668 5352 42674 5364
rect 43533 5355 43591 5361
rect 43533 5352 43545 5355
rect 42668 5324 43545 5352
rect 42668 5312 42674 5324
rect 33686 5284 33692 5296
rect 33336 5256 33692 5284
rect 30926 5176 30932 5228
rect 30984 5216 30990 5228
rect 31113 5219 31171 5225
rect 31113 5216 31125 5219
rect 30984 5188 31125 5216
rect 30984 5176 30990 5188
rect 31113 5185 31125 5188
rect 31159 5185 31171 5219
rect 31113 5179 31171 5185
rect 31202 5176 31208 5228
rect 31260 5176 31266 5228
rect 31481 5219 31539 5225
rect 31481 5185 31493 5219
rect 31527 5216 31539 5219
rect 32030 5216 32036 5228
rect 31527 5188 32036 5216
rect 31527 5185 31539 5188
rect 31481 5179 31539 5185
rect 32030 5176 32036 5188
rect 32088 5176 32094 5228
rect 33134 5176 33140 5228
rect 33192 5176 33198 5228
rect 33336 5225 33364 5256
rect 33686 5244 33692 5256
rect 33744 5244 33750 5296
rect 34422 5284 34428 5296
rect 34348 5256 34428 5284
rect 34348 5225 34376 5256
rect 34422 5244 34428 5256
rect 34480 5284 34486 5296
rect 34977 5287 35035 5293
rect 34977 5284 34989 5287
rect 34480 5256 34989 5284
rect 34480 5244 34486 5256
rect 34977 5253 34989 5256
rect 35023 5253 35035 5287
rect 36280 5284 36308 5312
rect 38378 5284 38384 5296
rect 36280 5256 38384 5284
rect 34977 5247 35035 5253
rect 33321 5219 33379 5225
rect 33321 5185 33333 5219
rect 33367 5185 33379 5219
rect 33321 5179 33379 5185
rect 34333 5219 34391 5225
rect 34333 5185 34345 5219
rect 34379 5185 34391 5219
rect 34333 5179 34391 5185
rect 34701 5219 34759 5225
rect 34701 5185 34713 5219
rect 34747 5185 34759 5219
rect 34701 5179 34759 5185
rect 31389 5151 31447 5157
rect 31389 5117 31401 5151
rect 31435 5148 31447 5151
rect 33336 5148 33364 5179
rect 31435 5120 33364 5148
rect 33413 5151 33471 5157
rect 31435 5117 31447 5120
rect 31389 5111 31447 5117
rect 33413 5117 33425 5151
rect 33459 5148 33471 5151
rect 33689 5151 33747 5157
rect 33689 5148 33701 5151
rect 33459 5120 33701 5148
rect 33459 5117 33471 5120
rect 33413 5111 33471 5117
rect 33689 5117 33701 5120
rect 33735 5117 33747 5151
rect 34716 5148 34744 5179
rect 34882 5176 34888 5228
rect 34940 5176 34946 5228
rect 35069 5219 35127 5225
rect 35069 5185 35081 5219
rect 35115 5216 35127 5219
rect 35158 5216 35164 5228
rect 35115 5188 35164 5216
rect 35115 5185 35127 5188
rect 35069 5179 35127 5185
rect 35158 5176 35164 5188
rect 35216 5216 35222 5228
rect 36170 5216 36176 5228
rect 35216 5188 36176 5216
rect 35216 5176 35222 5188
rect 36170 5176 36176 5188
rect 36228 5216 36234 5228
rect 36265 5219 36323 5225
rect 36265 5216 36277 5219
rect 36228 5188 36277 5216
rect 36228 5176 36234 5188
rect 36265 5185 36277 5188
rect 36311 5185 36323 5219
rect 36265 5179 36323 5185
rect 36354 5176 36360 5228
rect 36412 5176 36418 5228
rect 36449 5219 36507 5225
rect 36449 5185 36461 5219
rect 36495 5216 36507 5219
rect 36538 5216 36544 5228
rect 36495 5188 36544 5216
rect 36495 5185 36507 5188
rect 36449 5179 36507 5185
rect 36538 5176 36544 5188
rect 36596 5176 36602 5228
rect 36648 5225 36676 5256
rect 38378 5244 38384 5256
rect 38436 5284 38442 5296
rect 38436 5256 38884 5284
rect 38436 5244 38442 5256
rect 36633 5219 36691 5225
rect 36633 5185 36645 5219
rect 36679 5185 36691 5219
rect 36633 5179 36691 5185
rect 37001 5219 37059 5225
rect 37001 5185 37013 5219
rect 37047 5216 37059 5219
rect 37366 5216 37372 5228
rect 37047 5188 37372 5216
rect 37047 5185 37059 5188
rect 37001 5179 37059 5185
rect 37090 5148 37096 5160
rect 34716 5120 37096 5148
rect 33689 5111 33747 5117
rect 37090 5108 37096 5120
rect 37148 5108 37154 5160
rect 35986 5040 35992 5092
rect 36044 5080 36050 5092
rect 37200 5080 37228 5188
rect 37366 5176 37372 5188
rect 37424 5176 37430 5228
rect 37458 5176 37464 5228
rect 37516 5176 37522 5228
rect 38856 5225 38884 5256
rect 41874 5244 41880 5296
rect 41932 5284 41938 5296
rect 42886 5284 42892 5296
rect 41932 5256 42892 5284
rect 41932 5244 41938 5256
rect 42886 5244 42892 5256
rect 42944 5244 42950 5296
rect 42996 5293 43024 5324
rect 43533 5321 43545 5324
rect 43579 5321 43591 5355
rect 43533 5315 43591 5321
rect 43993 5355 44051 5361
rect 43993 5321 44005 5355
rect 44039 5352 44051 5355
rect 44174 5352 44180 5364
rect 44039 5324 44180 5352
rect 44039 5321 44051 5324
rect 43993 5315 44051 5321
rect 42981 5287 43039 5293
rect 42981 5253 42993 5287
rect 43027 5284 43039 5287
rect 44008 5284 44036 5315
rect 44174 5312 44180 5324
rect 44232 5312 44238 5364
rect 53098 5312 53104 5364
rect 53156 5352 53162 5364
rect 53156 5324 53328 5352
rect 53156 5312 53162 5324
rect 43027 5256 43061 5284
rect 43272 5256 44036 5284
rect 43027 5253 43039 5256
rect 42981 5247 43039 5253
rect 38841 5219 38899 5225
rect 38841 5185 38853 5219
rect 38887 5185 38899 5219
rect 38841 5179 38899 5185
rect 41782 5176 41788 5228
rect 41840 5216 41846 5228
rect 42751 5219 42809 5225
rect 42751 5216 42763 5219
rect 41840 5188 42763 5216
rect 41840 5176 41846 5188
rect 42751 5185 42763 5188
rect 42797 5185 42809 5219
rect 42751 5179 42809 5185
rect 43070 5176 43076 5228
rect 43128 5225 43134 5228
rect 43272 5225 43300 5256
rect 44542 5244 44548 5296
rect 44600 5284 44606 5296
rect 44600 5256 51120 5284
rect 44600 5244 44606 5256
rect 43128 5219 43167 5225
rect 43155 5185 43167 5219
rect 43128 5179 43167 5185
rect 43257 5219 43315 5225
rect 43257 5185 43269 5219
rect 43303 5185 43315 5219
rect 43257 5179 43315 5185
rect 43441 5219 43499 5225
rect 43441 5185 43453 5219
rect 43487 5216 43499 5219
rect 43898 5216 43904 5228
rect 43487 5188 43904 5216
rect 43487 5185 43499 5188
rect 43441 5179 43499 5185
rect 43128 5176 43152 5179
rect 43898 5176 43904 5188
rect 43956 5216 43962 5228
rect 44085 5219 44143 5225
rect 44085 5216 44097 5219
rect 43956 5188 44097 5216
rect 43956 5176 43962 5188
rect 44085 5185 44097 5188
rect 44131 5216 44143 5219
rect 49510 5216 49516 5228
rect 44131 5188 49516 5216
rect 44131 5185 44143 5188
rect 44085 5179 44143 5185
rect 49510 5176 49516 5188
rect 49568 5176 49574 5228
rect 49694 5176 49700 5228
rect 49752 5176 49758 5228
rect 50709 5219 50767 5225
rect 50709 5185 50721 5219
rect 50755 5216 50767 5219
rect 50982 5216 50988 5228
rect 50755 5188 50988 5216
rect 50755 5185 50767 5188
rect 50709 5179 50767 5185
rect 50982 5176 50988 5188
rect 51040 5176 51046 5228
rect 37737 5151 37795 5157
rect 37737 5117 37749 5151
rect 37783 5148 37795 5151
rect 38289 5151 38347 5157
rect 38289 5148 38301 5151
rect 37783 5120 38301 5148
rect 37783 5117 37795 5120
rect 37737 5111 37795 5117
rect 38289 5117 38301 5120
rect 38335 5117 38347 5151
rect 43124 5148 43152 5176
rect 45646 5148 45652 5160
rect 43124 5120 45652 5148
rect 38289 5111 38347 5117
rect 45646 5108 45652 5120
rect 45704 5108 45710 5160
rect 49786 5108 49792 5160
rect 49844 5148 49850 5160
rect 49881 5151 49939 5157
rect 49881 5148 49893 5151
rect 49844 5120 49893 5148
rect 49844 5108 49850 5120
rect 49881 5117 49893 5120
rect 49927 5117 49939 5151
rect 49881 5111 49939 5117
rect 49973 5151 50031 5157
rect 49973 5117 49985 5151
rect 50019 5148 50031 5151
rect 50065 5151 50123 5157
rect 50065 5148 50077 5151
rect 50019 5120 50077 5148
rect 50019 5117 50031 5120
rect 49973 5111 50031 5117
rect 50065 5117 50077 5120
rect 50111 5117 50123 5151
rect 50065 5111 50123 5117
rect 36044 5052 37228 5080
rect 36044 5040 36050 5052
rect 32306 4972 32312 5024
rect 32364 5012 32370 5024
rect 32953 5015 33011 5021
rect 32953 5012 32965 5015
rect 32364 4984 32965 5012
rect 32364 4972 32370 4984
rect 32953 4981 32965 4984
rect 32999 4981 33011 5015
rect 32953 4975 33011 4981
rect 35253 5015 35311 5021
rect 35253 4981 35265 5015
rect 35299 5012 35311 5015
rect 35526 5012 35532 5024
rect 35299 4984 35532 5012
rect 35299 4981 35311 4984
rect 35253 4975 35311 4981
rect 35526 4972 35532 4984
rect 35584 4972 35590 5024
rect 36081 5015 36139 5021
rect 36081 4981 36093 5015
rect 36127 5012 36139 5015
rect 36446 5012 36452 5024
rect 36127 4984 36452 5012
rect 36127 4981 36139 4984
rect 36081 4975 36139 4981
rect 36446 4972 36452 4984
rect 36504 4972 36510 5024
rect 37182 4972 37188 5024
rect 37240 5012 37246 5024
rect 37277 5015 37335 5021
rect 37277 5012 37289 5015
rect 37240 4984 37289 5012
rect 37240 4972 37246 4984
rect 37277 4981 37289 4984
rect 37323 4981 37335 5015
rect 37277 4975 37335 4981
rect 37550 4972 37556 5024
rect 37608 5012 37614 5024
rect 37645 5015 37703 5021
rect 37645 5012 37657 5015
rect 37608 4984 37657 5012
rect 37608 4972 37614 4984
rect 37645 4981 37657 4984
rect 37691 4981 37703 5015
rect 37645 4975 37703 4981
rect 42613 5015 42671 5021
rect 42613 4981 42625 5015
rect 42659 5012 42671 5015
rect 43438 5012 43444 5024
rect 42659 4984 43444 5012
rect 42659 4981 42671 4984
rect 42613 4975 42671 4981
rect 43438 4972 43444 4984
rect 43496 4972 43502 5024
rect 46290 4972 46296 5024
rect 46348 5012 46354 5024
rect 47394 5012 47400 5024
rect 46348 4984 47400 5012
rect 46348 4972 46354 4984
rect 47394 4972 47400 4984
rect 47452 4972 47458 5024
rect 49510 4972 49516 5024
rect 49568 4972 49574 5024
rect 49896 5012 49924 5111
rect 51092 5080 51120 5256
rect 51442 5244 51448 5296
rect 51500 5284 51506 5296
rect 53300 5293 53328 5324
rect 53285 5287 53343 5293
rect 51500 5256 52040 5284
rect 51500 5244 51506 5256
rect 51902 5176 51908 5228
rect 51960 5176 51966 5228
rect 52012 5225 52040 5256
rect 53285 5253 53297 5287
rect 53331 5253 53343 5287
rect 53285 5247 53343 5253
rect 51997 5219 52055 5225
rect 51997 5185 52009 5219
rect 52043 5185 52055 5219
rect 51997 5179 52055 5185
rect 52273 5219 52331 5225
rect 52273 5185 52285 5219
rect 52319 5216 52331 5219
rect 52822 5216 52828 5228
rect 52319 5188 52828 5216
rect 52319 5185 52331 5188
rect 52273 5179 52331 5185
rect 52822 5176 52828 5188
rect 52880 5176 52886 5228
rect 54665 5219 54723 5225
rect 54665 5185 54677 5219
rect 54711 5216 54723 5219
rect 55122 5216 55128 5228
rect 54711 5188 55128 5216
rect 54711 5185 54723 5188
rect 54665 5179 54723 5185
rect 55122 5176 55128 5188
rect 55180 5176 55186 5228
rect 78033 5219 78091 5225
rect 78033 5185 78045 5219
rect 78079 5216 78091 5219
rect 78306 5216 78312 5228
rect 78079 5188 78312 5216
rect 78079 5185 78091 5188
rect 78033 5179 78091 5185
rect 78306 5176 78312 5188
rect 78364 5176 78370 5228
rect 51718 5108 51724 5160
rect 51776 5108 51782 5160
rect 52086 5108 52092 5160
rect 52144 5148 52150 5160
rect 53374 5148 53380 5160
rect 52144 5120 53380 5148
rect 52144 5108 52150 5120
rect 53374 5108 53380 5120
rect 53432 5148 53438 5160
rect 54113 5151 54171 5157
rect 54113 5148 54125 5151
rect 53432 5120 54125 5148
rect 53432 5108 53438 5120
rect 54113 5117 54125 5120
rect 54159 5148 54171 5151
rect 56042 5148 56048 5160
rect 54159 5120 56048 5148
rect 54159 5117 54171 5120
rect 54113 5111 54171 5117
rect 56042 5108 56048 5120
rect 56100 5108 56106 5160
rect 54849 5083 54907 5089
rect 54849 5080 54861 5083
rect 51092 5052 54861 5080
rect 54849 5049 54861 5052
rect 54895 5080 54907 5083
rect 55398 5080 55404 5092
rect 54895 5052 55404 5080
rect 54895 5049 54907 5052
rect 54849 5043 54907 5049
rect 55398 5040 55404 5052
rect 55456 5040 55462 5092
rect 52181 5015 52239 5021
rect 52181 5012 52193 5015
rect 49896 4984 52193 5012
rect 52181 4981 52193 4984
rect 52227 5012 52239 5015
rect 52546 5012 52552 5024
rect 52227 4984 52552 5012
rect 52227 4981 52239 4984
rect 52181 4975 52239 4981
rect 52546 4972 52552 4984
rect 52604 4972 52610 5024
rect 78122 4972 78128 5024
rect 78180 4972 78186 5024
rect 1104 4922 78844 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 78844 4922
rect 1104 4848 78844 4870
rect 29917 4811 29975 4817
rect 29917 4777 29929 4811
rect 29963 4808 29975 4811
rect 30006 4808 30012 4820
rect 29963 4780 30012 4808
rect 29963 4777 29975 4780
rect 29917 4771 29975 4777
rect 30006 4768 30012 4780
rect 30064 4768 30070 4820
rect 43622 4808 43628 4820
rect 33704 4780 43628 4808
rect 30282 4632 30288 4684
rect 30340 4672 30346 4684
rect 32033 4675 32091 4681
rect 32033 4672 32045 4675
rect 30340 4644 32045 4672
rect 30340 4632 30346 4644
rect 32033 4641 32045 4644
rect 32079 4641 32091 4675
rect 32033 4635 32091 4641
rect 32306 4632 32312 4684
rect 32364 4632 32370 4684
rect 30006 4564 30012 4616
rect 30064 4564 30070 4616
rect 30193 4607 30251 4613
rect 30193 4573 30205 4607
rect 30239 4604 30251 4607
rect 31478 4604 31484 4616
rect 30239 4576 31484 4604
rect 30239 4573 30251 4576
rect 30193 4567 30251 4573
rect 31478 4564 31484 4576
rect 31536 4564 31542 4616
rect 33594 4536 33600 4548
rect 33534 4508 33600 4536
rect 33594 4496 33600 4508
rect 33652 4496 33658 4548
rect 30101 4471 30159 4477
rect 30101 4437 30113 4471
rect 30147 4468 30159 4471
rect 31662 4468 31668 4480
rect 30147 4440 31668 4468
rect 30147 4437 30159 4440
rect 30101 4431 30159 4437
rect 31662 4428 31668 4440
rect 31720 4468 31726 4480
rect 33704 4468 33732 4780
rect 43622 4768 43628 4780
rect 43680 4768 43686 4820
rect 44545 4811 44603 4817
rect 44545 4777 44557 4811
rect 44591 4808 44603 4811
rect 44726 4808 44732 4820
rect 44591 4780 44732 4808
rect 44591 4777 44603 4780
rect 44545 4771 44603 4777
rect 44726 4768 44732 4780
rect 44784 4768 44790 4820
rect 44818 4768 44824 4820
rect 44876 4808 44882 4820
rect 44876 4780 47164 4808
rect 44876 4768 44882 4780
rect 33781 4743 33839 4749
rect 33781 4709 33793 4743
rect 33827 4740 33839 4743
rect 34422 4740 34428 4752
rect 33827 4712 34428 4740
rect 33827 4709 33839 4712
rect 33781 4703 33839 4709
rect 34422 4700 34428 4712
rect 34480 4700 34486 4752
rect 34624 4712 35848 4740
rect 34054 4632 34060 4684
rect 34112 4672 34118 4684
rect 34624 4672 34652 4712
rect 35713 4675 35771 4681
rect 35713 4672 35725 4675
rect 34112 4644 34652 4672
rect 34716 4644 35725 4672
rect 34112 4632 34118 4644
rect 33778 4564 33784 4616
rect 33836 4604 33842 4616
rect 34716 4604 34744 4644
rect 35713 4641 35725 4644
rect 35759 4641 35771 4675
rect 35713 4635 35771 4641
rect 33836 4576 34744 4604
rect 35437 4607 35495 4613
rect 33836 4564 33842 4576
rect 35437 4573 35449 4607
rect 35483 4573 35495 4607
rect 35437 4567 35495 4573
rect 31720 4440 33732 4468
rect 31720 4428 31726 4440
rect 35250 4428 35256 4480
rect 35308 4428 35314 4480
rect 35452 4468 35480 4567
rect 35526 4564 35532 4616
rect 35584 4564 35590 4616
rect 35820 4613 35848 4712
rect 38378 4700 38384 4752
rect 38436 4740 38442 4752
rect 38657 4743 38715 4749
rect 38657 4740 38669 4743
rect 38436 4712 38669 4740
rect 38436 4700 38442 4712
rect 38657 4709 38669 4712
rect 38703 4709 38715 4743
rect 38657 4703 38715 4709
rect 41322 4700 41328 4752
rect 41380 4740 41386 4752
rect 41601 4743 41659 4749
rect 41601 4740 41613 4743
rect 41380 4712 41613 4740
rect 41380 4700 41386 4712
rect 41601 4709 41613 4712
rect 41647 4740 41659 4743
rect 41966 4740 41972 4752
rect 41647 4712 41972 4740
rect 41647 4709 41659 4712
rect 41601 4703 41659 4709
rect 41966 4700 41972 4712
rect 42024 4740 42030 4752
rect 42024 4712 42288 4740
rect 42024 4700 42030 4712
rect 37182 4632 37188 4684
rect 37240 4632 37246 4684
rect 40770 4632 40776 4684
rect 40828 4672 40834 4684
rect 42260 4681 42288 4712
rect 41693 4675 41751 4681
rect 41693 4672 41705 4675
rect 40828 4644 41705 4672
rect 40828 4632 40834 4644
rect 41693 4641 41705 4644
rect 41739 4641 41751 4675
rect 41693 4635 41751 4641
rect 42245 4675 42303 4681
rect 42245 4641 42257 4675
rect 42291 4641 42303 4675
rect 42245 4635 42303 4641
rect 44266 4632 44272 4684
rect 44324 4632 44330 4684
rect 45830 4672 45836 4684
rect 45204 4644 45836 4672
rect 35805 4607 35863 4613
rect 35805 4573 35817 4607
rect 35851 4604 35863 4607
rect 36354 4604 36360 4616
rect 35851 4576 36360 4604
rect 35851 4573 35863 4576
rect 35805 4567 35863 4573
rect 36354 4564 36360 4576
rect 36412 4564 36418 4616
rect 36909 4607 36967 4613
rect 36909 4573 36921 4607
rect 36955 4573 36967 4607
rect 36909 4567 36967 4573
rect 35897 4539 35955 4545
rect 35897 4505 35909 4539
rect 35943 4536 35955 4539
rect 35986 4536 35992 4548
rect 35943 4508 35992 4536
rect 35943 4505 35955 4508
rect 35897 4499 35955 4505
rect 35986 4496 35992 4508
rect 36044 4496 36050 4548
rect 36078 4496 36084 4548
rect 36136 4536 36142 4548
rect 36633 4539 36691 4545
rect 36633 4536 36645 4539
rect 36136 4508 36645 4536
rect 36136 4496 36142 4508
rect 36633 4505 36645 4508
rect 36679 4536 36691 4539
rect 36924 4536 36952 4567
rect 39850 4564 39856 4616
rect 39908 4564 39914 4616
rect 41230 4564 41236 4616
rect 41288 4564 41294 4616
rect 42794 4564 42800 4616
rect 42852 4564 42858 4616
rect 44284 4604 44312 4632
rect 44206 4576 44312 4604
rect 44818 4564 44824 4616
rect 44876 4604 44882 4616
rect 45204 4613 45232 4644
rect 45830 4632 45836 4644
rect 45888 4672 45894 4684
rect 46842 4672 46848 4684
rect 45888 4644 46848 4672
rect 45888 4632 45894 4644
rect 46842 4632 46848 4644
rect 46900 4632 46906 4684
rect 45005 4607 45063 4613
rect 45005 4604 45017 4607
rect 44876 4576 45017 4604
rect 44876 4564 44882 4576
rect 45005 4573 45017 4576
rect 45051 4573 45063 4607
rect 45005 4567 45063 4573
rect 45189 4607 45247 4613
rect 45189 4573 45201 4607
rect 45235 4573 45247 4607
rect 45189 4567 45247 4573
rect 45373 4607 45431 4613
rect 45373 4573 45385 4607
rect 45419 4604 45431 4607
rect 45554 4604 45560 4616
rect 45419 4576 45560 4604
rect 45419 4573 45431 4576
rect 45373 4567 45431 4573
rect 36679 4508 36952 4536
rect 36679 4505 36691 4508
rect 36633 4499 36691 4505
rect 37642 4496 37648 4548
rect 37700 4496 37706 4548
rect 40126 4496 40132 4548
rect 40184 4496 40190 4548
rect 36354 4468 36360 4480
rect 35452 4440 36360 4468
rect 36354 4428 36360 4440
rect 36412 4428 36418 4480
rect 41248 4468 41276 4564
rect 43070 4496 43076 4548
rect 43128 4496 43134 4548
rect 45281 4539 45339 4545
rect 45281 4505 45293 4539
rect 45327 4505 45339 4539
rect 45388 4536 45416 4567
rect 45554 4564 45560 4576
rect 45612 4564 45618 4616
rect 46106 4564 46112 4616
rect 46164 4604 46170 4616
rect 46661 4607 46719 4613
rect 46661 4604 46673 4607
rect 46164 4576 46673 4604
rect 46164 4564 46170 4576
rect 46661 4573 46673 4576
rect 46707 4573 46719 4607
rect 47029 4607 47087 4613
rect 47029 4604 47041 4607
rect 46661 4567 46719 4573
rect 46768 4576 47041 4604
rect 46768 4536 46796 4576
rect 47029 4573 47041 4576
rect 47075 4573 47087 4607
rect 47136 4604 47164 4780
rect 47394 4768 47400 4820
rect 47452 4768 47458 4820
rect 49510 4768 49516 4820
rect 49568 4808 49574 4820
rect 51641 4811 51699 4817
rect 51641 4808 51653 4811
rect 49568 4780 51653 4808
rect 49568 4768 49574 4780
rect 51641 4777 51653 4780
rect 51687 4777 51699 4811
rect 51641 4771 51699 4777
rect 53377 4811 53435 4817
rect 53377 4777 53389 4811
rect 53423 4808 53435 4811
rect 53558 4808 53564 4820
rect 53423 4780 53564 4808
rect 53423 4777 53435 4780
rect 53377 4771 53435 4777
rect 53558 4768 53564 4780
rect 53616 4768 53622 4820
rect 47213 4743 47271 4749
rect 47213 4709 47225 4743
rect 47259 4740 47271 4743
rect 47259 4712 47532 4740
rect 47259 4709 47271 4712
rect 47213 4703 47271 4709
rect 47302 4604 47308 4616
rect 47136 4576 47308 4604
rect 47029 4567 47087 4573
rect 47302 4564 47308 4576
rect 47360 4564 47366 4616
rect 47504 4604 47532 4712
rect 52546 4700 52552 4752
rect 52604 4740 52610 4752
rect 53837 4743 53895 4749
rect 53837 4740 53849 4743
rect 52604 4712 53849 4740
rect 52604 4700 52610 4712
rect 53837 4709 53849 4712
rect 53883 4709 53895 4743
rect 53837 4703 53895 4709
rect 50157 4675 50215 4681
rect 50157 4641 50169 4675
rect 50203 4672 50215 4675
rect 50982 4672 50988 4684
rect 50203 4644 50988 4672
rect 50203 4641 50215 4644
rect 50157 4635 50215 4641
rect 50982 4632 50988 4644
rect 51040 4632 51046 4684
rect 51905 4675 51963 4681
rect 51905 4641 51917 4675
rect 51951 4672 51963 4675
rect 52086 4672 52092 4684
rect 51951 4644 52092 4672
rect 51951 4641 51963 4644
rect 51905 4635 51963 4641
rect 52086 4632 52092 4644
rect 52144 4632 52150 4684
rect 54754 4672 54760 4684
rect 53576 4644 54760 4672
rect 47581 4607 47639 4613
rect 47581 4604 47593 4607
rect 47504 4576 47593 4604
rect 47581 4573 47593 4576
rect 47627 4573 47639 4607
rect 47581 4567 47639 4573
rect 47670 4564 47676 4616
rect 47728 4564 47734 4616
rect 51994 4564 52000 4616
rect 52052 4604 52058 4616
rect 53576 4613 53604 4644
rect 54754 4632 54760 4644
rect 54812 4632 54818 4684
rect 53561 4607 53619 4613
rect 53561 4604 53573 4607
rect 52052 4576 53573 4604
rect 52052 4564 52058 4576
rect 53561 4573 53573 4576
rect 53607 4573 53619 4607
rect 53561 4567 53619 4573
rect 53650 4564 53656 4616
rect 53708 4564 53714 4616
rect 53929 4607 53987 4613
rect 53929 4573 53941 4607
rect 53975 4604 53987 4607
rect 55030 4604 55036 4616
rect 53975 4576 55036 4604
rect 53975 4573 53987 4576
rect 53929 4567 53987 4573
rect 45388 4508 46796 4536
rect 45281 4499 45339 4505
rect 42978 4468 42984 4480
rect 41248 4440 42984 4468
rect 42978 4428 42984 4440
rect 43036 4428 43042 4480
rect 44726 4428 44732 4480
rect 44784 4468 44790 4480
rect 45296 4468 45324 4499
rect 46842 4496 46848 4548
rect 46900 4496 46906 4548
rect 46937 4539 46995 4545
rect 46937 4505 46949 4539
rect 46983 4505 46995 4539
rect 46937 4499 46995 4505
rect 44784 4440 45324 4468
rect 44784 4428 44790 4440
rect 45554 4428 45560 4480
rect 45612 4428 45618 4480
rect 45646 4428 45652 4480
rect 45704 4468 45710 4480
rect 46750 4468 46756 4480
rect 45704 4440 46756 4468
rect 45704 4428 45710 4440
rect 46750 4428 46756 4440
rect 46808 4468 46814 4480
rect 46952 4468 46980 4499
rect 49970 4496 49976 4548
rect 50028 4536 50034 4548
rect 50338 4536 50344 4548
rect 50028 4508 50344 4536
rect 50028 4496 50034 4508
rect 50338 4496 50344 4508
rect 50396 4536 50402 4548
rect 50396 4508 50462 4536
rect 50396 4496 50402 4508
rect 51534 4496 51540 4548
rect 51592 4536 51598 4548
rect 53944 4536 53972 4567
rect 55030 4564 55036 4576
rect 55088 4564 55094 4616
rect 78217 4607 78275 4613
rect 78217 4573 78229 4607
rect 78263 4604 78275 4607
rect 78490 4604 78496 4616
rect 78263 4576 78496 4604
rect 78263 4573 78275 4576
rect 78217 4567 78275 4573
rect 78490 4564 78496 4576
rect 78548 4564 78554 4616
rect 51592 4508 53972 4536
rect 51592 4496 51598 4508
rect 46808 4440 46980 4468
rect 47857 4471 47915 4477
rect 46808 4428 46814 4440
rect 47857 4437 47869 4471
rect 47903 4468 47915 4471
rect 49050 4468 49056 4480
rect 47903 4440 49056 4468
rect 47903 4437 47915 4440
rect 47857 4431 47915 4437
rect 49050 4428 49056 4440
rect 49108 4428 49114 4480
rect 78306 4428 78312 4480
rect 78364 4428 78370 4480
rect 1104 4378 78844 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 66314 4378
rect 66366 4326 66378 4378
rect 66430 4326 66442 4378
rect 66494 4326 66506 4378
rect 66558 4326 66570 4378
rect 66622 4326 78844 4378
rect 1104 4304 78844 4326
rect 34532 4236 35940 4264
rect 33594 4156 33600 4208
rect 33652 4196 33658 4208
rect 34532 4196 34560 4236
rect 35912 4196 35940 4236
rect 35986 4224 35992 4276
rect 36044 4264 36050 4276
rect 36909 4267 36967 4273
rect 36909 4264 36921 4267
rect 36044 4236 36921 4264
rect 36044 4224 36050 4236
rect 36909 4233 36921 4236
rect 36955 4264 36967 4267
rect 37826 4264 37832 4276
rect 36955 4236 37832 4264
rect 36955 4233 36967 4236
rect 36909 4227 36967 4233
rect 37826 4224 37832 4236
rect 37884 4224 37890 4276
rect 40126 4224 40132 4276
rect 40184 4264 40190 4276
rect 40497 4267 40555 4273
rect 40497 4264 40509 4267
rect 40184 4236 40509 4264
rect 40184 4224 40190 4236
rect 40497 4233 40509 4236
rect 40543 4233 40555 4267
rect 40497 4227 40555 4233
rect 43070 4224 43076 4276
rect 43128 4264 43134 4276
rect 43349 4267 43407 4273
rect 43349 4264 43361 4267
rect 43128 4236 43361 4264
rect 43128 4224 43134 4236
rect 43349 4233 43361 4236
rect 43395 4233 43407 4267
rect 43349 4227 43407 4233
rect 47302 4224 47308 4276
rect 47360 4264 47366 4276
rect 47581 4267 47639 4273
rect 47581 4264 47593 4267
rect 47360 4236 47593 4264
rect 47360 4224 47366 4236
rect 47581 4233 47593 4236
rect 47627 4233 47639 4267
rect 47581 4227 47639 4233
rect 36262 4196 36268 4208
rect 33652 4168 34638 4196
rect 35912 4168 36268 4196
rect 33652 4156 33658 4168
rect 36262 4156 36268 4168
rect 36320 4196 36326 4208
rect 37642 4196 37648 4208
rect 36320 4168 37648 4196
rect 36320 4156 36326 4168
rect 37642 4156 37648 4168
rect 37700 4196 37706 4208
rect 38194 4196 38200 4208
rect 37700 4168 38200 4196
rect 37700 4156 37706 4168
rect 38194 4156 38200 4168
rect 38252 4156 38258 4208
rect 39574 4156 39580 4208
rect 39632 4196 39638 4208
rect 39632 4168 41276 4196
rect 39632 4156 39638 4168
rect 30834 4088 30840 4140
rect 30892 4128 30898 4140
rect 31481 4131 31539 4137
rect 31481 4128 31493 4131
rect 30892 4100 31493 4128
rect 30892 4088 30898 4100
rect 31481 4097 31493 4100
rect 31527 4128 31539 4131
rect 31527 4100 31984 4128
rect 31527 4097 31539 4100
rect 31481 4091 31539 4097
rect 31956 3936 31984 4100
rect 36078 4088 36084 4140
rect 36136 4088 36142 4140
rect 36354 4088 36360 4140
rect 36412 4088 36418 4140
rect 36446 4088 36452 4140
rect 36504 4088 36510 4140
rect 36725 4131 36783 4137
rect 36725 4097 36737 4131
rect 36771 4128 36783 4131
rect 37277 4131 37335 4137
rect 37277 4128 37289 4131
rect 36771 4100 37289 4128
rect 36771 4097 36783 4100
rect 36725 4091 36783 4097
rect 37277 4097 37289 4100
rect 37323 4097 37335 4131
rect 37277 4091 37335 4097
rect 40681 4131 40739 4137
rect 40681 4097 40693 4131
rect 40727 4128 40739 4131
rect 41138 4128 41144 4140
rect 40727 4100 41144 4128
rect 40727 4097 40739 4100
rect 40681 4091 40739 4097
rect 41138 4088 41144 4100
rect 41196 4088 41202 4140
rect 41248 4137 41276 4168
rect 41782 4156 41788 4208
rect 41840 4196 41846 4208
rect 41840 4168 41920 4196
rect 41840 4156 41846 4168
rect 41892 4137 41920 4168
rect 41966 4156 41972 4208
rect 42024 4156 42030 4208
rect 42610 4196 42616 4208
rect 42076 4168 42616 4196
rect 42076 4137 42104 4168
rect 42610 4156 42616 4168
rect 42668 4156 42674 4208
rect 47762 4156 47768 4208
rect 47820 4196 47826 4208
rect 47820 4168 47886 4196
rect 47820 4156 47826 4168
rect 41233 4131 41291 4137
rect 41233 4097 41245 4131
rect 41279 4097 41291 4131
rect 41233 4091 41291 4097
rect 41325 4131 41383 4137
rect 41325 4097 41337 4131
rect 41371 4097 41383 4131
rect 41325 4091 41383 4097
rect 41601 4131 41659 4137
rect 41601 4097 41613 4131
rect 41647 4128 41659 4131
rect 41877 4131 41935 4137
rect 41647 4100 41828 4128
rect 41647 4097 41659 4100
rect 41601 4091 41659 4097
rect 34054 4020 34060 4072
rect 34112 4060 34118 4072
rect 34333 4063 34391 4069
rect 34333 4060 34345 4063
rect 34112 4032 34345 4060
rect 34112 4020 34118 4032
rect 34333 4029 34345 4032
rect 34379 4029 34391 4063
rect 34333 4023 34391 4029
rect 35250 4020 35256 4072
rect 35308 4060 35314 4072
rect 35805 4063 35863 4069
rect 35805 4060 35817 4063
rect 35308 4032 35817 4060
rect 35308 4020 35314 4032
rect 35805 4029 35817 4032
rect 35851 4029 35863 4063
rect 36372 4060 36400 4088
rect 36372 4032 36492 4060
rect 35805 4023 35863 4029
rect 19702 3884 19708 3936
rect 19760 3924 19766 3936
rect 31665 3927 31723 3933
rect 31665 3924 31677 3927
rect 19760 3896 31677 3924
rect 19760 3884 19766 3896
rect 31665 3893 31677 3896
rect 31711 3924 31723 3927
rect 31846 3924 31852 3936
rect 31711 3896 31852 3924
rect 31711 3893 31723 3896
rect 31665 3887 31723 3893
rect 31846 3884 31852 3896
rect 31904 3884 31910 3936
rect 31938 3884 31944 3936
rect 31996 3884 32002 3936
rect 36170 3884 36176 3936
rect 36228 3884 36234 3936
rect 36464 3924 36492 4032
rect 37090 4020 37096 4072
rect 37148 4060 37154 4072
rect 37829 4063 37887 4069
rect 37829 4060 37841 4063
rect 37148 4032 37841 4060
rect 37148 4020 37154 4032
rect 37829 4029 37841 4032
rect 37875 4029 37887 4063
rect 40957 4063 41015 4069
rect 37829 4023 37887 4029
rect 39684 4032 40908 4060
rect 36633 3995 36691 4001
rect 36633 3961 36645 3995
rect 36679 3992 36691 3995
rect 37550 3992 37556 4004
rect 36679 3964 37556 3992
rect 36679 3961 36691 3964
rect 36633 3955 36691 3961
rect 37550 3952 37556 3964
rect 37608 3992 37614 4004
rect 39684 3992 39712 4032
rect 40880 4004 40908 4032
rect 40957 4029 40969 4063
rect 41003 4029 41015 4063
rect 41340 4060 41368 4091
rect 41800 4060 41828 4100
rect 41877 4097 41889 4131
rect 41923 4097 41935 4131
rect 41877 4091 41935 4097
rect 42061 4131 42119 4137
rect 42061 4097 42073 4131
rect 42107 4097 42119 4131
rect 42061 4091 42119 4097
rect 42245 4131 42303 4137
rect 42245 4097 42257 4131
rect 42291 4128 42303 4131
rect 42291 4100 42840 4128
rect 42291 4097 42303 4100
rect 42245 4091 42303 4097
rect 42613 4063 42671 4069
rect 42613 4060 42625 4063
rect 41340 4032 41736 4060
rect 41800 4032 42625 4060
rect 40957 4023 41015 4029
rect 37608 3964 39712 3992
rect 37608 3952 37614 3964
rect 40862 3952 40868 4004
rect 40920 3952 40926 4004
rect 38838 3924 38844 3936
rect 36464 3896 38844 3924
rect 38838 3884 38844 3896
rect 38896 3924 38902 3936
rect 39574 3924 39580 3936
rect 38896 3896 39580 3924
rect 38896 3884 38902 3896
rect 39574 3884 39580 3896
rect 39632 3884 39638 3936
rect 40770 3884 40776 3936
rect 40828 3924 40834 3936
rect 40972 3924 41000 4023
rect 41708 4001 41736 4032
rect 42613 4029 42625 4032
rect 42659 4029 42671 4063
rect 42812 4060 42840 4100
rect 42886 4088 42892 4140
rect 42944 4128 42950 4140
rect 43165 4131 43223 4137
rect 43165 4128 43177 4131
rect 42944 4100 43177 4128
rect 42944 4088 42950 4100
rect 43165 4097 43177 4100
rect 43211 4097 43223 4131
rect 43165 4091 43223 4097
rect 43438 4088 43444 4140
rect 43496 4128 43502 4140
rect 43533 4131 43591 4137
rect 43533 4128 43545 4131
rect 43496 4100 43545 4128
rect 43496 4088 43502 4100
rect 43533 4097 43545 4100
rect 43579 4097 43591 4131
rect 44726 4128 44732 4140
rect 43533 4091 43591 4097
rect 43640 4100 44732 4128
rect 43640 4060 43668 4100
rect 44726 4088 44732 4100
rect 44784 4088 44790 4140
rect 45281 4131 45339 4137
rect 45281 4097 45293 4131
rect 45327 4097 45339 4131
rect 45281 4091 45339 4097
rect 45373 4131 45431 4137
rect 45373 4097 45385 4131
rect 45419 4128 45431 4131
rect 45554 4128 45560 4140
rect 45419 4100 45560 4128
rect 45419 4097 45431 4100
rect 45373 4091 45431 4097
rect 42812 4032 43668 4060
rect 43809 4063 43867 4069
rect 42613 4023 42671 4029
rect 43809 4029 43821 4063
rect 43855 4060 43867 4063
rect 44085 4063 44143 4069
rect 44085 4060 44097 4063
rect 43855 4032 44097 4060
rect 43855 4029 43867 4032
rect 43809 4023 43867 4029
rect 44085 4029 44097 4032
rect 44131 4029 44143 4063
rect 45296 4060 45324 4091
rect 45554 4088 45560 4100
rect 45612 4088 45618 4140
rect 45646 4088 45652 4140
rect 45704 4088 45710 4140
rect 54018 4088 54024 4140
rect 54076 4128 54082 4140
rect 58437 4131 58495 4137
rect 58437 4128 58449 4131
rect 54076 4100 58449 4128
rect 54076 4088 54082 4100
rect 58437 4097 58449 4100
rect 58483 4128 58495 4131
rect 58621 4131 58679 4137
rect 58621 4128 58633 4131
rect 58483 4100 58633 4128
rect 58483 4097 58495 4100
rect 58437 4091 58495 4097
rect 58621 4097 58633 4100
rect 58667 4128 58679 4131
rect 68186 4128 68192 4140
rect 58667 4100 68192 4128
rect 58667 4097 58679 4100
rect 58621 4091 58679 4097
rect 68186 4088 68192 4100
rect 68244 4088 68250 4140
rect 47118 4060 47124 4072
rect 45296 4032 47124 4060
rect 44085 4023 44143 4029
rect 47118 4020 47124 4032
rect 47176 4060 47182 4072
rect 47670 4060 47676 4072
rect 47176 4032 47676 4060
rect 47176 4020 47182 4032
rect 47670 4020 47676 4032
rect 47728 4020 47734 4072
rect 49050 4020 49056 4072
rect 49108 4020 49114 4072
rect 49329 4063 49387 4069
rect 49329 4029 49341 4063
rect 49375 4060 49387 4063
rect 51074 4060 51080 4072
rect 49375 4032 51080 4060
rect 49375 4029 49387 4032
rect 49329 4023 49387 4029
rect 51074 4020 51080 4032
rect 51132 4060 51138 4072
rect 52086 4060 52092 4072
rect 51132 4032 52092 4060
rect 51132 4020 51138 4032
rect 52086 4020 52092 4032
rect 52144 4020 52150 4072
rect 59354 4020 59360 4072
rect 59412 4060 59418 4072
rect 78306 4060 78312 4072
rect 59412 4032 78312 4060
rect 59412 4020 59418 4032
rect 78306 4020 78312 4032
rect 78364 4020 78370 4072
rect 41693 3995 41751 4001
rect 41693 3961 41705 3995
rect 41739 3961 41751 3995
rect 41693 3955 41751 3961
rect 43714 3952 43720 4004
rect 43772 3992 43778 4004
rect 45557 3995 45615 4001
rect 45557 3992 45569 3995
rect 43772 3964 45569 3992
rect 43772 3952 43778 3964
rect 45557 3961 45569 3964
rect 45603 3992 45615 3995
rect 46290 3992 46296 4004
rect 45603 3964 46296 3992
rect 45603 3961 45615 3964
rect 45557 3955 45615 3961
rect 46290 3952 46296 3964
rect 46348 3952 46354 4004
rect 51442 3952 51448 4004
rect 51500 3992 51506 4004
rect 58253 3995 58311 4001
rect 58253 3992 58265 3995
rect 51500 3964 58265 3992
rect 51500 3952 51506 3964
rect 58253 3961 58265 3964
rect 58299 3992 58311 3995
rect 58986 3992 58992 4004
rect 58299 3964 58992 3992
rect 58299 3961 58311 3964
rect 58253 3955 58311 3961
rect 58986 3952 58992 3964
rect 59044 3952 59050 4004
rect 40828 3896 41000 3924
rect 41049 3927 41107 3933
rect 40828 3884 40834 3896
rect 41049 3893 41061 3927
rect 41095 3924 41107 3927
rect 41414 3924 41420 3936
rect 41095 3896 41420 3924
rect 41095 3893 41107 3896
rect 41049 3887 41107 3893
rect 41414 3884 41420 3896
rect 41472 3884 41478 3936
rect 41506 3884 41512 3936
rect 41564 3884 41570 3936
rect 45097 3927 45155 3933
rect 45097 3893 45109 3927
rect 45143 3924 45155 3927
rect 45278 3924 45284 3936
rect 45143 3896 45284 3924
rect 45143 3893 45155 3896
rect 45097 3887 45155 3893
rect 45278 3884 45284 3896
rect 45336 3884 45342 3936
rect 56410 3884 56416 3936
rect 56468 3884 56474 3936
rect 1104 3834 78844 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 78844 3834
rect 1104 3760 78844 3782
rect 30006 3680 30012 3732
rect 30064 3680 30070 3732
rect 31938 3680 31944 3732
rect 31996 3720 32002 3732
rect 31996 3692 46336 3720
rect 31996 3680 32002 3692
rect 30024 3652 30052 3680
rect 30024 3624 30328 3652
rect 30190 3544 30196 3596
rect 30248 3544 30254 3596
rect 30300 3584 30328 3624
rect 31754 3612 31760 3664
rect 31812 3652 31818 3664
rect 32309 3655 32367 3661
rect 32309 3652 32321 3655
rect 31812 3624 32321 3652
rect 31812 3612 31818 3624
rect 32309 3621 32321 3624
rect 32355 3652 32367 3655
rect 32585 3655 32643 3661
rect 32585 3652 32597 3655
rect 32355 3624 32597 3652
rect 32355 3621 32367 3624
rect 32309 3615 32367 3621
rect 32585 3621 32597 3624
rect 32631 3621 32643 3655
rect 32585 3615 32643 3621
rect 38194 3612 38200 3664
rect 38252 3652 38258 3664
rect 38657 3655 38715 3661
rect 38657 3652 38669 3655
rect 38252 3624 38669 3652
rect 38252 3612 38258 3624
rect 38657 3621 38669 3624
rect 38703 3621 38715 3655
rect 38657 3615 38715 3621
rect 42886 3612 42892 3664
rect 42944 3612 42950 3664
rect 42978 3612 42984 3664
rect 43036 3652 43042 3664
rect 43254 3652 43260 3664
rect 43036 3624 43260 3652
rect 43036 3612 43042 3624
rect 43254 3612 43260 3624
rect 43312 3652 43318 3664
rect 44266 3652 44272 3664
rect 43312 3624 44272 3652
rect 43312 3612 43318 3624
rect 44266 3612 44272 3624
rect 44324 3612 44330 3664
rect 44542 3612 44548 3664
rect 44600 3652 44606 3664
rect 44637 3655 44695 3661
rect 44637 3652 44649 3655
rect 44600 3624 44649 3652
rect 44600 3612 44606 3624
rect 44637 3621 44649 3624
rect 44683 3621 44695 3655
rect 46308 3652 46336 3692
rect 46750 3680 46756 3732
rect 46808 3680 46814 3732
rect 50338 3680 50344 3732
rect 50396 3680 50402 3732
rect 50985 3723 51043 3729
rect 50985 3689 50997 3723
rect 51031 3720 51043 3723
rect 51350 3720 51356 3732
rect 51031 3692 51356 3720
rect 51031 3689 51043 3692
rect 50985 3683 51043 3689
rect 51350 3680 51356 3692
rect 51408 3680 51414 3732
rect 57149 3723 57207 3729
rect 57149 3689 57161 3723
rect 57195 3689 57207 3723
rect 59354 3720 59360 3732
rect 57149 3683 57207 3689
rect 58912 3692 59360 3720
rect 55306 3652 55312 3664
rect 46308 3624 55312 3652
rect 44637 3615 44695 3621
rect 55306 3612 55312 3624
rect 55364 3652 55370 3664
rect 56137 3655 56195 3661
rect 56137 3652 56149 3655
rect 55364 3624 56149 3652
rect 55364 3612 55370 3624
rect 56137 3621 56149 3624
rect 56183 3621 56195 3655
rect 56137 3615 56195 3621
rect 30469 3587 30527 3593
rect 30469 3584 30481 3587
rect 30300 3556 30481 3584
rect 30469 3553 30481 3556
rect 30515 3553 30527 3587
rect 30469 3547 30527 3553
rect 31772 3516 31800 3612
rect 41141 3587 41199 3593
rect 41141 3553 41153 3587
rect 41187 3584 41199 3587
rect 42794 3584 42800 3596
rect 41187 3556 42800 3584
rect 41187 3553 41199 3556
rect 41141 3547 41199 3553
rect 42794 3544 42800 3556
rect 42852 3584 42858 3596
rect 44818 3584 44824 3596
rect 42852 3556 44824 3584
rect 42852 3544 42858 3556
rect 44818 3544 44824 3556
rect 44876 3584 44882 3596
rect 45002 3584 45008 3596
rect 44876 3556 45008 3584
rect 44876 3544 44882 3556
rect 45002 3544 45008 3556
rect 45060 3544 45066 3596
rect 45278 3544 45284 3596
rect 45336 3544 45342 3596
rect 55398 3544 55404 3596
rect 55456 3584 55462 3596
rect 56410 3584 56416 3596
rect 55456 3556 56416 3584
rect 55456 3544 55462 3556
rect 56410 3544 56416 3556
rect 56468 3584 56474 3596
rect 57164 3584 57192 3683
rect 57790 3612 57796 3664
rect 57848 3652 57854 3664
rect 58912 3661 58940 3692
rect 59354 3680 59360 3692
rect 59412 3680 59418 3732
rect 72602 3680 72608 3732
rect 72660 3680 72666 3732
rect 58897 3655 58955 3661
rect 58897 3652 58909 3655
rect 57848 3624 58909 3652
rect 57848 3612 57854 3624
rect 58897 3621 58909 3624
rect 58943 3621 58955 3655
rect 58897 3615 58955 3621
rect 68922 3612 68928 3664
rect 68980 3652 68986 3664
rect 77662 3652 77668 3664
rect 68980 3624 77668 3652
rect 68980 3612 68986 3624
rect 77662 3612 77668 3624
rect 77720 3612 77726 3664
rect 57698 3584 57704 3596
rect 56468 3556 56640 3584
rect 57164 3556 57704 3584
rect 56468 3544 56474 3556
rect 31602 3488 31800 3516
rect 31846 3476 31852 3528
rect 31904 3516 31910 3528
rect 32125 3519 32183 3525
rect 32125 3516 32137 3519
rect 31904 3488 32137 3516
rect 31904 3476 31910 3488
rect 32125 3485 32137 3488
rect 32171 3485 32183 3519
rect 44269 3519 44327 3525
rect 44269 3516 44281 3519
rect 32125 3479 32183 3485
rect 42812 3488 44281 3516
rect 38930 3408 38936 3460
rect 38988 3408 38994 3460
rect 41414 3408 41420 3460
rect 41472 3408 41478 3460
rect 42702 3448 42708 3460
rect 42642 3420 42708 3448
rect 42702 3408 42708 3420
rect 42760 3408 42766 3460
rect 31938 3340 31944 3392
rect 31996 3340 32002 3392
rect 38948 3380 38976 3408
rect 42812 3380 42840 3488
rect 44269 3485 44281 3488
rect 44315 3516 44327 3519
rect 44910 3516 44916 3528
rect 44315 3488 44916 3516
rect 44315 3485 44327 3488
rect 44269 3479 44327 3485
rect 44910 3476 44916 3488
rect 44968 3476 44974 3528
rect 50617 3519 50675 3525
rect 50617 3485 50629 3519
rect 50663 3516 50675 3519
rect 51261 3519 51319 3525
rect 51261 3516 51273 3519
rect 50663 3488 51273 3516
rect 50663 3485 50675 3488
rect 50617 3479 50675 3485
rect 51261 3485 51273 3488
rect 51307 3516 51319 3519
rect 52914 3516 52920 3528
rect 51307 3488 52920 3516
rect 51307 3485 51319 3488
rect 51261 3479 51319 3485
rect 52914 3476 52920 3488
rect 52972 3476 52978 3528
rect 54294 3476 54300 3528
rect 54352 3516 54358 3528
rect 55309 3519 55367 3525
rect 55309 3516 55321 3519
rect 54352 3488 55321 3516
rect 54352 3476 54358 3488
rect 55309 3485 55321 3488
rect 55355 3485 55367 3519
rect 55309 3479 55367 3485
rect 55490 3476 55496 3528
rect 55548 3516 55554 3528
rect 56612 3525 56640 3556
rect 57698 3544 57704 3556
rect 57756 3584 57762 3596
rect 59081 3587 59139 3593
rect 59081 3584 59093 3587
rect 57756 3556 58388 3584
rect 57756 3544 57762 3556
rect 56321 3519 56379 3525
rect 56321 3516 56333 3519
rect 55548 3488 56333 3516
rect 55548 3476 55554 3488
rect 56321 3485 56333 3488
rect 56367 3485 56379 3519
rect 56321 3479 56379 3485
rect 56505 3519 56563 3525
rect 56505 3485 56517 3519
rect 56551 3485 56563 3519
rect 56505 3479 56563 3485
rect 56597 3519 56655 3525
rect 56597 3485 56609 3519
rect 56643 3485 56655 3519
rect 56597 3479 56655 3485
rect 57517 3519 57575 3525
rect 57517 3485 57529 3519
rect 57563 3516 57575 3519
rect 57609 3519 57667 3525
rect 57609 3516 57621 3519
rect 57563 3488 57621 3516
rect 57563 3485 57575 3488
rect 57517 3479 57575 3485
rect 57609 3485 57621 3488
rect 57655 3485 57667 3519
rect 57609 3479 57667 3485
rect 43622 3408 43628 3460
rect 43680 3408 43686 3460
rect 43809 3451 43867 3457
rect 43809 3417 43821 3451
rect 43855 3448 43867 3451
rect 43898 3448 43904 3460
rect 43855 3420 43904 3448
rect 43855 3417 43867 3420
rect 43809 3411 43867 3417
rect 43898 3408 43904 3420
rect 43956 3408 43962 3460
rect 44453 3451 44511 3457
rect 44453 3417 44465 3451
rect 44499 3448 44511 3451
rect 44542 3448 44548 3460
rect 44499 3420 44548 3448
rect 44499 3417 44511 3420
rect 44453 3411 44511 3417
rect 44542 3408 44548 3420
rect 44600 3408 44606 3460
rect 47762 3448 47768 3460
rect 46506 3420 47768 3448
rect 47762 3408 47768 3420
rect 47820 3408 47826 3460
rect 50338 3408 50344 3460
rect 50396 3448 50402 3460
rect 51169 3451 51227 3457
rect 51169 3448 51181 3451
rect 50396 3420 51181 3448
rect 50396 3408 50402 3420
rect 51169 3417 51181 3420
rect 51215 3417 51227 3451
rect 51169 3411 51227 3417
rect 55953 3451 56011 3457
rect 55953 3417 55965 3451
rect 55999 3448 56011 3451
rect 56520 3448 56548 3479
rect 58158 3476 58164 3528
rect 58216 3476 58222 3528
rect 58250 3448 58256 3460
rect 55999 3420 58256 3448
rect 55999 3417 56011 3420
rect 55953 3411 56011 3417
rect 58250 3408 58256 3420
rect 58308 3408 58314 3460
rect 58360 3448 58388 3556
rect 58544 3556 59093 3584
rect 58544 3525 58572 3556
rect 59081 3553 59093 3556
rect 59127 3553 59139 3587
rect 59081 3547 59139 3553
rect 72513 3587 72571 3593
rect 72513 3553 72525 3587
rect 72559 3584 72571 3587
rect 74442 3584 74448 3596
rect 72559 3556 74448 3584
rect 72559 3553 72571 3556
rect 72513 3547 72571 3553
rect 74442 3544 74448 3556
rect 74500 3544 74506 3596
rect 58529 3519 58587 3525
rect 58529 3485 58541 3519
rect 58575 3485 58587 3519
rect 58529 3479 58587 3485
rect 58986 3476 58992 3528
rect 59044 3476 59050 3528
rect 68462 3476 68468 3528
rect 68520 3516 68526 3528
rect 72329 3519 72387 3525
rect 72329 3516 72341 3519
rect 68520 3488 72341 3516
rect 68520 3476 68526 3488
rect 72329 3485 72341 3488
rect 72375 3485 72387 3519
rect 72329 3479 72387 3485
rect 72418 3476 72424 3528
rect 72476 3516 72482 3528
rect 72697 3519 72755 3525
rect 72697 3516 72709 3519
rect 72476 3488 72709 3516
rect 72476 3476 72482 3488
rect 72697 3485 72709 3488
rect 72743 3516 72755 3519
rect 72973 3519 73031 3525
rect 72973 3516 72985 3519
rect 72743 3488 72985 3516
rect 72743 3485 72755 3488
rect 72697 3479 72755 3485
rect 72973 3485 72985 3488
rect 73019 3516 73031 3519
rect 73522 3516 73528 3528
rect 73019 3488 73528 3516
rect 73019 3485 73031 3488
rect 72973 3479 73031 3485
rect 73522 3476 73528 3488
rect 73580 3516 73586 3528
rect 76190 3516 76196 3528
rect 73580 3488 76196 3516
rect 73580 3476 73586 3488
rect 76190 3476 76196 3488
rect 76248 3476 76254 3528
rect 58621 3451 58679 3457
rect 58360 3420 58572 3448
rect 38948 3352 42840 3380
rect 50798 3340 50804 3392
rect 50856 3340 50862 3392
rect 50982 3389 50988 3392
rect 50969 3383 50988 3389
rect 50969 3349 50981 3383
rect 50969 3343 50988 3349
rect 50982 3340 50988 3343
rect 51040 3340 51046 3392
rect 56778 3340 56784 3392
rect 56836 3340 56842 3392
rect 56962 3340 56968 3392
rect 57020 3340 57026 3392
rect 57149 3383 57207 3389
rect 57149 3349 57161 3383
rect 57195 3380 57207 3383
rect 57790 3380 57796 3392
rect 57195 3352 57796 3380
rect 57195 3349 57207 3352
rect 57149 3343 57207 3349
rect 57790 3340 57796 3352
rect 57848 3340 57854 3392
rect 58345 3383 58403 3389
rect 58345 3349 58357 3383
rect 58391 3380 58403 3383
rect 58434 3380 58440 3392
rect 58391 3352 58440 3380
rect 58391 3349 58403 3352
rect 58345 3343 58403 3349
rect 58434 3340 58440 3352
rect 58492 3340 58498 3392
rect 58544 3380 58572 3420
rect 58621 3417 58633 3451
rect 58667 3448 58679 3451
rect 59541 3451 59599 3457
rect 59541 3448 59553 3451
rect 58667 3420 58848 3448
rect 58667 3417 58679 3420
rect 58621 3411 58679 3417
rect 58713 3383 58771 3389
rect 58713 3380 58725 3383
rect 58544 3352 58725 3380
rect 58713 3349 58725 3352
rect 58759 3349 58771 3383
rect 58820 3380 58848 3420
rect 59188 3420 59553 3448
rect 59188 3380 59216 3420
rect 59541 3417 59553 3420
rect 59587 3448 59599 3451
rect 59587 3420 72464 3448
rect 59587 3417 59599 3420
rect 59541 3411 59599 3417
rect 58820 3352 59216 3380
rect 58713 3343 58771 3349
rect 72142 3340 72148 3392
rect 72200 3340 72206 3392
rect 72436 3380 72464 3420
rect 72510 3408 72516 3460
rect 72568 3448 72574 3460
rect 72605 3451 72663 3457
rect 72605 3448 72617 3451
rect 72568 3420 72617 3448
rect 72568 3408 72574 3420
rect 72605 3417 72617 3420
rect 72651 3417 72663 3451
rect 78122 3448 78128 3460
rect 72605 3411 72663 3417
rect 72712 3420 78128 3448
rect 72712 3380 72740 3420
rect 78122 3408 78128 3420
rect 78180 3408 78186 3460
rect 72436 3352 72740 3380
rect 72878 3340 72884 3392
rect 72936 3340 72942 3392
rect 73062 3340 73068 3392
rect 73120 3380 73126 3392
rect 77754 3380 77760 3392
rect 73120 3352 77760 3380
rect 73120 3340 73126 3352
rect 77754 3340 77760 3352
rect 77812 3340 77818 3392
rect 77938 3340 77944 3392
rect 77996 3380 78002 3392
rect 78033 3383 78091 3389
rect 78033 3380 78045 3383
rect 77996 3352 78045 3380
rect 77996 3340 78002 3352
rect 78033 3349 78045 3352
rect 78079 3349 78091 3383
rect 78033 3343 78091 3349
rect 78490 3340 78496 3392
rect 78548 3340 78554 3392
rect 1104 3290 78844 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 66314 3290
rect 66366 3238 66378 3290
rect 66430 3238 66442 3290
rect 66494 3238 66506 3290
rect 66558 3238 66570 3290
rect 66622 3238 78844 3290
rect 1104 3216 78844 3238
rect 31846 3136 31852 3188
rect 31904 3136 31910 3188
rect 35986 3136 35992 3188
rect 36044 3176 36050 3188
rect 36044 3148 37964 3176
rect 36044 3136 36050 3148
rect 36004 3108 36032 3136
rect 35360 3080 36032 3108
rect 31938 3000 31944 3052
rect 31996 3040 32002 3052
rect 35360 3049 35388 3080
rect 36262 3068 36268 3120
rect 36320 3068 36326 3120
rect 37936 3108 37964 3148
rect 44266 3136 44272 3188
rect 44324 3176 44330 3188
rect 45097 3179 45155 3185
rect 45097 3176 45109 3179
rect 44324 3148 45109 3176
rect 44324 3136 44330 3148
rect 45097 3145 45109 3148
rect 45143 3145 45155 3179
rect 54294 3176 54300 3188
rect 45097 3139 45155 3145
rect 53668 3148 54300 3176
rect 39850 3108 39856 3120
rect 37936 3080 39856 3108
rect 37936 3049 37964 3080
rect 39850 3068 39856 3080
rect 39908 3108 39914 3120
rect 39908 3080 39988 3108
rect 39908 3068 39914 3080
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 31996 3012 32321 3040
rect 31996 3000 32002 3012
rect 32309 3009 32321 3012
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 35345 3043 35403 3049
rect 35345 3009 35357 3043
rect 35391 3009 35403 3043
rect 35345 3003 35403 3009
rect 37921 3043 37979 3049
rect 37921 3009 37933 3043
rect 37967 3009 37979 3043
rect 37921 3003 37979 3009
rect 38188 3043 38246 3049
rect 38188 3009 38200 3043
rect 38234 3040 38246 3043
rect 38654 3040 38660 3052
rect 38234 3012 38660 3040
rect 38234 3009 38246 3012
rect 38188 3003 38246 3009
rect 38654 3000 38660 3012
rect 38712 3000 38718 3052
rect 39960 3049 39988 3080
rect 44910 3068 44916 3120
rect 44968 3108 44974 3120
rect 45005 3111 45063 3117
rect 45005 3108 45017 3111
rect 44968 3080 45017 3108
rect 44968 3068 44974 3080
rect 45005 3077 45017 3080
rect 45051 3077 45063 3111
rect 45005 3071 45063 3077
rect 50798 3068 50804 3120
rect 50856 3117 50862 3120
rect 53668 3117 53696 3148
rect 54294 3136 54300 3148
rect 54352 3136 54358 3188
rect 57885 3179 57943 3185
rect 57885 3176 57897 3179
rect 55784 3148 57897 3176
rect 50856 3108 50868 3117
rect 53653 3111 53711 3117
rect 50856 3080 50901 3108
rect 50856 3071 50868 3080
rect 53653 3077 53665 3111
rect 53699 3077 53711 3111
rect 53653 3071 53711 3077
rect 53837 3111 53895 3117
rect 53837 3077 53849 3111
rect 53883 3108 53895 3111
rect 54018 3108 54024 3120
rect 53883 3080 54024 3108
rect 53883 3077 53895 3080
rect 53837 3071 53895 3077
rect 50856 3068 50862 3071
rect 54018 3068 54024 3080
rect 54076 3068 54082 3120
rect 55490 3108 55496 3120
rect 55338 3080 55496 3108
rect 55490 3068 55496 3080
rect 55548 3068 55554 3120
rect 55784 3117 55812 3148
rect 57885 3145 57897 3148
rect 57931 3145 57943 3179
rect 57885 3139 57943 3145
rect 58250 3136 58256 3188
rect 58308 3136 58314 3188
rect 59357 3179 59415 3185
rect 59357 3145 59369 3179
rect 59403 3145 59415 3179
rect 66165 3179 66223 3185
rect 66165 3176 66177 3179
rect 59357 3139 59415 3145
rect 64846 3148 66177 3176
rect 55769 3111 55827 3117
rect 55769 3077 55781 3111
rect 55815 3077 55827 3111
rect 55769 3071 55827 3077
rect 56778 3068 56784 3120
rect 56836 3108 56842 3120
rect 59372 3108 59400 3139
rect 59909 3111 59967 3117
rect 59909 3108 59921 3111
rect 56836 3080 59124 3108
rect 59372 3080 59921 3108
rect 56836 3068 56842 3080
rect 39393 3043 39451 3049
rect 39393 3009 39405 3043
rect 39439 3009 39451 3043
rect 39393 3003 39451 3009
rect 39945 3043 40003 3049
rect 39945 3009 39957 3043
rect 39991 3009 40003 3043
rect 39945 3003 40003 3009
rect 35621 2975 35679 2981
rect 35621 2941 35633 2975
rect 35667 2972 35679 2975
rect 36170 2972 36176 2984
rect 35667 2944 36176 2972
rect 35667 2941 35679 2944
rect 35621 2935 35679 2941
rect 36170 2932 36176 2944
rect 36228 2932 36234 2984
rect 37090 2932 37096 2984
rect 37148 2932 37154 2984
rect 39301 2907 39359 2913
rect 39301 2873 39313 2907
rect 39347 2904 39359 2907
rect 39408 2904 39436 3003
rect 40034 3000 40040 3052
rect 40092 3040 40098 3052
rect 40201 3043 40259 3049
rect 40201 3040 40213 3043
rect 40092 3012 40213 3040
rect 40092 3000 40098 3012
rect 40201 3009 40213 3012
rect 40247 3009 40259 3043
rect 40201 3003 40259 3009
rect 44174 3000 44180 3052
rect 44232 3040 44238 3052
rect 44554 3043 44612 3049
rect 44554 3040 44566 3043
rect 44232 3012 44566 3040
rect 44232 3000 44238 3012
rect 44554 3009 44566 3012
rect 44600 3009 44612 3043
rect 44554 3003 44612 3009
rect 44818 3000 44824 3052
rect 44876 3000 44882 3052
rect 45554 3000 45560 3052
rect 45612 3040 45618 3052
rect 46201 3043 46259 3049
rect 46201 3040 46213 3043
rect 45612 3012 46213 3040
rect 45612 3000 45618 3012
rect 46201 3009 46213 3012
rect 46247 3040 46259 3043
rect 46845 3043 46903 3049
rect 46845 3040 46857 3043
rect 46247 3012 46857 3040
rect 46247 3009 46259 3012
rect 46201 3003 46259 3009
rect 46845 3009 46857 3012
rect 46891 3040 46903 3043
rect 47581 3043 47639 3049
rect 47581 3040 47593 3043
rect 46891 3012 47593 3040
rect 46891 3009 46903 3012
rect 46845 3003 46903 3009
rect 47581 3009 47593 3012
rect 47627 3040 47639 3043
rect 48777 3043 48835 3049
rect 48777 3040 48789 3043
rect 47627 3012 48789 3040
rect 47627 3009 47639 3012
rect 47581 3003 47639 3009
rect 48777 3009 48789 3012
rect 48823 3040 48835 3043
rect 49421 3043 49479 3049
rect 49421 3040 49433 3043
rect 48823 3012 49433 3040
rect 48823 3009 48835 3012
rect 48777 3003 48835 3009
rect 49421 3009 49433 3012
rect 49467 3040 49479 3043
rect 49467 3012 51028 3040
rect 49467 3009 49479 3012
rect 49421 3003 49479 3009
rect 42061 2975 42119 2981
rect 42061 2972 42073 2975
rect 41340 2944 42073 2972
rect 39482 2904 39488 2916
rect 39347 2876 39488 2904
rect 39347 2873 39359 2876
rect 39301 2867 39359 2873
rect 39482 2864 39488 2876
rect 39540 2864 39546 2916
rect 41340 2913 41368 2944
rect 42061 2941 42073 2944
rect 42107 2972 42119 2975
rect 51000 2972 51028 3012
rect 51074 3000 51080 3052
rect 51132 3000 51138 3052
rect 51353 3043 51411 3049
rect 51353 3009 51365 3043
rect 51399 3040 51411 3043
rect 51442 3040 51448 3052
rect 51399 3012 51448 3040
rect 51399 3009 51411 3012
rect 51353 3003 51411 3009
rect 51368 2972 51396 3003
rect 51442 3000 51448 3012
rect 51500 3000 51506 3052
rect 56137 3043 56195 3049
rect 56137 3009 56149 3043
rect 56183 3009 56195 3043
rect 56137 3003 56195 3009
rect 42107 2944 43668 2972
rect 51000 2944 51396 2972
rect 42107 2941 42119 2944
rect 42061 2935 42119 2941
rect 41325 2907 41383 2913
rect 41325 2873 41337 2907
rect 41371 2873 41383 2907
rect 41325 2867 41383 2873
rect 32493 2839 32551 2845
rect 32493 2805 32505 2839
rect 32539 2836 32551 2839
rect 32950 2836 32956 2848
rect 32539 2808 32956 2836
rect 32539 2805 32551 2808
rect 32493 2799 32551 2805
rect 32950 2796 32956 2808
rect 33008 2796 33014 2848
rect 39390 2796 39396 2848
rect 39448 2836 39454 2848
rect 39577 2839 39635 2845
rect 39577 2836 39589 2839
rect 39448 2808 39589 2836
rect 39448 2796 39454 2808
rect 39577 2805 39589 2808
rect 39623 2805 39635 2839
rect 39577 2799 39635 2805
rect 41414 2796 41420 2848
rect 41472 2796 41478 2848
rect 43346 2796 43352 2848
rect 43404 2796 43410 2848
rect 43441 2839 43499 2845
rect 43441 2805 43453 2839
rect 43487 2836 43499 2839
rect 43530 2836 43536 2848
rect 43487 2808 43536 2836
rect 43487 2805 43499 2808
rect 43441 2799 43499 2805
rect 43530 2796 43536 2808
rect 43588 2796 43594 2848
rect 43640 2836 43668 2944
rect 56042 2932 56048 2984
rect 56100 2932 56106 2984
rect 49605 2907 49663 2913
rect 49605 2873 49617 2907
rect 49651 2904 49663 2907
rect 49786 2904 49792 2916
rect 49651 2876 49792 2904
rect 49651 2873 49663 2876
rect 49605 2867 49663 2873
rect 49786 2864 49792 2876
rect 49844 2864 49850 2916
rect 45002 2836 45008 2848
rect 43640 2808 45008 2836
rect 45002 2796 45008 2808
rect 45060 2796 45066 2848
rect 45741 2839 45799 2845
rect 45741 2805 45753 2839
rect 45787 2836 45799 2839
rect 45830 2836 45836 2848
rect 45787 2808 45836 2836
rect 45787 2805 45799 2808
rect 45741 2799 45799 2805
rect 45830 2796 45836 2808
rect 45888 2796 45894 2848
rect 46385 2839 46443 2845
rect 46385 2805 46397 2839
rect 46431 2836 46443 2839
rect 46474 2836 46480 2848
rect 46431 2808 46480 2836
rect 46431 2805 46443 2808
rect 46385 2799 46443 2805
rect 46474 2796 46480 2808
rect 46532 2796 46538 2848
rect 47029 2839 47087 2845
rect 47029 2805 47041 2839
rect 47075 2836 47087 2839
rect 47118 2836 47124 2848
rect 47075 2808 47124 2836
rect 47075 2805 47087 2808
rect 47029 2799 47087 2805
rect 47118 2796 47124 2808
rect 47176 2796 47182 2848
rect 47762 2796 47768 2848
rect 47820 2796 47826 2848
rect 48961 2839 49019 2845
rect 48961 2805 48973 2839
rect 49007 2836 49019 2839
rect 49050 2836 49056 2848
rect 49007 2808 49056 2836
rect 49007 2805 49019 2808
rect 48961 2799 49019 2805
rect 49050 2796 49056 2808
rect 49108 2796 49114 2848
rect 49694 2796 49700 2848
rect 49752 2796 49758 2848
rect 51169 2839 51227 2845
rect 51169 2805 51181 2839
rect 51215 2836 51227 2839
rect 51258 2836 51264 2848
rect 51215 2808 51264 2836
rect 51215 2805 51227 2808
rect 51169 2799 51227 2805
rect 51258 2796 51264 2808
rect 51316 2796 51322 2848
rect 51626 2796 51632 2848
rect 51684 2796 51690 2848
rect 53469 2839 53527 2845
rect 53469 2805 53481 2839
rect 53515 2836 53527 2839
rect 53558 2836 53564 2848
rect 53515 2808 53564 2836
rect 53515 2805 53527 2808
rect 53469 2799 53527 2805
rect 53558 2796 53564 2808
rect 53616 2796 53622 2848
rect 54110 2796 54116 2848
rect 54168 2796 54174 2848
rect 55306 2796 55312 2848
rect 55364 2836 55370 2848
rect 56152 2836 56180 3003
rect 56318 3000 56324 3052
rect 56376 3040 56382 3052
rect 56413 3043 56471 3049
rect 56413 3040 56425 3043
rect 56376 3012 56425 3040
rect 56376 3000 56382 3012
rect 56413 3009 56425 3012
rect 56459 3040 56471 3043
rect 56689 3043 56747 3049
rect 56689 3040 56701 3043
rect 56459 3012 56701 3040
rect 56459 3009 56471 3012
rect 56413 3003 56471 3009
rect 56689 3009 56701 3012
rect 56735 3009 56747 3043
rect 56689 3003 56747 3009
rect 57701 3043 57759 3049
rect 57701 3009 57713 3043
rect 57747 3040 57759 3043
rect 57790 3040 57796 3052
rect 57747 3012 57796 3040
rect 57747 3009 57759 3012
rect 57701 3003 57759 3009
rect 57790 3000 57796 3012
rect 57848 3000 57854 3052
rect 58710 3000 58716 3052
rect 58768 3000 58774 3052
rect 58989 3043 59047 3049
rect 58989 3009 59001 3043
rect 59035 3009 59047 3043
rect 59096 3040 59124 3080
rect 59909 3077 59921 3080
rect 59955 3077 59967 3111
rect 64846 3108 64874 3148
rect 66165 3145 66177 3148
rect 66211 3145 66223 3179
rect 68373 3179 68431 3185
rect 68373 3176 68385 3179
rect 66165 3139 66223 3145
rect 66272 3148 68385 3176
rect 66272 3108 66300 3148
rect 68373 3145 68385 3148
rect 68419 3176 68431 3179
rect 68922 3176 68928 3188
rect 68419 3148 68928 3176
rect 68419 3145 68431 3148
rect 68373 3139 68431 3145
rect 68922 3136 68928 3148
rect 68980 3136 68986 3188
rect 72418 3176 72424 3188
rect 69124 3148 72424 3176
rect 59909 3071 59967 3077
rect 60706 3080 64874 3108
rect 66180 3080 66300 3108
rect 59541 3043 59599 3049
rect 59541 3040 59553 3043
rect 59096 3012 59553 3040
rect 58989 3003 59047 3009
rect 59541 3009 59553 3012
rect 59587 3009 59599 3043
rect 59541 3003 59599 3009
rect 56229 2975 56287 2981
rect 56229 2941 56241 2975
rect 56275 2972 56287 2975
rect 56594 2972 56600 2984
rect 56275 2944 56600 2972
rect 56275 2941 56287 2944
rect 56229 2935 56287 2941
rect 56594 2932 56600 2944
rect 56652 2932 56658 2984
rect 58342 2932 58348 2984
rect 58400 2932 58406 2984
rect 58434 2932 58440 2984
rect 58492 2932 58498 2984
rect 58802 2932 58808 2984
rect 58860 2932 58866 2984
rect 59004 2972 59032 3003
rect 59814 3000 59820 3052
rect 59872 3000 59878 3052
rect 60185 3043 60243 3049
rect 60185 3009 60197 3043
rect 60231 3040 60243 3043
rect 60706 3040 60734 3080
rect 60231 3012 60734 3040
rect 61565 3043 61623 3049
rect 60231 3009 60243 3012
rect 60185 3003 60243 3009
rect 61565 3009 61577 3043
rect 61611 3040 61623 3043
rect 61933 3043 61991 3049
rect 61933 3040 61945 3043
rect 61611 3012 61945 3040
rect 61611 3009 61623 3012
rect 61565 3003 61623 3009
rect 61933 3009 61945 3012
rect 61979 3040 61991 3043
rect 62209 3043 62267 3049
rect 62209 3040 62221 3043
rect 61979 3012 62221 3040
rect 61979 3009 61991 3012
rect 61933 3003 61991 3009
rect 62209 3009 62221 3012
rect 62255 3040 62267 3043
rect 62577 3043 62635 3049
rect 62577 3040 62589 3043
rect 62255 3012 62589 3040
rect 62255 3009 62267 3012
rect 62209 3003 62267 3009
rect 62577 3009 62589 3012
rect 62623 3040 62635 3043
rect 63037 3043 63095 3049
rect 63037 3040 63049 3043
rect 62623 3012 63049 3040
rect 62623 3009 62635 3012
rect 62577 3003 62635 3009
rect 63037 3009 63049 3012
rect 63083 3040 63095 3043
rect 63405 3043 63463 3049
rect 63405 3040 63417 3043
rect 63083 3012 63417 3040
rect 63083 3009 63095 3012
rect 63037 3003 63095 3009
rect 63405 3009 63417 3012
rect 63451 3040 63463 3043
rect 63497 3043 63555 3049
rect 63497 3040 63509 3043
rect 63451 3012 63509 3040
rect 63451 3009 63463 3012
rect 63405 3003 63463 3009
rect 63497 3009 63509 3012
rect 63543 3040 63555 3043
rect 63865 3043 63923 3049
rect 63865 3040 63877 3043
rect 63543 3012 63877 3040
rect 63543 3009 63555 3012
rect 63497 3003 63555 3009
rect 63865 3009 63877 3012
rect 63911 3040 63923 3043
rect 64141 3043 64199 3049
rect 64141 3040 64153 3043
rect 63911 3012 64153 3040
rect 63911 3009 63923 3012
rect 63865 3003 63923 3009
rect 64141 3009 64153 3012
rect 64187 3040 64199 3043
rect 64509 3043 64567 3049
rect 64509 3040 64521 3043
rect 64187 3012 64521 3040
rect 64187 3009 64199 3012
rect 64141 3003 64199 3009
rect 64509 3009 64521 3012
rect 64555 3040 64567 3043
rect 66180 3040 66208 3080
rect 66438 3068 66444 3120
rect 66496 3108 66502 3120
rect 69124 3117 69152 3148
rect 72418 3136 72424 3148
rect 72476 3136 72482 3188
rect 72510 3136 72516 3188
rect 72568 3136 72574 3188
rect 72602 3136 72608 3188
rect 72660 3136 72666 3188
rect 73522 3136 73528 3188
rect 73580 3136 73586 3188
rect 78125 3179 78183 3185
rect 78125 3176 78137 3179
rect 74280 3148 78137 3176
rect 66625 3111 66683 3117
rect 66625 3108 66637 3111
rect 66496 3080 66637 3108
rect 66496 3068 66502 3080
rect 66625 3077 66637 3080
rect 66671 3077 66683 3111
rect 69109 3111 69167 3117
rect 69109 3108 69121 3111
rect 66625 3071 66683 3077
rect 68204 3080 69121 3108
rect 68204 3052 68232 3080
rect 69109 3077 69121 3080
rect 69155 3077 69167 3111
rect 69109 3071 69167 3077
rect 71041 3111 71099 3117
rect 71041 3077 71053 3111
rect 71087 3108 71099 3111
rect 72053 3111 72111 3117
rect 72053 3108 72065 3111
rect 71087 3080 72065 3108
rect 71087 3077 71099 3080
rect 71041 3071 71099 3077
rect 72053 3077 72065 3080
rect 72099 3077 72111 3111
rect 72053 3071 72111 3077
rect 72142 3068 72148 3120
rect 72200 3108 72206 3120
rect 74280 3117 74308 3148
rect 78125 3145 78137 3148
rect 78171 3145 78183 3179
rect 78125 3139 78183 3145
rect 73433 3111 73491 3117
rect 73433 3108 73445 3111
rect 72200 3080 73445 3108
rect 72200 3068 72206 3080
rect 73433 3077 73445 3080
rect 73479 3077 73491 3111
rect 73433 3071 73491 3077
rect 74261 3111 74319 3117
rect 74261 3077 74273 3111
rect 74307 3077 74319 3111
rect 74261 3071 74319 3077
rect 74353 3111 74411 3117
rect 74353 3077 74365 3111
rect 74399 3108 74411 3111
rect 77386 3108 77392 3120
rect 74399 3080 77392 3108
rect 74399 3077 74411 3080
rect 74353 3071 74411 3077
rect 77386 3068 77392 3080
rect 77444 3068 77450 3120
rect 64555 3012 66208 3040
rect 66349 3043 66407 3049
rect 64555 3009 64567 3012
rect 64509 3003 64567 3009
rect 66349 3009 66361 3043
rect 66395 3040 66407 3043
rect 66395 3012 68140 3040
rect 66395 3009 66407 3012
rect 66349 3003 66407 3009
rect 59630 2972 59636 2984
rect 59004 2944 59636 2972
rect 59630 2932 59636 2944
rect 59688 2932 59694 2984
rect 59722 2932 59728 2984
rect 59780 2932 59786 2984
rect 59998 2932 60004 2984
rect 60056 2932 60062 2984
rect 66530 2932 66536 2984
rect 66588 2932 66594 2984
rect 68112 2972 68140 3012
rect 68186 3000 68192 3052
rect 68244 3000 68250 3052
rect 68741 3043 68799 3049
rect 68741 3009 68753 3043
rect 68787 3040 68799 3043
rect 68922 3040 68928 3052
rect 68787 3012 68928 3040
rect 68787 3009 68799 3012
rect 68741 3003 68799 3009
rect 68922 3000 68928 3012
rect 68980 3000 68986 3052
rect 69014 3000 69020 3052
rect 69072 3040 69078 3052
rect 70949 3043 71007 3049
rect 70949 3040 70961 3043
rect 69072 3012 70961 3040
rect 69072 3000 69078 3012
rect 70949 3009 70961 3012
rect 70995 3009 71007 3043
rect 70949 3003 71007 3009
rect 71130 3000 71136 3052
rect 71188 3000 71194 3052
rect 71222 3000 71228 3052
rect 71280 3040 71286 3052
rect 72329 3043 72387 3049
rect 72329 3040 72341 3043
rect 71280 3012 72341 3040
rect 71280 3000 71286 3012
rect 72329 3009 72341 3012
rect 72375 3009 72387 3043
rect 72329 3003 72387 3009
rect 72418 3000 72424 3052
rect 72476 3040 72482 3052
rect 72789 3043 72847 3049
rect 72789 3040 72801 3043
rect 72476 3012 72801 3040
rect 72476 3000 72482 3012
rect 72789 3009 72801 3012
rect 72835 3009 72847 3043
rect 73065 3043 73123 3049
rect 73065 3040 73077 3043
rect 72789 3003 72847 3009
rect 72896 3012 73077 3040
rect 69750 2972 69756 2984
rect 68112 2944 69756 2972
rect 69750 2932 69756 2944
rect 69808 2932 69814 2984
rect 72234 2932 72240 2984
rect 72292 2932 72298 2984
rect 72510 2932 72516 2984
rect 72568 2972 72574 2984
rect 72896 2972 72924 3012
rect 73065 3009 73077 3012
rect 73111 3009 73123 3043
rect 73065 3003 73123 3009
rect 73982 3000 73988 3052
rect 74040 3040 74046 3052
rect 74077 3043 74135 3049
rect 74077 3040 74089 3043
rect 74040 3012 74089 3040
rect 74040 3000 74046 3012
rect 74077 3009 74089 3012
rect 74123 3009 74135 3043
rect 74077 3003 74135 3009
rect 74166 3000 74172 3052
rect 74224 3000 74230 3052
rect 76190 3000 76196 3052
rect 76248 3040 76254 3052
rect 77846 3049 77852 3052
rect 76377 3043 76435 3049
rect 76377 3040 76389 3043
rect 76248 3012 76389 3040
rect 76248 3000 76254 3012
rect 76377 3009 76389 3012
rect 76423 3040 76435 3043
rect 77665 3043 77723 3049
rect 77665 3040 77677 3043
rect 76423 3012 77677 3040
rect 76423 3009 76435 3012
rect 76377 3003 76435 3009
rect 77665 3009 77677 3012
rect 77711 3040 77723 3043
rect 77841 3040 77852 3049
rect 77711 3012 77852 3040
rect 77711 3009 77723 3012
rect 77665 3003 77723 3009
rect 77841 3003 77852 3012
rect 77846 3000 77852 3003
rect 77904 3000 77910 3052
rect 78309 3043 78367 3049
rect 78309 3009 78321 3043
rect 78355 3040 78367 3043
rect 78490 3040 78496 3052
rect 78355 3012 78496 3040
rect 78355 3009 78367 3012
rect 78309 3003 78367 3009
rect 78490 3000 78496 3012
rect 78548 3040 78554 3052
rect 79226 3040 79232 3052
rect 78548 3012 79232 3040
rect 78548 3000 78554 3012
rect 79226 3000 79232 3012
rect 79284 3000 79290 3052
rect 72568 2944 72924 2972
rect 72973 2975 73031 2981
rect 72568 2932 72574 2944
rect 72973 2941 72985 2975
rect 73019 2972 73031 2975
rect 73019 2944 74212 2972
rect 73019 2941 73031 2944
rect 72973 2935 73031 2941
rect 59173 2907 59231 2913
rect 56612 2876 58940 2904
rect 56612 2845 56640 2876
rect 55364 2808 56180 2836
rect 56597 2839 56655 2845
rect 55364 2796 55370 2808
rect 56597 2805 56609 2839
rect 56643 2805 56655 2839
rect 56597 2799 56655 2805
rect 57422 2796 57428 2848
rect 57480 2796 57486 2848
rect 57974 2796 57980 2848
rect 58032 2836 58038 2848
rect 58713 2839 58771 2845
rect 58713 2836 58725 2839
rect 58032 2808 58725 2836
rect 58032 2796 58038 2808
rect 58713 2805 58725 2808
rect 58759 2805 58771 2839
rect 58912 2836 58940 2876
rect 59173 2873 59185 2907
rect 59219 2904 59231 2907
rect 60369 2907 60427 2913
rect 59219 2876 59952 2904
rect 59219 2873 59231 2876
rect 59173 2867 59231 2873
rect 59924 2845 59952 2876
rect 60369 2873 60381 2907
rect 60415 2904 60427 2907
rect 68462 2904 68468 2916
rect 60415 2876 68468 2904
rect 60415 2873 60427 2876
rect 60369 2867 60427 2873
rect 68462 2864 68468 2876
rect 68520 2864 68526 2916
rect 74184 2904 74212 2944
rect 74442 2932 74448 2984
rect 74500 2972 74506 2984
rect 74537 2975 74595 2981
rect 74537 2972 74549 2975
rect 74500 2944 74549 2972
rect 74500 2932 74506 2944
rect 74537 2941 74549 2944
rect 74583 2941 74595 2975
rect 74537 2935 74595 2941
rect 74258 2904 74264 2916
rect 73080 2876 73660 2904
rect 74184 2876 74264 2904
rect 59541 2839 59599 2845
rect 59541 2836 59553 2839
rect 58912 2808 59553 2836
rect 58713 2799 58771 2805
rect 59541 2805 59553 2808
rect 59587 2805 59599 2839
rect 59541 2799 59599 2805
rect 59909 2839 59967 2845
rect 59909 2805 59921 2839
rect 59955 2805 59967 2839
rect 59909 2799 59967 2805
rect 61746 2796 61752 2848
rect 61804 2796 61810 2848
rect 62390 2796 62396 2848
rect 62448 2796 62454 2848
rect 63218 2796 63224 2848
rect 63276 2796 63282 2848
rect 63678 2796 63684 2848
rect 63736 2796 63742 2848
rect 64322 2796 64328 2848
rect 64380 2796 64386 2848
rect 65978 2796 65984 2848
rect 66036 2836 66042 2848
rect 66438 2836 66444 2848
rect 66036 2808 66444 2836
rect 66036 2796 66042 2808
rect 66438 2796 66444 2808
rect 66496 2796 66502 2848
rect 66625 2839 66683 2845
rect 66625 2805 66637 2839
rect 66671 2836 66683 2839
rect 67634 2836 67640 2848
rect 66671 2808 67640 2836
rect 66671 2805 66683 2808
rect 66625 2799 66683 2805
rect 67634 2796 67640 2808
rect 67692 2796 67698 2848
rect 68557 2839 68615 2845
rect 68557 2805 68569 2839
rect 68603 2836 68615 2839
rect 68646 2836 68652 2848
rect 68603 2808 68652 2836
rect 68603 2805 68615 2808
rect 68557 2799 68615 2805
rect 68646 2796 68652 2808
rect 68704 2796 68710 2848
rect 72329 2839 72387 2845
rect 72329 2805 72341 2839
rect 72375 2836 72387 2839
rect 72970 2836 72976 2848
rect 72375 2808 72976 2836
rect 72375 2805 72387 2808
rect 72329 2799 72387 2805
rect 72970 2796 72976 2808
rect 73028 2796 73034 2848
rect 73080 2845 73108 2876
rect 73065 2839 73123 2845
rect 73065 2805 73077 2839
rect 73111 2805 73123 2839
rect 73632 2836 73660 2876
rect 74258 2864 74264 2876
rect 74316 2864 74322 2916
rect 76098 2836 76104 2848
rect 73632 2808 76104 2836
rect 73065 2799 73123 2805
rect 76098 2796 76104 2808
rect 76156 2796 76162 2848
rect 76561 2839 76619 2845
rect 76561 2805 76573 2839
rect 76607 2836 76619 2839
rect 76742 2836 76748 2848
rect 76607 2808 76748 2836
rect 76607 2805 76619 2808
rect 76561 2799 76619 2805
rect 76742 2796 76748 2808
rect 76800 2796 76806 2848
rect 78030 2796 78036 2848
rect 78088 2796 78094 2848
rect 1104 2746 78844 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 78844 2746
rect 1104 2672 78844 2694
rect 38654 2592 38660 2644
rect 38712 2592 38718 2644
rect 39945 2635 40003 2641
rect 39945 2601 39957 2635
rect 39991 2632 40003 2635
rect 40034 2632 40040 2644
rect 39991 2604 40040 2632
rect 39991 2601 40003 2604
rect 39945 2595 40003 2601
rect 40034 2592 40040 2604
rect 40092 2592 40098 2644
rect 43717 2635 43775 2641
rect 43717 2601 43729 2635
rect 43763 2632 43775 2635
rect 44174 2632 44180 2644
rect 43763 2604 44180 2632
rect 43763 2601 43775 2604
rect 43717 2595 43775 2601
rect 44174 2592 44180 2604
rect 44232 2592 44238 2644
rect 45554 2632 45560 2644
rect 44836 2604 45560 2632
rect 43162 2524 43168 2576
rect 43220 2564 43226 2576
rect 44637 2567 44695 2573
rect 44637 2564 44649 2567
rect 43220 2536 44649 2564
rect 43220 2524 43226 2536
rect 44637 2533 44649 2536
rect 44683 2533 44695 2567
rect 44637 2527 44695 2533
rect 39482 2456 39488 2508
rect 39540 2456 39546 2508
rect 40678 2496 40684 2508
rect 40144 2468 40684 2496
rect 32950 2388 32956 2440
rect 33008 2388 33014 2440
rect 38010 2388 38016 2440
rect 38068 2388 38074 2440
rect 38194 2388 38200 2440
rect 38252 2388 38258 2440
rect 40144 2437 40172 2468
rect 40678 2456 40684 2468
rect 40736 2456 40742 2508
rect 43530 2496 43536 2508
rect 42904 2468 43536 2496
rect 38289 2431 38347 2437
rect 38289 2397 38301 2431
rect 38335 2397 38347 2431
rect 38289 2391 38347 2397
rect 38381 2431 38439 2437
rect 38381 2397 38393 2431
rect 38427 2428 38439 2431
rect 38933 2431 38991 2437
rect 38933 2428 38945 2431
rect 38427 2400 38945 2428
rect 38427 2397 38439 2400
rect 38381 2391 38439 2397
rect 38933 2397 38945 2400
rect 38979 2397 38991 2431
rect 38933 2391 38991 2397
rect 40129 2431 40187 2437
rect 40129 2397 40141 2431
rect 40175 2397 40187 2431
rect 40129 2391 40187 2397
rect 40405 2431 40463 2437
rect 40405 2397 40417 2431
rect 40451 2397 40463 2431
rect 40405 2391 40463 2397
rect 40589 2431 40647 2437
rect 40589 2397 40601 2431
rect 40635 2428 40647 2431
rect 41414 2428 41420 2440
rect 40635 2400 41420 2428
rect 40635 2397 40647 2400
rect 40589 2391 40647 2397
rect 38304 2360 38332 2391
rect 38841 2363 38899 2369
rect 38841 2360 38853 2363
rect 38304 2332 38853 2360
rect 38841 2329 38853 2332
rect 38887 2360 38899 2363
rect 40420 2360 40448 2391
rect 41414 2388 41420 2400
rect 41472 2388 41478 2440
rect 42904 2437 42932 2468
rect 43530 2456 43536 2468
rect 43588 2496 43594 2508
rect 44361 2499 44419 2505
rect 44361 2496 44373 2499
rect 43588 2468 44373 2496
rect 43588 2456 43594 2468
rect 44361 2465 44373 2468
rect 44407 2465 44419 2499
rect 44361 2459 44419 2465
rect 42889 2431 42947 2437
rect 42889 2397 42901 2431
rect 42935 2397 42947 2431
rect 42889 2391 42947 2397
rect 43070 2388 43076 2440
rect 43128 2388 43134 2440
rect 43254 2388 43260 2440
rect 43312 2388 43318 2440
rect 43346 2388 43352 2440
rect 43404 2388 43410 2440
rect 44836 2437 44864 2604
rect 45554 2592 45560 2604
rect 45612 2592 45618 2644
rect 50525 2635 50583 2641
rect 50525 2601 50537 2635
rect 50571 2632 50583 2635
rect 50982 2632 50988 2644
rect 50571 2604 50988 2632
rect 50571 2601 50583 2604
rect 50525 2595 50583 2601
rect 50982 2592 50988 2604
rect 51040 2592 51046 2644
rect 54113 2635 54171 2641
rect 54113 2601 54125 2635
rect 54159 2632 54171 2635
rect 54573 2635 54631 2641
rect 54573 2632 54585 2635
rect 54159 2604 54585 2632
rect 54159 2601 54171 2604
rect 54113 2595 54171 2601
rect 54573 2601 54585 2604
rect 54619 2601 54631 2635
rect 54573 2595 54631 2601
rect 54662 2592 54668 2644
rect 54720 2632 54726 2644
rect 57974 2632 57980 2644
rect 54720 2604 57980 2632
rect 54720 2592 54726 2604
rect 57974 2592 57980 2604
rect 58032 2592 58038 2644
rect 58437 2635 58495 2641
rect 58437 2601 58449 2635
rect 58483 2632 58495 2635
rect 58710 2632 58716 2644
rect 58483 2604 58716 2632
rect 58483 2601 58495 2604
rect 58437 2595 58495 2601
rect 58710 2592 58716 2604
rect 58768 2592 58774 2644
rect 59814 2592 59820 2644
rect 59872 2632 59878 2644
rect 60001 2635 60059 2641
rect 60001 2632 60013 2635
rect 59872 2604 60013 2632
rect 59872 2592 59878 2604
rect 60001 2601 60013 2604
rect 60047 2601 60059 2635
rect 60001 2595 60059 2601
rect 66530 2592 66536 2644
rect 66588 2632 66594 2644
rect 66625 2635 66683 2641
rect 66625 2632 66637 2635
rect 66588 2604 66637 2632
rect 66588 2592 66594 2604
rect 66625 2601 66637 2604
rect 66671 2601 66683 2635
rect 66625 2595 66683 2601
rect 67634 2592 67640 2644
rect 67692 2632 67698 2644
rect 69661 2635 69719 2641
rect 69661 2632 69673 2635
rect 67692 2604 69673 2632
rect 67692 2592 67698 2604
rect 69661 2601 69673 2604
rect 69707 2601 69719 2635
rect 69661 2595 69719 2601
rect 69750 2592 69756 2644
rect 69808 2632 69814 2644
rect 70305 2635 70363 2641
rect 70305 2632 70317 2635
rect 69808 2604 70317 2632
rect 69808 2592 69814 2604
rect 70305 2601 70317 2604
rect 70351 2601 70363 2635
rect 70305 2595 70363 2601
rect 71130 2592 71136 2644
rect 71188 2632 71194 2644
rect 71593 2635 71651 2641
rect 71593 2632 71605 2635
rect 71188 2604 71605 2632
rect 71188 2592 71194 2604
rect 71593 2601 71605 2604
rect 71639 2601 71651 2635
rect 71593 2595 71651 2601
rect 72234 2592 72240 2644
rect 72292 2592 72298 2644
rect 72421 2635 72479 2641
rect 72421 2601 72433 2635
rect 72467 2601 72479 2635
rect 73525 2635 73583 2641
rect 73525 2632 73537 2635
rect 72421 2595 72479 2601
rect 72620 2604 73537 2632
rect 49694 2564 49700 2576
rect 48700 2536 49700 2564
rect 45094 2456 45100 2508
rect 45152 2496 45158 2508
rect 46845 2499 46903 2505
rect 46845 2496 46857 2499
rect 45152 2468 46857 2496
rect 45152 2456 45158 2468
rect 43441 2431 43499 2437
rect 43441 2397 43453 2431
rect 43487 2428 43499 2431
rect 43809 2431 43867 2437
rect 43809 2428 43821 2431
rect 43487 2400 43821 2428
rect 43487 2397 43499 2400
rect 43441 2391 43499 2397
rect 43809 2397 43821 2400
rect 43855 2397 43867 2431
rect 43809 2391 43867 2397
rect 44821 2431 44879 2437
rect 44821 2397 44833 2431
rect 44867 2397 44879 2431
rect 44821 2391 44879 2397
rect 45002 2388 45008 2440
rect 45060 2388 45066 2440
rect 45186 2388 45192 2440
rect 45244 2428 45250 2440
rect 45373 2431 45431 2437
rect 45373 2428 45385 2431
rect 45244 2400 45385 2428
rect 45244 2388 45250 2400
rect 45373 2397 45385 2400
rect 45419 2428 45431 2431
rect 45649 2431 45707 2437
rect 45649 2428 45661 2431
rect 45419 2400 45661 2428
rect 45419 2397 45431 2400
rect 45373 2391 45431 2397
rect 45649 2397 45661 2400
rect 45695 2397 45707 2431
rect 45649 2391 45707 2397
rect 45830 2388 45836 2440
rect 45888 2388 45894 2440
rect 46216 2437 46244 2468
rect 46845 2465 46857 2468
rect 46891 2465 46903 2499
rect 46845 2459 46903 2465
rect 46201 2431 46259 2437
rect 46201 2397 46213 2431
rect 46247 2397 46259 2431
rect 46201 2391 46259 2397
rect 46474 2388 46480 2440
rect 46532 2388 46538 2440
rect 47118 2388 47124 2440
rect 47176 2388 47182 2440
rect 47762 2388 47768 2440
rect 47820 2388 47826 2440
rect 48700 2437 48728 2536
rect 49694 2524 49700 2536
rect 49752 2524 49758 2576
rect 50801 2567 50859 2573
rect 50801 2533 50813 2567
rect 50847 2533 50859 2567
rect 50801 2527 50859 2533
rect 53101 2567 53159 2573
rect 53101 2533 53113 2567
rect 53147 2564 53159 2567
rect 54294 2564 54300 2576
rect 53147 2536 54300 2564
rect 53147 2533 53159 2536
rect 53101 2527 53159 2533
rect 49712 2496 49740 2524
rect 50816 2496 50844 2527
rect 54294 2524 54300 2536
rect 54352 2524 54358 2576
rect 54389 2567 54447 2573
rect 54389 2533 54401 2567
rect 54435 2564 54447 2567
rect 55401 2567 55459 2573
rect 54435 2536 54708 2564
rect 54435 2533 54447 2536
rect 54389 2527 54447 2533
rect 49712 2468 50384 2496
rect 50816 2468 54064 2496
rect 48685 2431 48743 2437
rect 48685 2397 48697 2431
rect 48731 2397 48743 2431
rect 48685 2391 48743 2397
rect 49050 2388 49056 2440
rect 49108 2388 49114 2440
rect 49697 2431 49755 2437
rect 49697 2397 49709 2431
rect 49743 2428 49755 2431
rect 49786 2428 49792 2440
rect 49743 2400 49792 2428
rect 49743 2397 49755 2400
rect 49697 2391 49755 2397
rect 49786 2388 49792 2400
rect 49844 2388 49850 2440
rect 50356 2437 50384 2468
rect 50341 2431 50399 2437
rect 50341 2397 50353 2431
rect 50387 2397 50399 2431
rect 50341 2391 50399 2397
rect 50617 2431 50675 2437
rect 50617 2397 50629 2431
rect 50663 2397 50675 2431
rect 50617 2391 50675 2397
rect 40773 2363 40831 2369
rect 40773 2360 40785 2363
rect 38887 2332 40785 2360
rect 38887 2329 38899 2332
rect 38841 2323 38899 2329
rect 40773 2329 40785 2332
rect 40819 2360 40831 2363
rect 43364 2360 43392 2388
rect 49513 2363 49571 2369
rect 40819 2332 43392 2360
rect 43824 2332 45232 2360
rect 40819 2329 40831 2332
rect 40773 2323 40831 2329
rect 43824 2304 43852 2332
rect 32858 2252 32864 2304
rect 32916 2292 32922 2304
rect 33137 2295 33195 2301
rect 33137 2292 33149 2295
rect 32916 2264 33149 2292
rect 32916 2252 32922 2264
rect 33137 2261 33149 2264
rect 33183 2261 33195 2295
rect 33137 2255 33195 2261
rect 42518 2252 42524 2304
rect 42576 2292 42582 2304
rect 42705 2295 42763 2301
rect 42705 2292 42717 2295
rect 42576 2264 42717 2292
rect 42576 2252 42582 2264
rect 42705 2261 42717 2264
rect 42751 2261 42763 2295
rect 42705 2255 42763 2261
rect 43806 2252 43812 2304
rect 43864 2252 43870 2304
rect 45204 2301 45232 2332
rect 49513 2329 49525 2363
rect 49559 2360 49571 2363
rect 50154 2360 50160 2372
rect 49559 2332 50160 2360
rect 49559 2329 49571 2332
rect 49513 2323 49571 2329
rect 50154 2320 50160 2332
rect 50212 2320 50218 2372
rect 50246 2320 50252 2372
rect 50304 2360 50310 2372
rect 50632 2360 50660 2391
rect 51258 2388 51264 2440
rect 51316 2388 51322 2440
rect 51626 2388 51632 2440
rect 51684 2388 51690 2440
rect 52273 2431 52331 2437
rect 52273 2428 52285 2431
rect 52196 2400 52285 2428
rect 51353 2363 51411 2369
rect 51353 2360 51365 2363
rect 50304 2332 51365 2360
rect 50304 2320 50310 2332
rect 51353 2329 51365 2332
rect 51399 2329 51411 2363
rect 51353 2323 51411 2329
rect 52196 2304 52224 2400
rect 52273 2397 52285 2400
rect 52319 2397 52331 2431
rect 52917 2431 52975 2437
rect 52917 2428 52929 2431
rect 52273 2391 52331 2397
rect 52840 2400 52929 2428
rect 52840 2304 52868 2400
rect 52917 2397 52929 2400
rect 52963 2397 52975 2431
rect 52917 2391 52975 2397
rect 53558 2388 53564 2440
rect 53616 2388 53622 2440
rect 53929 2431 53987 2437
rect 53929 2397 53941 2431
rect 53975 2397 53987 2431
rect 53929 2391 53987 2397
rect 53377 2363 53435 2369
rect 53377 2329 53389 2363
rect 53423 2360 53435 2363
rect 53944 2360 53972 2391
rect 53423 2332 53972 2360
rect 54036 2360 54064 2468
rect 54478 2456 54484 2508
rect 54536 2496 54542 2508
rect 54680 2505 54708 2536
rect 55401 2533 55413 2567
rect 55447 2564 55459 2567
rect 55490 2564 55496 2576
rect 55447 2536 55496 2564
rect 55447 2533 55459 2536
rect 55401 2527 55459 2533
rect 55490 2524 55496 2536
rect 55548 2524 55554 2576
rect 57330 2524 57336 2576
rect 57388 2564 57394 2576
rect 58069 2567 58127 2573
rect 58069 2564 58081 2567
rect 57388 2536 58081 2564
rect 57388 2524 57394 2536
rect 58069 2533 58081 2536
rect 58115 2533 58127 2567
rect 58069 2527 58127 2533
rect 59722 2524 59728 2576
rect 59780 2564 59786 2576
rect 60645 2567 60703 2573
rect 60645 2564 60657 2567
rect 59780 2536 60657 2564
rect 59780 2524 59786 2536
rect 60645 2533 60657 2536
rect 60691 2533 60703 2567
rect 60645 2527 60703 2533
rect 61289 2567 61347 2573
rect 61289 2533 61301 2567
rect 61335 2533 61347 2567
rect 61289 2527 61347 2533
rect 67269 2567 67327 2573
rect 67269 2533 67281 2567
rect 67315 2533 67327 2567
rect 67269 2527 67327 2533
rect 67913 2567 67971 2573
rect 67913 2533 67925 2567
rect 67959 2564 67971 2567
rect 69014 2564 69020 2576
rect 67959 2536 69020 2564
rect 67959 2533 67971 2536
rect 67913 2527 67971 2533
rect 54665 2499 54723 2505
rect 54536 2468 54616 2496
rect 54536 2456 54542 2468
rect 54110 2388 54116 2440
rect 54168 2428 54174 2440
rect 54588 2437 54616 2468
rect 54665 2465 54677 2499
rect 54711 2465 54723 2499
rect 54665 2459 54723 2465
rect 55677 2499 55735 2505
rect 55677 2465 55689 2499
rect 55723 2496 55735 2499
rect 56042 2496 56048 2508
rect 55723 2468 56048 2496
rect 55723 2465 55735 2468
rect 55677 2459 55735 2465
rect 56042 2456 56048 2468
rect 56100 2456 56106 2508
rect 56686 2456 56692 2508
rect 56744 2496 56750 2508
rect 57422 2496 57428 2508
rect 56744 2468 57428 2496
rect 56744 2456 56750 2468
rect 57422 2456 57428 2468
rect 57480 2496 57486 2508
rect 58158 2496 58164 2508
rect 57480 2468 57560 2496
rect 57480 2456 57486 2468
rect 54205 2431 54263 2437
rect 54205 2428 54217 2431
rect 54168 2400 54217 2428
rect 54168 2388 54174 2400
rect 54205 2397 54217 2400
rect 54251 2397 54263 2431
rect 54205 2391 54263 2397
rect 54573 2431 54631 2437
rect 54573 2397 54585 2431
rect 54619 2397 54631 2431
rect 54573 2391 54631 2397
rect 54846 2388 54852 2440
rect 54904 2388 54910 2440
rect 55306 2428 55312 2440
rect 55186 2400 55312 2428
rect 55186 2360 55214 2400
rect 55306 2388 55312 2400
rect 55364 2388 55370 2440
rect 57532 2437 57560 2468
rect 57900 2468 58164 2496
rect 57900 2437 57928 2468
rect 58158 2456 58164 2468
rect 58216 2456 58222 2508
rect 59630 2456 59636 2508
rect 59688 2496 59694 2508
rect 61304 2496 61332 2527
rect 59688 2468 61332 2496
rect 67284 2496 67312 2527
rect 69014 2524 69020 2536
rect 69072 2524 69078 2576
rect 69201 2567 69259 2573
rect 69201 2533 69213 2567
rect 69247 2564 69259 2567
rect 71222 2564 71228 2576
rect 69247 2536 71228 2564
rect 69247 2533 69259 2536
rect 69201 2527 69259 2533
rect 71222 2524 71228 2536
rect 71280 2524 71286 2576
rect 72436 2496 72464 2595
rect 72620 2505 72648 2604
rect 73525 2601 73537 2604
rect 73571 2601 73583 2635
rect 73525 2595 73583 2601
rect 74074 2592 74080 2644
rect 74132 2632 74138 2644
rect 74169 2635 74227 2641
rect 74169 2632 74181 2635
rect 74132 2604 74181 2632
rect 74132 2592 74138 2604
rect 74169 2601 74181 2604
rect 74215 2601 74227 2635
rect 74169 2595 74227 2601
rect 74258 2592 74264 2644
rect 74316 2632 74322 2644
rect 75457 2635 75515 2641
rect 75457 2632 75469 2635
rect 74316 2604 75469 2632
rect 74316 2592 74322 2604
rect 75457 2601 75469 2604
rect 75503 2601 75515 2635
rect 75457 2595 75515 2601
rect 76098 2592 76104 2644
rect 76156 2592 76162 2644
rect 77386 2592 77392 2644
rect 77444 2592 77450 2644
rect 77754 2592 77760 2644
rect 77812 2592 77818 2644
rect 74813 2567 74871 2573
rect 74813 2564 74825 2567
rect 72712 2536 74825 2564
rect 67284 2468 72464 2496
rect 72605 2499 72663 2505
rect 59688 2456 59694 2468
rect 72605 2465 72617 2499
rect 72651 2465 72663 2499
rect 72605 2459 72663 2465
rect 57517 2431 57575 2437
rect 57517 2397 57529 2431
rect 57563 2397 57575 2431
rect 57517 2391 57575 2397
rect 57885 2431 57943 2437
rect 57885 2397 57897 2431
rect 57931 2397 57943 2431
rect 57885 2391 57943 2397
rect 54036 2332 55214 2360
rect 55953 2363 56011 2369
rect 53423 2329 53435 2332
rect 53377 2323 53435 2329
rect 45189 2295 45247 2301
rect 45189 2261 45201 2295
rect 45235 2261 45247 2295
rect 45189 2255 45247 2261
rect 45554 2252 45560 2304
rect 45612 2252 45618 2304
rect 45738 2252 45744 2304
rect 45796 2292 45802 2304
rect 46017 2295 46075 2301
rect 46017 2292 46029 2295
rect 45796 2264 46029 2292
rect 45796 2252 45802 2264
rect 46017 2261 46029 2264
rect 46063 2261 46075 2295
rect 46017 2255 46075 2261
rect 46382 2252 46388 2304
rect 46440 2252 46446 2304
rect 46474 2252 46480 2304
rect 46532 2292 46538 2304
rect 46661 2295 46719 2301
rect 46661 2292 46673 2295
rect 46532 2264 46673 2292
rect 46532 2252 46538 2264
rect 46661 2261 46673 2264
rect 46707 2261 46719 2295
rect 46661 2255 46719 2261
rect 47026 2252 47032 2304
rect 47084 2292 47090 2304
rect 47305 2295 47363 2301
rect 47305 2292 47317 2295
rect 47084 2264 47317 2292
rect 47084 2252 47090 2264
rect 47305 2261 47317 2264
rect 47351 2261 47363 2295
rect 47305 2255 47363 2261
rect 47670 2252 47676 2304
rect 47728 2292 47734 2304
rect 47949 2295 48007 2301
rect 47949 2292 47961 2295
rect 47728 2264 47961 2292
rect 47728 2252 47734 2264
rect 47949 2261 47961 2264
rect 47995 2261 48007 2295
rect 47949 2255 48007 2261
rect 48314 2252 48320 2304
rect 48372 2292 48378 2304
rect 48501 2295 48559 2301
rect 48501 2292 48513 2295
rect 48372 2264 48513 2292
rect 48372 2252 48378 2264
rect 48501 2261 48513 2264
rect 48547 2261 48559 2295
rect 48501 2255 48559 2261
rect 48958 2252 48964 2304
rect 49016 2292 49022 2304
rect 49237 2295 49295 2301
rect 49237 2292 49249 2295
rect 49016 2264 49249 2292
rect 49016 2252 49022 2264
rect 49237 2261 49249 2264
rect 49283 2261 49295 2295
rect 49237 2255 49295 2261
rect 49602 2252 49608 2304
rect 49660 2292 49666 2304
rect 49881 2295 49939 2301
rect 49881 2292 49893 2295
rect 49660 2264 49893 2292
rect 49660 2252 49666 2264
rect 49881 2261 49893 2264
rect 49927 2261 49939 2295
rect 49881 2255 49939 2261
rect 50890 2252 50896 2304
rect 50948 2292 50954 2304
rect 51077 2295 51135 2301
rect 51077 2292 51089 2295
rect 50948 2264 51089 2292
rect 50948 2252 50954 2264
rect 51077 2261 51089 2264
rect 51123 2261 51135 2295
rect 51077 2255 51135 2261
rect 51534 2252 51540 2304
rect 51592 2292 51598 2304
rect 51813 2295 51871 2301
rect 51813 2292 51825 2295
rect 51592 2264 51825 2292
rect 51592 2252 51598 2264
rect 51813 2261 51825 2264
rect 51859 2261 51871 2295
rect 51813 2255 51871 2261
rect 52178 2252 52184 2304
rect 52236 2252 52242 2304
rect 52454 2252 52460 2304
rect 52512 2252 52518 2304
rect 52822 2252 52828 2304
rect 52880 2252 52886 2304
rect 53466 2252 53472 2304
rect 53524 2292 53530 2304
rect 53745 2295 53803 2301
rect 53745 2292 53757 2295
rect 53524 2264 53757 2292
rect 53524 2252 53530 2264
rect 53745 2261 53757 2264
rect 53791 2261 53803 2295
rect 53944 2292 53972 2332
rect 55953 2329 55965 2363
rect 55999 2329 56011 2363
rect 55953 2323 56011 2329
rect 54754 2292 54760 2304
rect 53944 2264 54760 2292
rect 53745 2255 53803 2261
rect 54754 2252 54760 2264
rect 54812 2252 54818 2304
rect 55030 2252 55036 2304
rect 55088 2252 55094 2304
rect 55968 2292 55996 2323
rect 56594 2320 56600 2372
rect 56652 2320 56658 2372
rect 57900 2360 57928 2391
rect 57974 2388 57980 2440
rect 58032 2428 58038 2440
rect 58253 2431 58311 2437
rect 58253 2428 58265 2431
rect 58032 2400 58265 2428
rect 58032 2388 58038 2400
rect 58253 2397 58265 2400
rect 58299 2428 58311 2431
rect 58529 2431 58587 2437
rect 58529 2428 58541 2431
rect 58299 2400 58541 2428
rect 58299 2397 58311 2400
rect 58253 2391 58311 2397
rect 58529 2397 58541 2400
rect 58575 2397 58587 2431
rect 58529 2391 58587 2397
rect 58897 2431 58955 2437
rect 58897 2397 58909 2431
rect 58943 2428 58955 2431
rect 59541 2431 59599 2437
rect 59541 2428 59553 2431
rect 58943 2400 58977 2428
rect 59280 2400 59553 2428
rect 58943 2397 58955 2400
rect 58897 2391 58955 2397
rect 57440 2332 57928 2360
rect 56962 2292 56968 2304
rect 55968 2264 56968 2292
rect 56962 2252 56968 2264
rect 57020 2252 57026 2304
rect 57440 2301 57468 2332
rect 58618 2320 58624 2372
rect 58676 2360 58682 2372
rect 58912 2360 58940 2391
rect 58989 2363 59047 2369
rect 58989 2360 59001 2363
rect 58676 2332 59001 2360
rect 58676 2320 58682 2332
rect 58989 2329 59001 2332
rect 59035 2329 59047 2363
rect 58989 2323 59047 2329
rect 59280 2304 59308 2400
rect 59541 2397 59553 2400
rect 59587 2397 59599 2431
rect 60185 2431 60243 2437
rect 60185 2428 60197 2431
rect 59541 2391 59599 2397
rect 59924 2400 60197 2428
rect 59924 2304 59952 2400
rect 60185 2397 60197 2400
rect 60231 2397 60243 2431
rect 60829 2431 60887 2437
rect 60829 2428 60841 2431
rect 60185 2391 60243 2397
rect 60568 2400 60841 2428
rect 60568 2304 60596 2400
rect 60829 2397 60841 2400
rect 60875 2397 60887 2431
rect 61473 2431 61531 2437
rect 61473 2428 61485 2431
rect 60829 2391 60887 2397
rect 61212 2400 61485 2428
rect 61212 2304 61240 2400
rect 61473 2397 61485 2400
rect 61519 2397 61531 2431
rect 61473 2391 61531 2397
rect 61746 2388 61752 2440
rect 61804 2428 61810 2440
rect 61933 2431 61991 2437
rect 61933 2428 61945 2431
rect 61804 2400 61945 2428
rect 61804 2388 61810 2400
rect 61933 2397 61945 2400
rect 61979 2397 61991 2431
rect 61933 2391 61991 2397
rect 62390 2388 62396 2440
rect 62448 2428 62454 2440
rect 62577 2431 62635 2437
rect 62577 2428 62589 2431
rect 62448 2400 62589 2428
rect 62448 2388 62454 2400
rect 62577 2397 62589 2400
rect 62623 2397 62635 2431
rect 62577 2391 62635 2397
rect 63218 2388 63224 2440
rect 63276 2388 63282 2440
rect 63678 2388 63684 2440
rect 63736 2428 63742 2440
rect 63865 2431 63923 2437
rect 63865 2428 63877 2431
rect 63736 2400 63877 2428
rect 63736 2388 63742 2400
rect 63865 2397 63877 2400
rect 63911 2397 63923 2431
rect 63865 2391 63923 2397
rect 64322 2388 64328 2440
rect 64380 2428 64386 2440
rect 64509 2431 64567 2437
rect 64509 2428 64521 2431
rect 64380 2400 64521 2428
rect 64380 2388 64386 2400
rect 64509 2397 64521 2400
rect 64555 2397 64567 2431
rect 65153 2431 65211 2437
rect 65153 2428 65165 2431
rect 64509 2391 64567 2397
rect 65076 2400 65165 2428
rect 65076 2304 65104 2400
rect 65153 2397 65165 2400
rect 65199 2397 65211 2431
rect 65797 2431 65855 2437
rect 65797 2428 65809 2431
rect 65153 2391 65211 2397
rect 65720 2400 65809 2428
rect 65720 2304 65748 2400
rect 65797 2397 65809 2400
rect 65843 2397 65855 2431
rect 66441 2431 66499 2437
rect 66441 2428 66453 2431
rect 65797 2391 65855 2397
rect 66272 2400 66453 2428
rect 66272 2304 66300 2400
rect 66441 2397 66453 2400
rect 66487 2397 66499 2431
rect 67085 2431 67143 2437
rect 67085 2428 67097 2431
rect 66441 2391 66499 2397
rect 67008 2400 67097 2428
rect 67008 2304 67036 2400
rect 67085 2397 67097 2400
rect 67131 2397 67143 2431
rect 67729 2431 67787 2437
rect 67729 2428 67741 2431
rect 67085 2391 67143 2397
rect 67652 2400 67741 2428
rect 67652 2304 67680 2400
rect 67729 2397 67741 2400
rect 67775 2397 67787 2431
rect 67729 2391 67787 2397
rect 68646 2388 68652 2440
rect 68704 2388 68710 2440
rect 69017 2431 69075 2437
rect 69017 2428 69029 2431
rect 68940 2400 69029 2428
rect 68940 2304 68968 2400
rect 69017 2397 69029 2400
rect 69063 2397 69075 2431
rect 69845 2431 69903 2437
rect 69845 2428 69857 2431
rect 69017 2391 69075 2397
rect 69584 2400 69857 2428
rect 69584 2304 69612 2400
rect 69845 2397 69857 2400
rect 69891 2397 69903 2431
rect 70489 2431 70547 2437
rect 70489 2428 70501 2431
rect 69845 2391 69903 2397
rect 70228 2400 70501 2428
rect 70228 2304 70256 2400
rect 70489 2397 70501 2400
rect 70535 2397 70547 2431
rect 70949 2431 71007 2437
rect 70949 2428 70961 2431
rect 70489 2391 70547 2397
rect 70872 2400 70961 2428
rect 70872 2304 70900 2400
rect 70949 2397 70961 2400
rect 70995 2397 71007 2431
rect 71777 2431 71835 2437
rect 71777 2428 71789 2431
rect 70949 2391 71007 2397
rect 71516 2400 71789 2428
rect 71516 2304 71544 2400
rect 71777 2397 71789 2400
rect 71823 2397 71835 2431
rect 71777 2391 71835 2397
rect 71961 2431 72019 2437
rect 71961 2397 71973 2431
rect 72007 2428 72019 2431
rect 72050 2428 72056 2440
rect 72007 2400 72056 2428
rect 72007 2397 72019 2400
rect 71961 2391 72019 2397
rect 72050 2388 72056 2400
rect 72108 2388 72114 2440
rect 72712 2437 72740 2536
rect 74813 2533 74825 2536
rect 74859 2533 74871 2567
rect 74813 2527 74871 2533
rect 72421 2431 72479 2437
rect 72421 2428 72433 2431
rect 72160 2400 72433 2428
rect 57425 2295 57483 2301
rect 57425 2261 57437 2295
rect 57471 2261 57483 2295
rect 57425 2255 57483 2261
rect 57698 2252 57704 2304
rect 57756 2252 57762 2304
rect 58342 2252 58348 2304
rect 58400 2292 58406 2304
rect 58713 2295 58771 2301
rect 58713 2292 58725 2295
rect 58400 2264 58725 2292
rect 58400 2252 58406 2264
rect 58713 2261 58725 2264
rect 58759 2261 58771 2295
rect 58713 2255 58771 2261
rect 59262 2252 59268 2304
rect 59320 2252 59326 2304
rect 59354 2252 59360 2304
rect 59412 2252 59418 2304
rect 59906 2252 59912 2304
rect 59964 2252 59970 2304
rect 60550 2252 60556 2304
rect 60608 2252 60614 2304
rect 61194 2252 61200 2304
rect 61252 2252 61258 2304
rect 61838 2252 61844 2304
rect 61896 2292 61902 2304
rect 62117 2295 62175 2301
rect 62117 2292 62129 2295
rect 61896 2264 62129 2292
rect 61896 2252 61902 2264
rect 62117 2261 62129 2264
rect 62163 2261 62175 2295
rect 62117 2255 62175 2261
rect 62482 2252 62488 2304
rect 62540 2292 62546 2304
rect 62761 2295 62819 2301
rect 62761 2292 62773 2295
rect 62540 2264 62773 2292
rect 62540 2252 62546 2264
rect 62761 2261 62773 2264
rect 62807 2261 62819 2295
rect 62761 2255 62819 2261
rect 63126 2252 63132 2304
rect 63184 2292 63190 2304
rect 63405 2295 63463 2301
rect 63405 2292 63417 2295
rect 63184 2264 63417 2292
rect 63184 2252 63190 2264
rect 63405 2261 63417 2264
rect 63451 2261 63463 2295
rect 63405 2255 63463 2261
rect 63770 2252 63776 2304
rect 63828 2292 63834 2304
rect 64049 2295 64107 2301
rect 64049 2292 64061 2295
rect 63828 2264 64061 2292
rect 63828 2252 63834 2264
rect 64049 2261 64061 2264
rect 64095 2261 64107 2295
rect 64049 2255 64107 2261
rect 64414 2252 64420 2304
rect 64472 2292 64478 2304
rect 64693 2295 64751 2301
rect 64693 2292 64705 2295
rect 64472 2264 64705 2292
rect 64472 2252 64478 2264
rect 64693 2261 64705 2264
rect 64739 2261 64751 2295
rect 64693 2255 64751 2261
rect 65058 2252 65064 2304
rect 65116 2252 65122 2304
rect 65334 2252 65340 2304
rect 65392 2252 65398 2304
rect 65702 2252 65708 2304
rect 65760 2252 65766 2304
rect 65981 2295 66039 2301
rect 65981 2261 65993 2295
rect 66027 2292 66039 2295
rect 66070 2292 66076 2304
rect 66027 2264 66076 2292
rect 66027 2261 66039 2264
rect 65981 2255 66039 2261
rect 66070 2252 66076 2264
rect 66128 2252 66134 2304
rect 66254 2252 66260 2304
rect 66312 2252 66318 2304
rect 66990 2252 66996 2304
rect 67048 2252 67054 2304
rect 67634 2252 67640 2304
rect 67692 2252 67698 2304
rect 68278 2252 68284 2304
rect 68336 2292 68342 2304
rect 68465 2295 68523 2301
rect 68465 2292 68477 2295
rect 68336 2264 68477 2292
rect 68336 2252 68342 2264
rect 68465 2261 68477 2264
rect 68511 2261 68523 2295
rect 68465 2255 68523 2261
rect 68922 2252 68928 2304
rect 68980 2252 68986 2304
rect 69566 2252 69572 2304
rect 69624 2252 69630 2304
rect 70210 2252 70216 2304
rect 70268 2252 70274 2304
rect 70854 2252 70860 2304
rect 70912 2252 70918 2304
rect 71130 2252 71136 2304
rect 71188 2252 71194 2304
rect 71498 2252 71504 2304
rect 71556 2252 71562 2304
rect 72160 2301 72188 2400
rect 72421 2397 72433 2400
rect 72467 2397 72479 2431
rect 72421 2391 72479 2397
rect 72697 2431 72755 2437
rect 72697 2397 72709 2431
rect 72743 2397 72755 2431
rect 72697 2391 72755 2397
rect 72878 2388 72884 2440
rect 72936 2388 72942 2440
rect 73709 2431 73767 2437
rect 73709 2397 73721 2431
rect 73755 2428 73767 2431
rect 74353 2431 74411 2437
rect 74353 2428 74365 2431
rect 73755 2400 73789 2428
rect 74092 2400 74365 2428
rect 73755 2397 73767 2400
rect 73709 2391 73767 2397
rect 72234 2320 72240 2372
rect 72292 2360 72298 2372
rect 73341 2363 73399 2369
rect 73341 2360 73353 2363
rect 72292 2332 73353 2360
rect 72292 2320 72298 2332
rect 73341 2329 73353 2332
rect 73387 2329 73399 2363
rect 73341 2323 73399 2329
rect 73430 2320 73436 2372
rect 73488 2360 73494 2372
rect 73724 2360 73752 2391
rect 73801 2363 73859 2369
rect 73801 2360 73813 2363
rect 73488 2332 73813 2360
rect 73488 2320 73494 2332
rect 73801 2329 73813 2332
rect 73847 2329 73859 2363
rect 73801 2323 73859 2329
rect 74092 2304 74120 2400
rect 74353 2397 74365 2400
rect 74399 2397 74411 2431
rect 74997 2431 75055 2437
rect 74997 2428 75009 2431
rect 74353 2391 74411 2397
rect 74736 2400 75009 2428
rect 74736 2304 74764 2400
rect 74997 2397 75009 2400
rect 75043 2397 75055 2431
rect 75641 2431 75699 2437
rect 75641 2428 75653 2431
rect 74997 2391 75055 2397
rect 75380 2400 75653 2428
rect 75380 2304 75408 2400
rect 75641 2397 75653 2400
rect 75687 2397 75699 2431
rect 76285 2431 76343 2437
rect 76285 2428 76297 2431
rect 75641 2391 75699 2397
rect 76024 2400 76297 2428
rect 76024 2304 76052 2400
rect 76285 2397 76297 2400
rect 76331 2397 76343 2431
rect 76285 2391 76343 2397
rect 76742 2388 76748 2440
rect 76800 2388 76806 2440
rect 77573 2431 77631 2437
rect 77573 2428 77585 2431
rect 77312 2400 77585 2428
rect 77312 2304 77340 2400
rect 77573 2397 77585 2400
rect 77619 2397 77631 2431
rect 77573 2391 77631 2397
rect 77938 2388 77944 2440
rect 77996 2388 78002 2440
rect 78030 2388 78036 2440
rect 78088 2388 78094 2440
rect 72145 2295 72203 2301
rect 72145 2261 72157 2295
rect 72191 2261 72203 2295
rect 72145 2255 72203 2261
rect 72786 2252 72792 2304
rect 72844 2292 72850 2304
rect 73065 2295 73123 2301
rect 73065 2292 73077 2295
rect 72844 2264 73077 2292
rect 72844 2252 72850 2264
rect 73065 2261 73077 2264
rect 73111 2261 73123 2295
rect 73065 2255 73123 2261
rect 74074 2252 74080 2304
rect 74132 2252 74138 2304
rect 74718 2252 74724 2304
rect 74776 2252 74782 2304
rect 75362 2252 75368 2304
rect 75420 2252 75426 2304
rect 76006 2252 76012 2304
rect 76064 2252 76070 2304
rect 76650 2252 76656 2304
rect 76708 2292 76714 2304
rect 76929 2295 76987 2301
rect 76929 2292 76941 2295
rect 76708 2264 76941 2292
rect 76708 2252 76714 2264
rect 76929 2261 76941 2264
rect 76975 2261 76987 2295
rect 76929 2255 76987 2261
rect 77294 2252 77300 2304
rect 77352 2252 77358 2304
rect 78217 2295 78275 2301
rect 78217 2261 78229 2295
rect 78263 2292 78275 2295
rect 78582 2292 78588 2304
rect 78263 2264 78588 2292
rect 78263 2261 78275 2264
rect 78217 2255 78275 2261
rect 78582 2252 78588 2264
rect 78640 2252 78646 2304
rect 1104 2202 78844 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 66314 2202
rect 66366 2150 66378 2202
rect 66430 2150 66442 2202
rect 66494 2150 66506 2202
rect 66558 2150 66570 2202
rect 66622 2150 78844 2202
rect 1104 2128 78844 2150
rect 44450 2048 44456 2100
rect 44508 2088 44514 2100
rect 45186 2088 45192 2100
rect 44508 2060 45192 2088
rect 44508 2048 44514 2060
rect 45186 2048 45192 2060
rect 45244 2048 45250 2100
rect 45554 2048 45560 2100
rect 45612 2088 45618 2100
rect 54846 2088 54852 2100
rect 45612 2060 54852 2088
rect 45612 2048 45618 2060
rect 54846 2048 54852 2060
rect 54904 2048 54910 2100
rect 55030 2048 55036 2100
rect 55088 2088 55094 2100
rect 59998 2088 60004 2100
rect 55088 2060 60004 2088
rect 55088 2048 55094 2060
rect 59998 2048 60004 2060
rect 60056 2048 60062 2100
rect 65334 2048 65340 2100
rect 65392 2088 65398 2100
rect 65392 2060 66116 2088
rect 65392 2048 65398 2060
rect 43346 1980 43352 2032
rect 43404 2020 43410 2032
rect 43404 1992 45554 2020
rect 43404 1980 43410 1992
rect 45526 1952 45554 1992
rect 46382 1980 46388 2032
rect 46440 2020 46446 2032
rect 65978 2020 65984 2032
rect 46440 1992 65984 2020
rect 46440 1980 46446 1992
rect 65978 1980 65984 1992
rect 66036 1980 66042 2032
rect 66088 2020 66116 2060
rect 72418 2020 72424 2032
rect 66088 1992 72424 2020
rect 72418 1980 72424 1992
rect 72476 1980 72482 2032
rect 50154 1952 50160 1964
rect 45526 1924 50160 1952
rect 50154 1912 50160 1924
rect 50212 1912 50218 1964
rect 54478 1912 54484 1964
rect 54536 1952 54542 1964
rect 59354 1952 59360 1964
rect 54536 1924 59360 1952
rect 54536 1912 54542 1924
rect 59354 1912 59360 1924
rect 59412 1912 59418 1964
rect 66070 1912 66076 1964
rect 66128 1952 66134 1964
rect 72510 1952 72516 1964
rect 66128 1924 72516 1952
rect 66128 1912 66134 1924
rect 72510 1912 72516 1924
rect 72568 1912 72574 1964
rect 52454 1844 52460 1896
rect 52512 1884 52518 1896
rect 58802 1884 58808 1896
rect 52512 1856 58808 1884
rect 52512 1844 52518 1856
rect 58802 1844 58808 1856
rect 58860 1844 58866 1896
rect 50154 1776 50160 1828
rect 50212 1816 50218 1828
rect 55214 1816 55220 1828
rect 50212 1788 55220 1816
rect 50212 1776 50218 1788
rect 55214 1776 55220 1788
rect 55272 1776 55278 1828
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 38660 37408 38712 37460
rect 45100 37408 45152 37460
rect 46388 37408 46440 37460
rect 43812 37340 43864 37392
rect 36268 37247 36320 37256
rect 36268 37213 36277 37247
rect 36277 37213 36311 37247
rect 36311 37213 36320 37247
rect 36268 37204 36320 37213
rect 40500 37247 40552 37256
rect 40500 37213 40509 37247
rect 40509 37213 40543 37247
rect 40543 37213 40552 37247
rect 40500 37204 40552 37213
rect 40868 37204 40920 37256
rect 39396 37136 39448 37188
rect 43904 37136 43956 37188
rect 44364 37136 44416 37188
rect 46112 37136 46164 37188
rect 35440 37068 35492 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 66314 36966 66366 37018
rect 66378 36966 66430 37018
rect 66442 36966 66494 37018
rect 66506 36966 66558 37018
rect 66570 36966 66622 37018
rect 36268 36864 36320 36916
rect 39948 36864 40000 36916
rect 40592 36864 40644 36916
rect 41236 36864 41288 36916
rect 41880 36864 41932 36916
rect 42524 36864 42576 36916
rect 43168 36864 43220 36916
rect 44456 36864 44508 36916
rect 45744 36864 45796 36916
rect 46112 36907 46164 36916
rect 46112 36873 46121 36907
rect 46121 36873 46155 36907
rect 46155 36873 46164 36907
rect 46112 36864 46164 36873
rect 47032 36864 47084 36916
rect 47676 36907 47728 36916
rect 47676 36873 47685 36907
rect 47685 36873 47719 36907
rect 47719 36873 47728 36907
rect 47676 36864 47728 36873
rect 48320 36864 48372 36916
rect 48964 36907 49016 36916
rect 48964 36873 48973 36907
rect 48973 36873 49007 36907
rect 49007 36873 49016 36907
rect 48964 36864 49016 36873
rect 49608 36864 49660 36916
rect 50252 36864 50304 36916
rect 50896 36864 50948 36916
rect 51540 36864 51592 36916
rect 52184 36864 52236 36916
rect 52828 36907 52880 36916
rect 52828 36873 52837 36907
rect 52837 36873 52871 36907
rect 52871 36873 52880 36907
rect 52828 36864 52880 36873
rect 53472 36907 53524 36916
rect 53472 36873 53481 36907
rect 53481 36873 53515 36907
rect 53515 36873 53524 36907
rect 53472 36864 53524 36873
rect 54116 36864 54168 36916
rect 54760 36864 54812 36916
rect 55404 36864 55456 36916
rect 56048 36864 56100 36916
rect 56692 36864 56744 36916
rect 57336 36864 57388 36916
rect 57980 36907 58032 36916
rect 57980 36873 57989 36907
rect 57989 36873 58023 36907
rect 58023 36873 58032 36907
rect 57980 36864 58032 36873
rect 58624 36864 58676 36916
rect 59268 36864 59320 36916
rect 59912 36907 59964 36916
rect 59912 36873 59921 36907
rect 59921 36873 59955 36907
rect 59955 36873 59964 36907
rect 59912 36864 59964 36873
rect 60556 36864 60608 36916
rect 61200 36907 61252 36916
rect 61200 36873 61209 36907
rect 61209 36873 61243 36907
rect 61243 36873 61252 36907
rect 61200 36864 61252 36873
rect 61844 36864 61896 36916
rect 62488 36864 62540 36916
rect 63132 36864 63184 36916
rect 63776 36864 63828 36916
rect 64420 36864 64472 36916
rect 65064 36864 65116 36916
rect 65524 36864 65576 36916
rect 66260 36907 66312 36916
rect 66260 36873 66269 36907
rect 66269 36873 66303 36907
rect 66303 36873 66312 36907
rect 66260 36864 66312 36873
rect 66996 36864 67048 36916
rect 67640 36864 67692 36916
rect 68284 36864 68336 36916
rect 68928 36864 68980 36916
rect 69572 36864 69624 36916
rect 70216 36864 70268 36916
rect 70860 36864 70912 36916
rect 71504 36864 71556 36916
rect 72148 36864 72200 36916
rect 72792 36864 72844 36916
rect 73436 36864 73488 36916
rect 35440 36728 35492 36780
rect 36360 36796 36412 36848
rect 36820 36796 36872 36848
rect 40408 36796 40460 36848
rect 44916 36796 44968 36848
rect 2136 36660 2188 36712
rect 32220 36703 32272 36712
rect 32220 36669 32229 36703
rect 32229 36669 32263 36703
rect 32263 36669 32272 36703
rect 32220 36660 32272 36669
rect 33232 36703 33284 36712
rect 33232 36669 33241 36703
rect 33241 36669 33275 36703
rect 33275 36669 33284 36703
rect 33232 36660 33284 36669
rect 33876 36703 33928 36712
rect 33876 36669 33885 36703
rect 33885 36669 33919 36703
rect 33919 36669 33928 36703
rect 33876 36660 33928 36669
rect 34152 36703 34204 36712
rect 34152 36669 34161 36703
rect 34161 36669 34195 36703
rect 34195 36669 34204 36703
rect 34152 36660 34204 36669
rect 37464 36728 37516 36780
rect 40500 36771 40552 36780
rect 40500 36737 40509 36771
rect 40509 36737 40543 36771
rect 40543 36737 40552 36771
rect 40500 36728 40552 36737
rect 40868 36771 40920 36780
rect 40868 36737 40877 36771
rect 40877 36737 40911 36771
rect 40911 36737 40920 36771
rect 40868 36728 40920 36737
rect 42524 36728 42576 36780
rect 43076 36771 43128 36780
rect 43076 36737 43085 36771
rect 43085 36737 43119 36771
rect 43119 36737 43128 36771
rect 43076 36728 43128 36737
rect 45008 36771 45060 36780
rect 45008 36737 45017 36771
rect 45017 36737 45051 36771
rect 45051 36737 45060 36771
rect 45008 36728 45060 36737
rect 36176 36660 36228 36712
rect 38476 36703 38528 36712
rect 38476 36669 38485 36703
rect 38485 36669 38519 36703
rect 38519 36669 38528 36703
rect 38476 36660 38528 36669
rect 42248 36660 42300 36712
rect 43536 36660 43588 36712
rect 45928 36771 45980 36780
rect 45928 36737 45937 36771
rect 45937 36737 45971 36771
rect 45971 36737 45980 36771
rect 45928 36728 45980 36737
rect 47768 36728 47820 36780
rect 48780 36771 48832 36780
rect 48780 36737 48789 36771
rect 48789 36737 48823 36771
rect 48823 36737 48832 36771
rect 48780 36728 48832 36737
rect 52920 36728 52972 36780
rect 53288 36771 53340 36780
rect 53288 36737 53297 36771
rect 53297 36737 53331 36771
rect 53331 36737 53340 36771
rect 53288 36728 53340 36737
rect 58072 36728 58124 36780
rect 60648 36771 60700 36780
rect 60648 36737 60657 36771
rect 60657 36737 60691 36771
rect 60691 36737 60700 36771
rect 60648 36728 60700 36737
rect 61016 36771 61068 36780
rect 61016 36737 61025 36771
rect 61025 36737 61059 36771
rect 61059 36737 61068 36771
rect 61016 36728 61068 36737
rect 63132 36728 63184 36780
rect 68284 36728 68336 36780
rect 72240 36771 72292 36780
rect 72240 36737 72249 36771
rect 72249 36737 72283 36771
rect 72283 36737 72292 36771
rect 72240 36728 72292 36737
rect 36084 36592 36136 36644
rect 33508 36524 33560 36576
rect 35716 36524 35768 36576
rect 37280 36524 37332 36576
rect 39488 36524 39540 36576
rect 44548 36524 44600 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 1308 36320 1360 36372
rect 32220 36320 32272 36372
rect 34152 36320 34204 36372
rect 34704 36295 34756 36304
rect 34704 36261 34713 36295
rect 34713 36261 34747 36295
rect 34747 36261 34756 36295
rect 34704 36252 34756 36261
rect 38476 36320 38528 36372
rect 39212 36320 39264 36372
rect 42524 36363 42576 36372
rect 42524 36329 42533 36363
rect 42533 36329 42567 36363
rect 42567 36329 42576 36363
rect 42524 36320 42576 36329
rect 43076 36363 43128 36372
rect 43076 36329 43085 36363
rect 43085 36329 43119 36363
rect 43119 36329 43128 36363
rect 43076 36320 43128 36329
rect 43536 36363 43588 36372
rect 43536 36329 43545 36363
rect 43545 36329 43579 36363
rect 43579 36329 43588 36363
rect 43536 36320 43588 36329
rect 43720 36363 43772 36372
rect 43720 36329 43729 36363
rect 43729 36329 43763 36363
rect 43763 36329 43772 36363
rect 43720 36320 43772 36329
rect 44364 36363 44416 36372
rect 44364 36329 44373 36363
rect 44373 36329 44407 36363
rect 44407 36329 44416 36363
rect 44364 36320 44416 36329
rect 45008 36320 45060 36372
rect 47768 36363 47820 36372
rect 47768 36329 47777 36363
rect 47777 36329 47811 36363
rect 47811 36329 47820 36363
rect 47768 36320 47820 36329
rect 48780 36363 48832 36372
rect 48780 36329 48789 36363
rect 48789 36329 48823 36363
rect 48823 36329 48832 36363
rect 48780 36320 48832 36329
rect 52920 36363 52972 36372
rect 52920 36329 52929 36363
rect 52929 36329 52963 36363
rect 52963 36329 52972 36363
rect 52920 36320 52972 36329
rect 53288 36363 53340 36372
rect 53288 36329 53297 36363
rect 53297 36329 53331 36363
rect 53331 36329 53340 36363
rect 53288 36320 53340 36329
rect 58072 36363 58124 36372
rect 58072 36329 58081 36363
rect 58081 36329 58115 36363
rect 58115 36329 58124 36363
rect 58072 36320 58124 36329
rect 60648 36363 60700 36372
rect 60648 36329 60657 36363
rect 60657 36329 60691 36363
rect 60691 36329 60700 36363
rect 60648 36320 60700 36329
rect 61016 36363 61068 36372
rect 61016 36329 61025 36363
rect 61025 36329 61059 36363
rect 61059 36329 61068 36363
rect 61016 36320 61068 36329
rect 63132 36363 63184 36372
rect 63132 36329 63141 36363
rect 63141 36329 63175 36363
rect 63175 36329 63184 36363
rect 63132 36320 63184 36329
rect 68284 36363 68336 36372
rect 68284 36329 68293 36363
rect 68293 36329 68327 36363
rect 68327 36329 68336 36363
rect 68284 36320 68336 36329
rect 72240 36363 72292 36372
rect 72240 36329 72249 36363
rect 72249 36329 72283 36363
rect 72283 36329 72292 36363
rect 72240 36320 72292 36329
rect 33508 36227 33560 36236
rect 33508 36193 33517 36227
rect 33517 36193 33551 36227
rect 33551 36193 33560 36227
rect 33508 36184 33560 36193
rect 33876 36184 33928 36236
rect 36176 36227 36228 36236
rect 36176 36193 36185 36227
rect 36185 36193 36219 36227
rect 36219 36193 36228 36227
rect 36176 36184 36228 36193
rect 39028 36252 39080 36304
rect 38200 36184 38252 36236
rect 2136 36159 2188 36168
rect 2136 36125 2145 36159
rect 2145 36125 2179 36159
rect 2179 36125 2188 36159
rect 2136 36116 2188 36125
rect 35164 36159 35216 36168
rect 35164 36125 35173 36159
rect 35173 36125 35207 36159
rect 35207 36125 35216 36159
rect 35164 36116 35216 36125
rect 940 35980 992 36032
rect 35716 36048 35768 36100
rect 36084 36159 36136 36168
rect 36084 36125 36093 36159
rect 36093 36125 36127 36159
rect 36127 36125 36136 36159
rect 36084 36116 36136 36125
rect 36728 36048 36780 36100
rect 37464 36048 37516 36100
rect 34612 35980 34664 36032
rect 36360 35980 36412 36032
rect 39028 36116 39080 36168
rect 39212 36159 39264 36168
rect 39212 36125 39221 36159
rect 39221 36125 39255 36159
rect 39255 36125 39264 36159
rect 39212 36116 39264 36125
rect 42248 36227 42300 36236
rect 42248 36193 42257 36227
rect 42257 36193 42291 36227
rect 42291 36193 42300 36227
rect 42248 36184 42300 36193
rect 45744 36184 45796 36236
rect 44088 36159 44140 36168
rect 44088 36125 44097 36159
rect 44097 36125 44131 36159
rect 44131 36125 44140 36159
rect 44088 36116 44140 36125
rect 44364 36116 44416 36168
rect 46112 36159 46164 36168
rect 46112 36125 46121 36159
rect 46121 36125 46155 36159
rect 46155 36125 46164 36159
rect 46112 36116 46164 36125
rect 46480 36116 46532 36168
rect 38384 36048 38436 36100
rect 38016 36023 38068 36032
rect 38016 35989 38025 36023
rect 38025 35989 38059 36023
rect 38059 35989 38068 36023
rect 38016 35980 38068 35989
rect 39120 36023 39172 36032
rect 39120 35989 39129 36023
rect 39129 35989 39163 36023
rect 39163 35989 39172 36023
rect 39120 35980 39172 35989
rect 39488 36091 39540 36100
rect 39488 36057 39497 36091
rect 39497 36057 39531 36091
rect 39531 36057 39540 36091
rect 39488 36048 39540 36057
rect 40408 36048 40460 36100
rect 41972 36091 42024 36100
rect 41972 36057 41981 36091
rect 41981 36057 42015 36091
rect 42015 36057 42024 36091
rect 41972 36048 42024 36057
rect 40684 35980 40736 36032
rect 44272 35980 44324 36032
rect 45928 36023 45980 36032
rect 45928 35989 45937 36023
rect 45937 35989 45971 36023
rect 45971 35989 45980 36023
rect 45928 35980 45980 35989
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 66314 35878 66366 35930
rect 66378 35878 66430 35930
rect 66442 35878 66494 35930
rect 66506 35878 66558 35930
rect 66570 35878 66622 35930
rect 32680 35776 32732 35828
rect 33232 35776 33284 35828
rect 35164 35776 35216 35828
rect 35348 35776 35400 35828
rect 36268 35776 36320 35828
rect 36820 35819 36872 35828
rect 36820 35785 36829 35819
rect 36829 35785 36863 35819
rect 36863 35785 36872 35819
rect 36820 35776 36872 35785
rect 32404 35640 32456 35692
rect 38016 35708 38068 35760
rect 39120 35776 39172 35828
rect 41972 35776 42024 35828
rect 44272 35776 44324 35828
rect 46480 35776 46532 35828
rect 41328 35751 41380 35760
rect 32772 35683 32824 35692
rect 32772 35649 32781 35683
rect 32781 35649 32815 35683
rect 32815 35649 32824 35683
rect 32772 35640 32824 35649
rect 36360 35640 36412 35692
rect 37280 35640 37332 35692
rect 38200 35683 38252 35692
rect 38200 35649 38209 35683
rect 38209 35649 38243 35683
rect 38243 35649 38252 35683
rect 38200 35640 38252 35649
rect 38384 35683 38436 35692
rect 38384 35649 38393 35683
rect 38393 35649 38427 35683
rect 38427 35649 38436 35683
rect 38384 35640 38436 35649
rect 41328 35717 41337 35751
rect 41337 35717 41371 35751
rect 41371 35717 41380 35751
rect 41328 35708 41380 35717
rect 43720 35708 43772 35760
rect 40684 35640 40736 35692
rect 40868 35683 40920 35692
rect 40868 35649 40877 35683
rect 40877 35649 40911 35683
rect 40911 35649 40920 35683
rect 40868 35640 40920 35649
rect 44548 35683 44600 35692
rect 44548 35649 44557 35683
rect 44557 35649 44591 35683
rect 44591 35649 44600 35683
rect 44548 35640 44600 35649
rect 44732 35683 44784 35692
rect 44732 35649 44741 35683
rect 44741 35649 44775 35683
rect 44775 35649 44784 35683
rect 44732 35640 44784 35649
rect 45744 35708 45796 35760
rect 45928 35708 45980 35760
rect 42248 35572 42300 35624
rect 45928 35572 45980 35624
rect 36728 35504 36780 35556
rect 940 35436 992 35488
rect 31484 35436 31536 35488
rect 48780 35436 48832 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 34704 35275 34756 35284
rect 34704 35241 34713 35275
rect 34713 35241 34747 35275
rect 34747 35241 34756 35275
rect 34704 35232 34756 35241
rect 44732 35232 44784 35284
rect 43720 35164 43772 35216
rect 28632 35096 28684 35148
rect 28724 35139 28776 35148
rect 28724 35105 28733 35139
rect 28733 35105 28767 35139
rect 28767 35105 28776 35139
rect 28724 35096 28776 35105
rect 31484 35139 31536 35148
rect 31484 35105 31493 35139
rect 31493 35105 31527 35139
rect 31527 35105 31536 35139
rect 31484 35096 31536 35105
rect 36176 35096 36228 35148
rect 44088 35096 44140 35148
rect 29920 35028 29972 35080
rect 30196 35028 30248 35080
rect 31576 34960 31628 35012
rect 35440 35028 35492 35080
rect 38568 35028 38620 35080
rect 43352 35071 43404 35080
rect 43352 35037 43361 35071
rect 43361 35037 43395 35071
rect 43395 35037 43404 35071
rect 43352 35028 43404 35037
rect 43536 35071 43588 35080
rect 43536 35037 43545 35071
rect 43545 35037 43579 35071
rect 43579 35037 43588 35071
rect 43536 35028 43588 35037
rect 44272 35028 44324 35080
rect 46112 35232 46164 35284
rect 46480 35096 46532 35148
rect 36268 34960 36320 35012
rect 44640 34960 44692 35012
rect 2044 34935 2096 34944
rect 2044 34901 2053 34935
rect 2053 34901 2087 34935
rect 2087 34901 2096 34935
rect 2044 34892 2096 34901
rect 32496 34892 32548 34944
rect 32772 34892 32824 34944
rect 34520 34892 34572 34944
rect 35256 34892 35308 34944
rect 38752 34892 38804 34944
rect 42800 34892 42852 34944
rect 44088 34892 44140 34944
rect 45744 34892 45796 34944
rect 46848 35028 46900 35080
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 66314 34790 66366 34842
rect 66378 34790 66430 34842
rect 66442 34790 66494 34842
rect 66506 34790 66558 34842
rect 66570 34790 66622 34842
rect 1308 34688 1360 34740
rect 2044 34595 2096 34604
rect 2044 34561 2053 34595
rect 2053 34561 2087 34595
rect 2087 34561 2096 34595
rect 2044 34552 2096 34561
rect 30196 34688 30248 34740
rect 34612 34688 34664 34740
rect 28724 34663 28776 34672
rect 28724 34629 28733 34663
rect 28733 34629 28767 34663
rect 28767 34629 28776 34663
rect 28724 34620 28776 34629
rect 2136 34527 2188 34536
rect 2136 34493 2145 34527
rect 2145 34493 2179 34527
rect 2179 34493 2188 34527
rect 2136 34484 2188 34493
rect 31576 34620 31628 34672
rect 32220 34552 32272 34604
rect 33876 34620 33928 34672
rect 36176 34688 36228 34740
rect 36268 34731 36320 34740
rect 36268 34697 36277 34731
rect 36277 34697 36311 34731
rect 36311 34697 36320 34731
rect 36268 34688 36320 34697
rect 35256 34620 35308 34672
rect 35348 34620 35400 34672
rect 35532 34552 35584 34604
rect 28356 34416 28408 34468
rect 29736 34416 29788 34468
rect 29920 34348 29972 34400
rect 32312 34527 32364 34536
rect 32312 34493 32321 34527
rect 32321 34493 32355 34527
rect 32355 34493 32364 34527
rect 32312 34484 32364 34493
rect 32496 34527 32548 34536
rect 32496 34493 32505 34527
rect 32505 34493 32539 34527
rect 32539 34493 32548 34527
rect 32496 34484 32548 34493
rect 32588 34527 32640 34536
rect 32588 34493 32597 34527
rect 32597 34493 32631 34527
rect 32631 34493 32640 34527
rect 32588 34484 32640 34493
rect 35348 34484 35400 34536
rect 38200 34552 38252 34604
rect 40408 34552 40460 34604
rect 41236 34552 41288 34604
rect 42800 34620 42852 34672
rect 45836 34688 45888 34740
rect 44640 34620 44692 34672
rect 42248 34552 42300 34604
rect 44272 34552 44324 34604
rect 46112 34552 46164 34604
rect 31944 34348 31996 34400
rect 34520 34348 34572 34400
rect 37280 34391 37332 34400
rect 37280 34357 37289 34391
rect 37289 34357 37323 34391
rect 37323 34357 37332 34391
rect 37280 34348 37332 34357
rect 39488 34348 39540 34400
rect 40040 34348 40092 34400
rect 44272 34348 44324 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 38200 34144 38252 34196
rect 39120 34144 39172 34196
rect 39488 34187 39540 34196
rect 39488 34153 39497 34187
rect 39497 34153 39531 34187
rect 39531 34153 39540 34187
rect 39488 34144 39540 34153
rect 41144 34144 41196 34196
rect 43352 34187 43404 34196
rect 43352 34153 43361 34187
rect 43361 34153 43395 34187
rect 43395 34153 43404 34187
rect 43352 34144 43404 34153
rect 940 34076 992 34128
rect 28448 34076 28500 34128
rect 30196 34051 30248 34060
rect 30196 34017 30205 34051
rect 30205 34017 30239 34051
rect 30239 34017 30248 34051
rect 30196 34008 30248 34017
rect 2136 33940 2188 33992
rect 26976 33983 27028 33992
rect 26976 33949 26985 33983
rect 26985 33949 27019 33983
rect 27019 33949 27028 33983
rect 26976 33940 27028 33949
rect 28356 33940 28408 33992
rect 28632 33940 28684 33992
rect 29736 33940 29788 33992
rect 31576 33940 31628 33992
rect 32220 33940 32272 33992
rect 32588 34008 32640 34060
rect 35532 34076 35584 34128
rect 38568 34076 38620 34128
rect 45100 34076 45152 34128
rect 37280 34008 37332 34060
rect 40960 34008 41012 34060
rect 27252 33915 27304 33924
rect 27252 33881 27261 33915
rect 27261 33881 27295 33915
rect 27295 33881 27304 33915
rect 27252 33872 27304 33881
rect 29092 33915 29144 33924
rect 29092 33881 29101 33915
rect 29101 33881 29135 33915
rect 29135 33881 29144 33915
rect 29092 33872 29144 33881
rect 30380 33872 30432 33924
rect 29460 33804 29512 33856
rect 32036 33847 32088 33856
rect 32036 33813 32045 33847
rect 32045 33813 32079 33847
rect 32079 33813 32088 33847
rect 32036 33804 32088 33813
rect 32312 33804 32364 33856
rect 32404 33804 32456 33856
rect 35348 33940 35400 33992
rect 35532 33983 35584 33992
rect 35532 33949 35541 33983
rect 35541 33949 35575 33983
rect 35575 33949 35584 33983
rect 35532 33940 35584 33949
rect 33048 33872 33100 33924
rect 35256 33915 35308 33924
rect 35256 33881 35265 33915
rect 35265 33881 35299 33915
rect 35299 33881 35308 33915
rect 35256 33872 35308 33881
rect 33692 33804 33744 33856
rect 35440 33804 35492 33856
rect 36084 33983 36136 33992
rect 36084 33949 36093 33983
rect 36093 33949 36127 33983
rect 36127 33949 36136 33983
rect 36084 33940 36136 33949
rect 36176 33940 36228 33992
rect 38936 33983 38988 33992
rect 38936 33949 38945 33983
rect 38945 33949 38979 33983
rect 38979 33949 38988 33983
rect 38936 33940 38988 33949
rect 39948 33940 40000 33992
rect 40868 33983 40920 33992
rect 40868 33949 40877 33983
rect 40877 33949 40911 33983
rect 40911 33949 40920 33983
rect 40868 33940 40920 33949
rect 41052 33940 41104 33992
rect 37372 33872 37424 33924
rect 40040 33915 40092 33924
rect 40040 33881 40049 33915
rect 40049 33881 40083 33915
rect 40083 33881 40092 33915
rect 41328 33940 41380 33992
rect 42432 33940 42484 33992
rect 43536 33940 43588 33992
rect 40040 33872 40092 33881
rect 36360 33804 36412 33856
rect 40684 33804 40736 33856
rect 42156 33872 42208 33924
rect 44272 33804 44324 33856
rect 45100 33847 45152 33856
rect 45100 33813 45109 33847
rect 45109 33813 45143 33847
rect 45143 33813 45152 33847
rect 45100 33804 45152 33813
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 66314 33702 66366 33754
rect 66378 33702 66430 33754
rect 66442 33702 66494 33754
rect 66506 33702 66558 33754
rect 66570 33702 66622 33754
rect 27252 33600 27304 33652
rect 29092 33600 29144 33652
rect 29000 33532 29052 33584
rect 30380 33643 30432 33652
rect 30380 33609 30389 33643
rect 30389 33609 30423 33643
rect 30423 33609 30432 33643
rect 30380 33600 30432 33609
rect 38936 33600 38988 33652
rect 39948 33600 40000 33652
rect 28448 33507 28500 33516
rect 28448 33473 28457 33507
rect 28457 33473 28491 33507
rect 28491 33473 28500 33507
rect 28448 33464 28500 33473
rect 28632 33464 28684 33516
rect 29920 33575 29972 33584
rect 29920 33541 29929 33575
rect 29929 33541 29963 33575
rect 29963 33541 29972 33575
rect 29920 33532 29972 33541
rect 32220 33532 32272 33584
rect 35256 33532 35308 33584
rect 32036 33464 32088 33516
rect 32404 33464 32456 33516
rect 32588 33464 32640 33516
rect 35440 33507 35492 33516
rect 35440 33473 35449 33507
rect 35449 33473 35483 33507
rect 35483 33473 35492 33507
rect 35440 33464 35492 33473
rect 35992 33464 36044 33516
rect 36360 33507 36412 33516
rect 36360 33473 36369 33507
rect 36369 33473 36403 33507
rect 36403 33473 36412 33507
rect 36360 33464 36412 33473
rect 29460 33439 29512 33448
rect 29460 33405 29469 33439
rect 29469 33405 29503 33439
rect 29503 33405 29512 33439
rect 29460 33396 29512 33405
rect 36084 33396 36136 33448
rect 37004 33464 37056 33516
rect 38108 33507 38160 33516
rect 38108 33473 38117 33507
rect 38117 33473 38151 33507
rect 38151 33473 38160 33507
rect 38108 33464 38160 33473
rect 39488 33532 39540 33584
rect 39212 33396 39264 33448
rect 40868 33600 40920 33652
rect 40684 33575 40736 33584
rect 40684 33541 40693 33575
rect 40693 33541 40727 33575
rect 40727 33541 40736 33575
rect 41052 33600 41104 33652
rect 40684 33532 40736 33541
rect 43812 33600 43864 33652
rect 44180 33600 44232 33652
rect 40960 33464 41012 33516
rect 41328 33464 41380 33516
rect 42156 33507 42208 33516
rect 42156 33473 42165 33507
rect 42165 33473 42199 33507
rect 42199 33473 42208 33507
rect 42156 33464 42208 33473
rect 42432 33507 42484 33516
rect 42432 33473 42441 33507
rect 42441 33473 42475 33507
rect 42475 33473 42484 33507
rect 42432 33464 42484 33473
rect 44272 33507 44324 33516
rect 44272 33473 44281 33507
rect 44281 33473 44315 33507
rect 44315 33473 44324 33507
rect 44272 33464 44324 33473
rect 45928 33600 45980 33652
rect 46112 33643 46164 33652
rect 46112 33609 46121 33643
rect 46121 33609 46155 33643
rect 46155 33609 46164 33643
rect 46112 33600 46164 33609
rect 46204 33600 46256 33652
rect 45100 33575 45152 33584
rect 45100 33541 45109 33575
rect 45109 33541 45143 33575
rect 45143 33541 45152 33575
rect 45100 33532 45152 33541
rect 44732 33464 44784 33516
rect 940 33328 992 33380
rect 31944 33328 31996 33380
rect 41604 33328 41656 33380
rect 29736 33303 29788 33312
rect 29736 33269 29745 33303
rect 29745 33269 29779 33303
rect 29779 33269 29788 33303
rect 29736 33260 29788 33269
rect 32036 33260 32088 33312
rect 33048 33260 33100 33312
rect 37280 33260 37332 33312
rect 37740 33260 37792 33312
rect 39672 33303 39724 33312
rect 39672 33269 39681 33303
rect 39681 33269 39715 33303
rect 39715 33269 39724 33303
rect 39672 33260 39724 33269
rect 39856 33303 39908 33312
rect 39856 33269 39865 33303
rect 39865 33269 39899 33303
rect 39899 33269 39908 33303
rect 39856 33260 39908 33269
rect 40592 33260 40644 33312
rect 41144 33303 41196 33312
rect 41144 33269 41153 33303
rect 41153 33269 41187 33303
rect 41187 33269 41196 33303
rect 41144 33260 41196 33269
rect 46388 33507 46440 33516
rect 46388 33473 46397 33507
rect 46397 33473 46431 33507
rect 46431 33473 46440 33507
rect 46388 33464 46440 33473
rect 47676 33532 47728 33584
rect 48780 33532 48832 33584
rect 46020 33396 46072 33448
rect 46848 33464 46900 33516
rect 44732 33328 44784 33380
rect 45192 33328 45244 33380
rect 47768 33439 47820 33448
rect 47768 33405 47777 33439
rect 47777 33405 47811 33439
rect 47811 33405 47820 33439
rect 47768 33396 47820 33405
rect 48044 33439 48096 33448
rect 48044 33405 48053 33439
rect 48053 33405 48087 33439
rect 48087 33405 48096 33439
rect 48044 33396 48096 33405
rect 42156 33260 42208 33312
rect 44640 33303 44692 33312
rect 44640 33269 44649 33303
rect 44649 33269 44683 33303
rect 44683 33269 44692 33303
rect 44640 33260 44692 33269
rect 46020 33260 46072 33312
rect 47492 33260 47544 33312
rect 47676 33260 47728 33312
rect 49608 33260 49660 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 30288 33056 30340 33108
rect 33968 33056 34020 33108
rect 36360 33056 36412 33108
rect 36912 33056 36964 33108
rect 37004 33099 37056 33108
rect 37004 33065 37013 33099
rect 37013 33065 37047 33099
rect 37047 33065 37056 33099
rect 37004 33056 37056 33065
rect 38108 33056 38160 33108
rect 38936 33056 38988 33108
rect 40684 33056 40736 33108
rect 43812 33099 43864 33108
rect 43812 33065 43821 33099
rect 43821 33065 43855 33099
rect 43855 33065 43864 33099
rect 43812 33056 43864 33065
rect 44272 33056 44324 33108
rect 29000 32920 29052 32972
rect 30196 32920 30248 32972
rect 33048 32963 33100 32972
rect 33048 32929 33057 32963
rect 33057 32929 33091 32963
rect 33091 32929 33100 32963
rect 33048 32920 33100 32929
rect 29184 32895 29236 32904
rect 29184 32861 29193 32895
rect 29193 32861 29227 32895
rect 29227 32861 29236 32895
rect 29184 32852 29236 32861
rect 32036 32895 32088 32904
rect 32036 32861 32045 32895
rect 32045 32861 32079 32895
rect 32079 32861 32088 32895
rect 32036 32852 32088 32861
rect 32128 32895 32180 32904
rect 32128 32861 32137 32895
rect 32137 32861 32171 32895
rect 32171 32861 32180 32895
rect 32128 32852 32180 32861
rect 33692 32895 33744 32904
rect 33692 32861 33701 32895
rect 33701 32861 33735 32895
rect 33735 32861 33744 32895
rect 33692 32852 33744 32861
rect 39212 33031 39264 33040
rect 39212 32997 39221 33031
rect 39221 32997 39255 33031
rect 39255 32997 39264 33031
rect 39212 32988 39264 32997
rect 36176 32920 36228 32972
rect 37740 32963 37792 32972
rect 37740 32929 37749 32963
rect 37749 32929 37783 32963
rect 37783 32929 37792 32963
rect 37740 32920 37792 32929
rect 38752 32920 38804 32972
rect 29368 32784 29420 32836
rect 940 32716 992 32768
rect 27988 32716 28040 32768
rect 35348 32716 35400 32768
rect 37096 32895 37148 32904
rect 37096 32861 37105 32895
rect 37105 32861 37139 32895
rect 37139 32861 37148 32895
rect 37096 32852 37148 32861
rect 39488 32895 39540 32904
rect 39488 32861 39497 32895
rect 39497 32861 39531 32895
rect 39531 32861 39540 32895
rect 39488 32852 39540 32861
rect 39856 32920 39908 32972
rect 42248 32920 42300 32972
rect 42708 32920 42760 32972
rect 45192 33099 45244 33108
rect 45192 33065 45201 33099
rect 45201 33065 45235 33099
rect 45235 33065 45244 33099
rect 45192 33056 45244 33065
rect 45376 32988 45428 33040
rect 41236 32852 41288 32904
rect 44548 32852 44600 32904
rect 45192 32920 45244 32972
rect 48044 33056 48096 33108
rect 46848 32988 46900 33040
rect 45928 32920 45980 32972
rect 44732 32852 44784 32904
rect 45376 32852 45428 32904
rect 46020 32852 46072 32904
rect 39672 32716 39724 32768
rect 39948 32759 40000 32768
rect 39948 32725 39957 32759
rect 39957 32725 39991 32759
rect 39991 32725 40000 32759
rect 39948 32716 40000 32725
rect 41604 32716 41656 32768
rect 44364 32759 44416 32768
rect 44364 32725 44373 32759
rect 44373 32725 44407 32759
rect 44407 32725 44416 32759
rect 44364 32716 44416 32725
rect 44456 32716 44508 32768
rect 46204 32784 46256 32836
rect 47768 32920 47820 32972
rect 48780 32920 48832 32972
rect 49608 32920 49660 32972
rect 47216 32895 47268 32904
rect 47216 32861 47225 32895
rect 47225 32861 47259 32895
rect 47259 32861 47268 32895
rect 47216 32852 47268 32861
rect 47308 32895 47360 32904
rect 47308 32861 47317 32895
rect 47317 32861 47351 32895
rect 47351 32861 47360 32895
rect 47308 32852 47360 32861
rect 47492 32895 47544 32904
rect 47492 32861 47501 32895
rect 47501 32861 47535 32895
rect 47535 32861 47544 32895
rect 47492 32852 47544 32861
rect 47584 32895 47636 32904
rect 47584 32861 47593 32895
rect 47593 32861 47627 32895
rect 47627 32861 47636 32895
rect 47584 32852 47636 32861
rect 47676 32895 47728 32904
rect 47676 32861 47685 32895
rect 47685 32861 47719 32895
rect 47719 32861 47728 32895
rect 47676 32852 47728 32861
rect 48780 32784 48832 32836
rect 46112 32716 46164 32768
rect 46572 32759 46624 32768
rect 46572 32725 46599 32759
rect 46599 32725 46624 32759
rect 46572 32716 46624 32725
rect 49792 32759 49844 32768
rect 49792 32725 49801 32759
rect 49801 32725 49835 32759
rect 49835 32725 49844 32759
rect 49792 32716 49844 32725
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 66314 32614 66366 32666
rect 66378 32614 66430 32666
rect 66442 32614 66494 32666
rect 66506 32614 66558 32666
rect 66570 32614 66622 32666
rect 17684 32444 17736 32496
rect 18696 32444 18748 32496
rect 27344 32512 27396 32564
rect 30196 32512 30248 32564
rect 30288 32555 30340 32564
rect 30288 32521 30297 32555
rect 30297 32521 30331 32555
rect 30331 32521 30340 32555
rect 30288 32512 30340 32521
rect 33048 32512 33100 32564
rect 33968 32487 34020 32496
rect 33968 32453 33977 32487
rect 33977 32453 34011 32487
rect 34011 32453 34020 32487
rect 33968 32444 34020 32453
rect 28356 32376 28408 32428
rect 29000 32419 29052 32428
rect 29000 32385 29009 32419
rect 29009 32385 29043 32419
rect 29043 32385 29052 32419
rect 29000 32376 29052 32385
rect 29736 32419 29788 32428
rect 29736 32385 29745 32419
rect 29745 32385 29779 32419
rect 29779 32385 29788 32419
rect 29736 32376 29788 32385
rect 30012 32376 30064 32428
rect 31300 32419 31352 32428
rect 31300 32385 31309 32419
rect 31309 32385 31343 32419
rect 31343 32385 31352 32419
rect 31300 32376 31352 32385
rect 32864 32376 32916 32428
rect 36176 32512 36228 32564
rect 45192 32555 45244 32564
rect 45192 32521 45201 32555
rect 45201 32521 45235 32555
rect 45235 32521 45244 32555
rect 45192 32512 45244 32521
rect 46388 32512 46440 32564
rect 47584 32555 47636 32564
rect 47584 32521 47593 32555
rect 47593 32521 47627 32555
rect 47627 32521 47636 32555
rect 47584 32512 47636 32521
rect 37372 32444 37424 32496
rect 43812 32376 43864 32428
rect 44180 32376 44232 32428
rect 44456 32419 44508 32428
rect 44456 32385 44465 32419
rect 44465 32385 44499 32419
rect 44499 32385 44508 32419
rect 44456 32376 44508 32385
rect 44640 32419 44692 32428
rect 44640 32385 44649 32419
rect 44649 32385 44683 32419
rect 44683 32385 44692 32419
rect 44640 32376 44692 32385
rect 45560 32487 45612 32496
rect 45560 32453 45569 32487
rect 45569 32453 45603 32487
rect 45603 32453 45612 32487
rect 45560 32444 45612 32453
rect 45928 32444 45980 32496
rect 46020 32487 46072 32496
rect 46020 32453 46061 32487
rect 46061 32453 46072 32487
rect 46020 32444 46072 32453
rect 2044 32351 2096 32360
rect 2044 32317 2053 32351
rect 2053 32317 2087 32351
rect 2087 32317 2096 32351
rect 2044 32308 2096 32317
rect 17408 32351 17460 32360
rect 17408 32317 17417 32351
rect 17417 32317 17451 32351
rect 17451 32317 17460 32351
rect 17408 32308 17460 32317
rect 27252 32351 27304 32360
rect 27252 32317 27261 32351
rect 27261 32317 27295 32351
rect 27295 32317 27304 32351
rect 27252 32308 27304 32317
rect 29184 32351 29236 32360
rect 29184 32317 29193 32351
rect 29193 32317 29227 32351
rect 29227 32317 29236 32351
rect 29184 32308 29236 32317
rect 29920 32308 29972 32360
rect 30380 32351 30432 32360
rect 30380 32317 30389 32351
rect 30389 32317 30423 32351
rect 30423 32317 30432 32351
rect 30380 32308 30432 32317
rect 34704 32308 34756 32360
rect 35992 32308 36044 32360
rect 39672 32308 39724 32360
rect 46572 32308 46624 32360
rect 47216 32444 47268 32496
rect 47768 32419 47820 32428
rect 47768 32385 47777 32419
rect 47777 32385 47811 32419
rect 47811 32385 47820 32419
rect 47768 32376 47820 32385
rect 18512 32172 18564 32224
rect 27712 32172 27764 32224
rect 28816 32215 28868 32224
rect 28816 32181 28825 32215
rect 28825 32181 28859 32215
rect 28859 32181 28868 32215
rect 28816 32172 28868 32181
rect 29368 32215 29420 32224
rect 29368 32181 29377 32215
rect 29377 32181 29411 32215
rect 29411 32181 29420 32215
rect 29368 32172 29420 32181
rect 43536 32283 43588 32292
rect 43536 32249 43545 32283
rect 43545 32249 43579 32283
rect 43579 32249 43588 32283
rect 43536 32240 43588 32249
rect 31392 32172 31444 32224
rect 36176 32215 36228 32224
rect 36176 32181 36185 32215
rect 36185 32181 36219 32215
rect 36219 32181 36228 32215
rect 36176 32172 36228 32181
rect 46204 32240 46256 32292
rect 48044 32351 48096 32360
rect 48044 32317 48053 32351
rect 48053 32317 48087 32351
rect 48087 32317 48096 32351
rect 48044 32308 48096 32317
rect 49792 32376 49844 32428
rect 45560 32172 45612 32224
rect 46112 32172 46164 32224
rect 46388 32172 46440 32224
rect 47308 32172 47360 32224
rect 48044 32172 48096 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 1308 31968 1360 32020
rect 17408 31968 17460 32020
rect 27252 31968 27304 32020
rect 30380 31968 30432 32020
rect 31392 32011 31444 32020
rect 31392 31977 31413 32011
rect 31413 31977 31444 32011
rect 31392 31968 31444 31977
rect 34704 32011 34756 32020
rect 34704 31977 34713 32011
rect 34713 31977 34747 32011
rect 34747 31977 34756 32011
rect 34704 31968 34756 31977
rect 35440 31968 35492 32020
rect 44456 31968 44508 32020
rect 46388 31968 46440 32020
rect 47124 31968 47176 32020
rect 47768 31968 47820 32020
rect 28356 31900 28408 31952
rect 2044 31807 2096 31816
rect 2044 31773 2053 31807
rect 2053 31773 2087 31807
rect 2087 31773 2096 31807
rect 2044 31764 2096 31773
rect 11336 31764 11388 31816
rect 15384 31807 15436 31816
rect 15384 31773 15393 31807
rect 15393 31773 15427 31807
rect 15427 31773 15436 31807
rect 15384 31764 15436 31773
rect 17684 31832 17736 31884
rect 21456 31875 21508 31884
rect 21456 31841 21465 31875
rect 21465 31841 21499 31875
rect 21499 31841 21508 31875
rect 21456 31832 21508 31841
rect 26976 31832 27028 31884
rect 12348 31739 12400 31748
rect 12348 31705 12357 31739
rect 12357 31705 12391 31739
rect 12391 31705 12400 31739
rect 12348 31696 12400 31705
rect 13636 31696 13688 31748
rect 14740 31696 14792 31748
rect 16304 31696 16356 31748
rect 18512 31807 18564 31816
rect 18512 31773 18521 31807
rect 18521 31773 18555 31807
rect 18555 31773 18564 31807
rect 18512 31764 18564 31773
rect 18788 31764 18840 31816
rect 27712 31764 27764 31816
rect 27988 31807 28040 31816
rect 27988 31773 27997 31807
rect 27997 31773 28031 31807
rect 28031 31773 28040 31807
rect 27988 31764 28040 31773
rect 28816 31764 28868 31816
rect 44180 31900 44232 31952
rect 44548 31900 44600 31952
rect 30380 31832 30432 31884
rect 36176 31832 36228 31884
rect 40684 31832 40736 31884
rect 44640 31832 44692 31884
rect 17132 31696 17184 31748
rect 20168 31696 20220 31748
rect 30012 31696 30064 31748
rect 2044 31628 2096 31680
rect 13820 31671 13872 31680
rect 13820 31637 13829 31671
rect 13829 31637 13863 31671
rect 13863 31637 13872 31671
rect 13820 31628 13872 31637
rect 15292 31628 15344 31680
rect 29920 31671 29972 31680
rect 29920 31637 29929 31671
rect 29929 31637 29963 31671
rect 29963 31637 29972 31671
rect 29920 31628 29972 31637
rect 35348 31764 35400 31816
rect 37280 31807 37332 31816
rect 37280 31773 37289 31807
rect 37289 31773 37323 31807
rect 37323 31773 37332 31807
rect 37280 31764 37332 31773
rect 41420 31764 41472 31816
rect 41696 31764 41748 31816
rect 43812 31764 43864 31816
rect 44364 31764 44416 31816
rect 45376 31764 45428 31816
rect 46112 31739 46164 31748
rect 46112 31705 46121 31739
rect 46121 31705 46155 31739
rect 46155 31705 46164 31739
rect 46112 31696 46164 31705
rect 46296 31739 46348 31748
rect 46296 31705 46337 31739
rect 46337 31705 46348 31739
rect 46296 31696 46348 31705
rect 46572 31696 46624 31748
rect 30748 31628 30800 31680
rect 36728 31628 36780 31680
rect 39120 31628 39172 31680
rect 40500 31628 40552 31680
rect 45100 31628 45152 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 66314 31526 66366 31578
rect 66378 31526 66430 31578
rect 66442 31526 66494 31578
rect 66506 31526 66558 31578
rect 66570 31526 66622 31578
rect 940 31424 992 31476
rect 11612 31356 11664 31408
rect 13636 31424 13688 31476
rect 15292 31356 15344 31408
rect 16304 31356 16356 31408
rect 18696 31424 18748 31476
rect 28816 31424 28868 31476
rect 30748 31424 30800 31476
rect 20352 31356 20404 31408
rect 30012 31399 30064 31408
rect 2044 31331 2096 31340
rect 2044 31297 2053 31331
rect 2053 31297 2087 31331
rect 2087 31297 2096 31331
rect 2044 31288 2096 31297
rect 11428 31288 11480 31340
rect 17684 31331 17736 31340
rect 17684 31297 17693 31331
rect 17693 31297 17727 31331
rect 17727 31297 17736 31331
rect 17684 31288 17736 31297
rect 29092 31288 29144 31340
rect 30012 31365 30021 31399
rect 30021 31365 30055 31399
rect 30055 31365 30064 31399
rect 30012 31356 30064 31365
rect 35992 31356 36044 31408
rect 36728 31399 36780 31408
rect 36728 31365 36737 31399
rect 36737 31365 36771 31399
rect 36771 31365 36780 31399
rect 36728 31356 36780 31365
rect 37372 31356 37424 31408
rect 37280 31288 37332 31340
rect 40500 31399 40552 31408
rect 40500 31365 40509 31399
rect 40509 31365 40543 31399
rect 40543 31365 40552 31399
rect 40500 31356 40552 31365
rect 40684 31467 40736 31476
rect 40684 31433 40709 31467
rect 40709 31433 40736 31467
rect 40684 31424 40736 31433
rect 40868 31424 40920 31476
rect 42892 31356 42944 31408
rect 44548 31356 44600 31408
rect 9864 31263 9916 31272
rect 9864 31229 9873 31263
rect 9873 31229 9907 31263
rect 9907 31229 9916 31263
rect 9864 31220 9916 31229
rect 11888 31220 11940 31272
rect 12256 31220 12308 31272
rect 13820 31220 13872 31272
rect 18512 31220 18564 31272
rect 18696 31220 18748 31272
rect 27712 31263 27764 31272
rect 27712 31229 27721 31263
rect 27721 31229 27755 31263
rect 27755 31229 27764 31263
rect 27712 31220 27764 31229
rect 29920 31220 29972 31272
rect 31576 31220 31628 31272
rect 29736 31152 29788 31204
rect 31300 31152 31352 31204
rect 9680 31084 9732 31136
rect 11336 31084 11388 31136
rect 11428 31084 11480 31136
rect 12808 31127 12860 31136
rect 12808 31093 12817 31127
rect 12817 31093 12851 31127
rect 12851 31093 12860 31127
rect 12808 31084 12860 31093
rect 13544 31127 13596 31136
rect 13544 31093 13553 31127
rect 13553 31093 13587 31127
rect 13587 31093 13596 31127
rect 13544 31084 13596 31093
rect 16488 31127 16540 31136
rect 16488 31093 16497 31127
rect 16497 31093 16531 31127
rect 16531 31093 16540 31127
rect 16488 31084 16540 31093
rect 16672 31127 16724 31136
rect 16672 31093 16681 31127
rect 16681 31093 16715 31127
rect 16715 31093 16724 31127
rect 16672 31084 16724 31093
rect 19524 31127 19576 31136
rect 19524 31093 19533 31127
rect 19533 31093 19567 31127
rect 19567 31093 19576 31127
rect 19524 31084 19576 31093
rect 20352 31127 20404 31136
rect 20352 31093 20361 31127
rect 20361 31093 20395 31127
rect 20395 31093 20404 31127
rect 20352 31084 20404 31093
rect 27620 31084 27672 31136
rect 29920 31084 29972 31136
rect 36912 31127 36964 31136
rect 36912 31093 36921 31127
rect 36921 31093 36955 31127
rect 36955 31093 36964 31127
rect 36912 31084 36964 31093
rect 37464 31084 37516 31136
rect 38660 31084 38712 31136
rect 40684 31220 40736 31272
rect 41696 31331 41748 31340
rect 41696 31297 41705 31331
rect 41705 31297 41739 31331
rect 41739 31297 41748 31331
rect 41696 31288 41748 31297
rect 42524 31331 42576 31340
rect 42524 31297 42533 31331
rect 42533 31297 42567 31331
rect 42567 31297 42576 31331
rect 42524 31288 42576 31297
rect 44272 31288 44324 31340
rect 46296 31288 46348 31340
rect 46388 31288 46440 31340
rect 46572 31331 46624 31340
rect 46572 31297 46581 31331
rect 46581 31297 46615 31331
rect 46615 31297 46624 31331
rect 46572 31288 46624 31297
rect 47124 31331 47176 31340
rect 47124 31297 47133 31331
rect 47133 31297 47167 31331
rect 47167 31297 47176 31331
rect 47124 31288 47176 31297
rect 46112 31220 46164 31272
rect 46756 31220 46808 31272
rect 40592 31084 40644 31136
rect 40960 31152 41012 31204
rect 47308 31220 47360 31272
rect 40776 31084 40828 31136
rect 42800 31084 42852 31136
rect 45100 31127 45152 31136
rect 45100 31093 45109 31127
rect 45109 31093 45143 31127
rect 45143 31093 45152 31127
rect 45100 31084 45152 31093
rect 45284 31127 45336 31136
rect 45284 31093 45293 31127
rect 45293 31093 45327 31127
rect 45327 31093 45336 31127
rect 45284 31084 45336 31093
rect 47216 31084 47268 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 9864 30880 9916 30932
rect 12348 30880 12400 30932
rect 15384 30880 15436 30932
rect 18512 30923 18564 30932
rect 18512 30889 18521 30923
rect 18521 30889 18555 30923
rect 18555 30889 18564 30923
rect 18512 30880 18564 30889
rect 29092 30923 29144 30932
rect 29092 30889 29101 30923
rect 29101 30889 29135 30923
rect 29135 30889 29144 30923
rect 29092 30880 29144 30889
rect 31576 30923 31628 30932
rect 31576 30889 31585 30923
rect 31585 30889 31619 30923
rect 31619 30889 31628 30923
rect 31576 30880 31628 30889
rect 36912 30880 36964 30932
rect 37372 30880 37424 30932
rect 40684 30923 40736 30932
rect 40684 30889 40693 30923
rect 40693 30889 40727 30923
rect 40727 30889 40736 30923
rect 40684 30880 40736 30889
rect 42524 30880 42576 30932
rect 46756 30923 46808 30932
rect 46756 30889 46765 30923
rect 46765 30889 46799 30923
rect 46799 30889 46808 30923
rect 46756 30880 46808 30889
rect 11704 30787 11756 30796
rect 11704 30753 11713 30787
rect 11713 30753 11747 30787
rect 11747 30753 11756 30787
rect 11704 30744 11756 30753
rect 32128 30812 32180 30864
rect 46572 30812 46624 30864
rect 11244 30719 11296 30728
rect 11244 30685 11253 30719
rect 11253 30685 11287 30719
rect 11287 30685 11296 30719
rect 11244 30676 11296 30685
rect 11428 30719 11480 30728
rect 11428 30685 11437 30719
rect 11437 30685 11471 30719
rect 11471 30685 11480 30719
rect 11428 30676 11480 30685
rect 12808 30676 12860 30728
rect 15200 30719 15252 30728
rect 15200 30685 15209 30719
rect 15209 30685 15243 30719
rect 15243 30685 15252 30719
rect 15200 30676 15252 30685
rect 16672 30676 16724 30728
rect 17132 30719 17184 30728
rect 17132 30685 17141 30719
rect 17141 30685 17175 30719
rect 17175 30685 17184 30719
rect 17132 30676 17184 30685
rect 19524 30744 19576 30796
rect 27344 30787 27396 30796
rect 27344 30753 27353 30787
rect 27353 30753 27387 30787
rect 27387 30753 27396 30787
rect 27344 30744 27396 30753
rect 27620 30787 27672 30796
rect 27620 30753 27629 30787
rect 27629 30753 27663 30787
rect 27663 30753 27672 30787
rect 27620 30744 27672 30753
rect 18420 30676 18472 30728
rect 31300 30676 31352 30728
rect 11704 30608 11756 30660
rect 28356 30608 28408 30660
rect 940 30540 992 30592
rect 15292 30583 15344 30592
rect 15292 30549 15301 30583
rect 15301 30549 15335 30583
rect 15335 30549 15344 30583
rect 15292 30540 15344 30549
rect 17960 30540 18012 30592
rect 30380 30540 30432 30592
rect 32128 30676 32180 30728
rect 34244 30719 34296 30728
rect 34244 30685 34253 30719
rect 34253 30685 34287 30719
rect 34287 30685 34296 30719
rect 34244 30676 34296 30685
rect 37464 30719 37516 30728
rect 37464 30685 37473 30719
rect 37473 30685 37507 30719
rect 37507 30685 37516 30719
rect 37464 30676 37516 30685
rect 37740 30719 37792 30728
rect 32956 30608 33008 30660
rect 33968 30651 34020 30660
rect 33968 30617 33977 30651
rect 33977 30617 34011 30651
rect 34011 30617 34020 30651
rect 33968 30608 34020 30617
rect 33140 30540 33192 30592
rect 36084 30583 36136 30592
rect 36084 30549 36093 30583
rect 36093 30549 36127 30583
rect 36127 30549 36136 30583
rect 36084 30540 36136 30549
rect 36452 30651 36504 30660
rect 36452 30617 36461 30651
rect 36461 30617 36495 30651
rect 36495 30617 36504 30651
rect 37740 30685 37749 30719
rect 37749 30685 37783 30719
rect 37783 30685 37792 30719
rect 37740 30676 37792 30685
rect 37832 30719 37884 30728
rect 37832 30685 37841 30719
rect 37841 30685 37875 30719
rect 37875 30685 37884 30719
rect 37832 30676 37884 30685
rect 42708 30744 42760 30796
rect 47216 30787 47268 30796
rect 47216 30753 47225 30787
rect 47225 30753 47259 30787
rect 47259 30753 47268 30787
rect 47216 30744 47268 30753
rect 40592 30719 40644 30728
rect 40592 30685 40601 30719
rect 40601 30685 40635 30719
rect 40635 30685 40644 30719
rect 40592 30676 40644 30685
rect 36452 30608 36504 30617
rect 36544 30540 36596 30592
rect 37648 30583 37700 30592
rect 37648 30549 37657 30583
rect 37657 30549 37691 30583
rect 37691 30549 37700 30583
rect 37648 30540 37700 30549
rect 37740 30540 37792 30592
rect 40224 30608 40276 30660
rect 41236 30608 41288 30660
rect 43076 30651 43128 30660
rect 43076 30617 43085 30651
rect 43085 30617 43119 30651
rect 43119 30617 43128 30651
rect 43076 30608 43128 30617
rect 45284 30651 45336 30660
rect 45284 30617 45293 30651
rect 45293 30617 45327 30651
rect 45327 30617 45336 30651
rect 45284 30608 45336 30617
rect 46940 30608 46992 30660
rect 43628 30540 43680 30592
rect 48228 30540 48280 30592
rect 48780 30583 48832 30592
rect 48780 30549 48789 30583
rect 48789 30549 48823 30583
rect 48823 30549 48832 30583
rect 48780 30540 48832 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 66314 30438 66366 30490
rect 66378 30438 66430 30490
rect 66442 30438 66494 30490
rect 66506 30438 66558 30490
rect 66570 30438 66622 30490
rect 11244 30336 11296 30388
rect 13544 30336 13596 30388
rect 15200 30336 15252 30388
rect 17960 30336 18012 30388
rect 18788 30336 18840 30388
rect 11888 30243 11940 30252
rect 11888 30209 11897 30243
rect 11897 30209 11931 30243
rect 11931 30209 11940 30243
rect 15476 30268 15528 30320
rect 11888 30200 11940 30209
rect 12532 30243 12584 30252
rect 12532 30209 12541 30243
rect 12541 30209 12575 30243
rect 12575 30209 12584 30243
rect 12532 30200 12584 30209
rect 11704 30064 11756 30116
rect 12256 30107 12308 30116
rect 12256 30073 12265 30107
rect 12265 30073 12299 30107
rect 12299 30073 12308 30107
rect 12256 30064 12308 30073
rect 13084 30064 13136 30116
rect 13360 30107 13412 30116
rect 13360 30073 13369 30107
rect 13369 30073 13403 30107
rect 13403 30073 13412 30107
rect 13360 30064 13412 30073
rect 940 29996 992 30048
rect 13544 30243 13596 30252
rect 13544 30209 13553 30243
rect 13553 30209 13587 30243
rect 13587 30209 13596 30243
rect 13544 30200 13596 30209
rect 15200 30200 15252 30252
rect 18696 30268 18748 30320
rect 16488 30200 16540 30252
rect 17408 30243 17460 30252
rect 17408 30209 17417 30243
rect 17417 30209 17451 30243
rect 17451 30209 17460 30243
rect 17408 30200 17460 30209
rect 18420 30243 18472 30252
rect 18420 30209 18429 30243
rect 18429 30209 18463 30243
rect 18463 30209 18472 30243
rect 18420 30200 18472 30209
rect 29736 30200 29788 30252
rect 30380 30200 30432 30252
rect 32956 30268 33008 30320
rect 35992 30268 36044 30320
rect 39948 30336 40000 30388
rect 40224 30268 40276 30320
rect 40776 30268 40828 30320
rect 43076 30379 43128 30388
rect 43076 30345 43085 30379
rect 43085 30345 43119 30379
rect 43119 30345 43128 30379
rect 43076 30336 43128 30345
rect 44916 30268 44968 30320
rect 32128 30243 32180 30252
rect 32128 30209 32137 30243
rect 32137 30209 32171 30243
rect 32171 30209 32180 30243
rect 32128 30200 32180 30209
rect 14556 30175 14608 30184
rect 14556 30141 14565 30175
rect 14565 30141 14599 30175
rect 14599 30141 14608 30175
rect 14556 30132 14608 30141
rect 19064 30132 19116 30184
rect 31300 30132 31352 30184
rect 17132 30064 17184 30116
rect 28356 30064 28408 30116
rect 15292 29996 15344 30048
rect 15844 29996 15896 30048
rect 17684 29996 17736 30048
rect 19248 29996 19300 30048
rect 29552 30039 29604 30048
rect 29552 30005 29561 30039
rect 29561 30005 29595 30039
rect 29595 30005 29604 30039
rect 29552 29996 29604 30005
rect 33140 30243 33192 30252
rect 33140 30209 33149 30243
rect 33149 30209 33183 30243
rect 33183 30209 33192 30243
rect 33140 30200 33192 30209
rect 34244 30243 34296 30252
rect 34244 30209 34253 30243
rect 34253 30209 34287 30243
rect 34287 30209 34296 30243
rect 34244 30200 34296 30209
rect 36544 30243 36596 30252
rect 36544 30209 36553 30243
rect 36553 30209 36587 30243
rect 36587 30209 36596 30243
rect 36544 30200 36596 30209
rect 34520 30175 34572 30184
rect 34520 30141 34529 30175
rect 34529 30141 34563 30175
rect 34563 30141 34572 30175
rect 34520 30132 34572 30141
rect 30288 29996 30340 30048
rect 31760 29996 31812 30048
rect 33968 29996 34020 30048
rect 35900 29996 35952 30048
rect 36452 30132 36504 30184
rect 42800 30243 42852 30252
rect 42800 30209 42809 30243
rect 42809 30209 42843 30243
rect 42843 30209 42852 30243
rect 42800 30200 42852 30209
rect 42892 30243 42944 30252
rect 42892 30209 42901 30243
rect 42901 30209 42935 30243
rect 42935 30209 42944 30243
rect 42892 30200 42944 30209
rect 43628 30243 43680 30252
rect 43628 30209 43637 30243
rect 43637 30209 43671 30243
rect 43671 30209 43680 30243
rect 43628 30200 43680 30209
rect 44824 30200 44876 30252
rect 40592 30132 40644 30184
rect 42432 30175 42484 30184
rect 42432 30141 42441 30175
rect 42441 30141 42475 30175
rect 42475 30141 42484 30175
rect 42432 30132 42484 30141
rect 43444 30175 43496 30184
rect 43444 30141 43453 30175
rect 43453 30141 43487 30175
rect 43487 30141 43496 30175
rect 43444 30132 43496 30141
rect 36084 29996 36136 30048
rect 36360 29996 36412 30048
rect 37280 29996 37332 30048
rect 38660 29996 38712 30048
rect 40960 29996 41012 30048
rect 43812 30039 43864 30048
rect 43812 30005 43821 30039
rect 43821 30005 43855 30039
rect 43855 30005 43864 30039
rect 43812 29996 43864 30005
rect 44824 30039 44876 30048
rect 44824 30005 44833 30039
rect 44833 30005 44867 30039
rect 44867 30005 44876 30039
rect 44824 29996 44876 30005
rect 46940 30039 46992 30048
rect 46940 30005 46949 30039
rect 46949 30005 46983 30039
rect 46983 30005 46992 30039
rect 46940 29996 46992 30005
rect 48228 29996 48280 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 11612 29835 11664 29844
rect 11612 29801 11621 29835
rect 11621 29801 11655 29835
rect 11655 29801 11664 29835
rect 11612 29792 11664 29801
rect 15476 29835 15528 29844
rect 15476 29801 15485 29835
rect 15485 29801 15519 29835
rect 15519 29801 15528 29835
rect 15476 29792 15528 29801
rect 15844 29835 15896 29844
rect 15844 29801 15853 29835
rect 15853 29801 15887 29835
rect 15887 29801 15896 29835
rect 15844 29792 15896 29801
rect 16488 29792 16540 29844
rect 17776 29792 17828 29844
rect 18420 29792 18472 29844
rect 18788 29835 18840 29844
rect 18788 29801 18797 29835
rect 18797 29801 18831 29835
rect 18831 29801 18840 29835
rect 18788 29792 18840 29801
rect 20260 29792 20312 29844
rect 22376 29792 22428 29844
rect 31300 29835 31352 29844
rect 31300 29801 31309 29835
rect 31309 29801 31343 29835
rect 31343 29801 31352 29835
rect 31300 29792 31352 29801
rect 34520 29792 34572 29844
rect 37648 29792 37700 29844
rect 9680 29656 9732 29708
rect 10232 29656 10284 29708
rect 11152 29656 11204 29708
rect 14648 29588 14700 29640
rect 15844 29588 15896 29640
rect 17408 29656 17460 29708
rect 9220 29563 9272 29572
rect 9220 29529 9229 29563
rect 9229 29529 9263 29563
rect 9263 29529 9272 29563
rect 9220 29520 9272 29529
rect 11612 29520 11664 29572
rect 16304 29520 16356 29572
rect 2044 29495 2096 29504
rect 2044 29461 2053 29495
rect 2053 29461 2087 29495
rect 2087 29461 2096 29495
rect 2044 29452 2096 29461
rect 10784 29495 10836 29504
rect 10784 29461 10793 29495
rect 10793 29461 10827 29495
rect 10827 29461 10836 29495
rect 10784 29452 10836 29461
rect 14556 29452 14608 29504
rect 17684 29563 17736 29572
rect 17684 29529 17714 29563
rect 17714 29529 17736 29563
rect 18696 29588 18748 29640
rect 35992 29724 36044 29776
rect 19984 29699 20036 29708
rect 19064 29631 19116 29640
rect 19064 29597 19073 29631
rect 19073 29597 19107 29631
rect 19107 29597 19116 29631
rect 19064 29588 19116 29597
rect 19248 29631 19300 29640
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 19984 29665 19993 29699
rect 19993 29665 20027 29699
rect 20027 29665 20036 29699
rect 19984 29656 20036 29665
rect 17684 29520 17736 29529
rect 17960 29563 18012 29572
rect 17960 29529 17969 29563
rect 17969 29529 18003 29563
rect 18003 29529 18012 29563
rect 17960 29520 18012 29529
rect 20076 29631 20128 29640
rect 20076 29597 20085 29631
rect 20085 29597 20119 29631
rect 20119 29597 20128 29631
rect 20076 29588 20128 29597
rect 20812 29656 20864 29708
rect 21456 29656 21508 29708
rect 30196 29656 30248 29708
rect 32128 29656 32180 29708
rect 35900 29656 35952 29708
rect 36360 29656 36412 29708
rect 40960 29656 41012 29708
rect 34244 29588 34296 29640
rect 35992 29631 36044 29640
rect 35992 29597 36001 29631
rect 36001 29597 36035 29631
rect 36035 29597 36044 29631
rect 35992 29588 36044 29597
rect 18052 29452 18104 29504
rect 28356 29520 28408 29572
rect 30104 29520 30156 29572
rect 30288 29520 30340 29572
rect 32956 29520 33008 29572
rect 20444 29452 20496 29504
rect 31576 29452 31628 29504
rect 37280 29452 37332 29504
rect 38660 29520 38712 29572
rect 42616 29520 42668 29572
rect 38476 29452 38528 29504
rect 38844 29495 38896 29504
rect 38844 29461 38853 29495
rect 38853 29461 38887 29495
rect 38887 29461 38896 29495
rect 38844 29452 38896 29461
rect 40224 29452 40276 29504
rect 43812 29588 43864 29640
rect 44364 29520 44416 29572
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 66314 29350 66366 29402
rect 66378 29350 66430 29402
rect 66442 29350 66494 29402
rect 66506 29350 66558 29402
rect 66570 29350 66622 29402
rect 1308 29248 1360 29300
rect 11152 29248 11204 29300
rect 13360 29248 13412 29300
rect 14740 29291 14792 29300
rect 14740 29257 14749 29291
rect 14749 29257 14783 29291
rect 14783 29257 14792 29291
rect 14740 29248 14792 29257
rect 19064 29248 19116 29300
rect 20076 29248 20128 29300
rect 30104 29291 30156 29300
rect 30104 29257 30113 29291
rect 30113 29257 30147 29291
rect 30147 29257 30156 29291
rect 30104 29248 30156 29257
rect 32128 29291 32180 29300
rect 32128 29257 32137 29291
rect 32137 29257 32171 29291
rect 32171 29257 32180 29291
rect 32128 29248 32180 29257
rect 39396 29291 39448 29300
rect 39396 29257 39405 29291
rect 39405 29257 39439 29291
rect 39439 29257 39448 29291
rect 39396 29248 39448 29257
rect 42616 29291 42668 29300
rect 42616 29257 42625 29291
rect 42625 29257 42659 29291
rect 42659 29257 42668 29291
rect 42616 29248 42668 29257
rect 42984 29291 43036 29300
rect 42984 29257 42993 29291
rect 42993 29257 43027 29291
rect 43027 29257 43036 29291
rect 42984 29248 43036 29257
rect 44364 29248 44416 29300
rect 2044 29155 2096 29164
rect 2044 29121 2053 29155
rect 2053 29121 2087 29155
rect 2087 29121 2096 29155
rect 2044 29112 2096 29121
rect 10784 29112 10836 29164
rect 10876 29155 10928 29164
rect 10876 29121 10885 29155
rect 10885 29121 10919 29155
rect 10919 29121 10928 29155
rect 10876 29112 10928 29121
rect 11244 29112 11296 29164
rect 11336 29112 11388 29164
rect 11888 29155 11940 29164
rect 11888 29121 11897 29155
rect 11897 29121 11931 29155
rect 11931 29121 11940 29155
rect 11888 29112 11940 29121
rect 13268 29180 13320 29232
rect 20444 29223 20496 29232
rect 20444 29189 20453 29223
rect 20453 29189 20487 29223
rect 20487 29189 20496 29223
rect 20444 29180 20496 29189
rect 32956 29180 33008 29232
rect 15200 29112 15252 29164
rect 2136 29087 2188 29096
rect 2136 29053 2145 29087
rect 2145 29053 2179 29087
rect 2179 29053 2188 29087
rect 2136 29044 2188 29053
rect 9220 29044 9272 29096
rect 10232 28976 10284 29028
rect 13268 29044 13320 29096
rect 14648 29087 14700 29096
rect 14648 29053 14657 29087
rect 14657 29053 14691 29087
rect 14691 29053 14700 29087
rect 14648 29044 14700 29053
rect 15844 29112 15896 29164
rect 16672 29155 16724 29164
rect 16672 29121 16681 29155
rect 16681 29121 16715 29155
rect 16715 29121 16724 29155
rect 16672 29112 16724 29121
rect 19340 29112 19392 29164
rect 20812 29112 20864 29164
rect 22376 29155 22428 29164
rect 22376 29121 22385 29155
rect 22385 29121 22419 29155
rect 22419 29121 22428 29155
rect 22376 29112 22428 29121
rect 29552 29112 29604 29164
rect 16488 29044 16540 29096
rect 20352 29044 20404 29096
rect 31576 29155 31628 29164
rect 31576 29121 31585 29155
rect 31585 29121 31619 29155
rect 31619 29121 31628 29155
rect 31576 29112 31628 29121
rect 31760 29112 31812 29164
rect 34244 29112 34296 29164
rect 15292 28976 15344 29028
rect 16304 28976 16356 29028
rect 35992 29044 36044 29096
rect 38660 29180 38712 29232
rect 38292 29155 38344 29164
rect 38292 29121 38326 29155
rect 38326 29121 38344 29155
rect 38292 29112 38344 29121
rect 41144 29180 41196 29232
rect 40868 29155 40920 29164
rect 40868 29121 40877 29155
rect 40877 29121 40911 29155
rect 40911 29121 40920 29155
rect 40868 29112 40920 29121
rect 42708 29112 42760 29164
rect 41144 29087 41196 29096
rect 41144 29053 41153 29087
rect 41153 29053 41187 29087
rect 41187 29053 41196 29087
rect 41144 29044 41196 29053
rect 43076 29087 43128 29096
rect 43076 29053 43085 29087
rect 43085 29053 43119 29087
rect 43119 29053 43128 29087
rect 43076 29044 43128 29053
rect 43444 29180 43496 29232
rect 47676 29180 47728 29232
rect 30380 28976 30432 29028
rect 42800 28976 42852 29028
rect 43996 29044 44048 29096
rect 44272 29112 44324 29164
rect 45100 29112 45152 29164
rect 46204 29112 46256 29164
rect 47492 29112 47544 29164
rect 48504 29155 48556 29164
rect 48504 29121 48513 29155
rect 48513 29121 48547 29155
rect 48547 29121 48556 29155
rect 48504 29112 48556 29121
rect 44364 29044 44416 29096
rect 45836 29044 45888 29096
rect 46020 29087 46072 29096
rect 46020 29053 46029 29087
rect 46029 29053 46063 29087
rect 46063 29053 46072 29087
rect 46020 29044 46072 29053
rect 44548 28976 44600 29028
rect 12256 28908 12308 28960
rect 15660 28908 15712 28960
rect 15936 28908 15988 28960
rect 38384 28908 38436 28960
rect 40132 28908 40184 28960
rect 46480 28951 46532 28960
rect 46480 28917 46489 28951
rect 46489 28917 46523 28951
rect 46523 28917 46532 28951
rect 46480 28908 46532 28917
rect 48320 28951 48372 28960
rect 48320 28917 48329 28951
rect 48329 28917 48363 28951
rect 48363 28917 48372 28951
rect 48320 28908 48372 28917
rect 49240 28908 49292 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 10784 28704 10836 28756
rect 940 28636 992 28688
rect 11244 28704 11296 28756
rect 14556 28747 14608 28756
rect 14556 28713 14565 28747
rect 14565 28713 14599 28747
rect 14599 28713 14608 28747
rect 14556 28704 14608 28713
rect 11152 28679 11204 28688
rect 11152 28645 11161 28679
rect 11161 28645 11195 28679
rect 11195 28645 11204 28679
rect 11152 28636 11204 28645
rect 11428 28568 11480 28620
rect 2136 28500 2188 28552
rect 9496 28543 9548 28552
rect 9496 28509 9505 28543
rect 9505 28509 9539 28543
rect 9539 28509 9548 28543
rect 9496 28500 9548 28509
rect 13268 28611 13320 28620
rect 13268 28577 13277 28611
rect 13277 28577 13311 28611
rect 13311 28577 13320 28611
rect 13268 28568 13320 28577
rect 15200 28568 15252 28620
rect 19340 28636 19392 28688
rect 20168 28636 20220 28688
rect 20444 28679 20496 28688
rect 20444 28645 20453 28679
rect 20453 28645 20487 28679
rect 20487 28645 20496 28679
rect 20444 28636 20496 28645
rect 20628 28679 20680 28688
rect 20628 28645 20637 28679
rect 20637 28645 20671 28679
rect 20671 28645 20680 28679
rect 20628 28636 20680 28645
rect 10876 28475 10928 28484
rect 10508 28364 10560 28416
rect 10876 28441 10903 28475
rect 10903 28441 10928 28475
rect 13360 28500 13412 28552
rect 14648 28500 14700 28552
rect 15292 28543 15344 28552
rect 15292 28509 15301 28543
rect 15301 28509 15335 28543
rect 15335 28509 15344 28543
rect 15292 28500 15344 28509
rect 15752 28500 15804 28552
rect 16672 28568 16724 28620
rect 20352 28568 20404 28620
rect 38292 28747 38344 28756
rect 38292 28713 38301 28747
rect 38301 28713 38335 28747
rect 38335 28713 38344 28747
rect 38292 28704 38344 28713
rect 35992 28568 36044 28620
rect 17408 28543 17460 28552
rect 17408 28509 17417 28543
rect 17417 28509 17451 28543
rect 17451 28509 17460 28543
rect 17408 28500 17460 28509
rect 17592 28500 17644 28552
rect 19984 28500 20036 28552
rect 10876 28432 10928 28441
rect 11336 28475 11388 28484
rect 11336 28441 11345 28475
rect 11345 28441 11379 28475
rect 11379 28441 11388 28475
rect 11336 28432 11388 28441
rect 15476 28432 15528 28484
rect 15936 28432 15988 28484
rect 16304 28475 16356 28484
rect 16304 28441 16313 28475
rect 16313 28441 16347 28475
rect 16347 28441 16356 28475
rect 16304 28432 16356 28441
rect 16488 28475 16540 28484
rect 16488 28441 16497 28475
rect 16497 28441 16531 28475
rect 16531 28441 16540 28475
rect 16488 28432 16540 28441
rect 20260 28475 20312 28484
rect 20260 28441 20269 28475
rect 20269 28441 20303 28475
rect 20303 28441 20312 28475
rect 20260 28432 20312 28441
rect 20536 28432 20588 28484
rect 36728 28543 36780 28552
rect 36728 28509 36737 28543
rect 36737 28509 36771 28543
rect 36771 28509 36780 28543
rect 36728 28500 36780 28509
rect 38384 28500 38436 28552
rect 43444 28704 43496 28756
rect 38752 28636 38804 28688
rect 42800 28636 42852 28688
rect 40132 28611 40184 28620
rect 40132 28577 40141 28611
rect 40141 28577 40175 28611
rect 40175 28577 40184 28611
rect 40132 28568 40184 28577
rect 40868 28568 40920 28620
rect 11428 28407 11480 28416
rect 11428 28373 11437 28407
rect 11437 28373 11471 28407
rect 11471 28373 11480 28407
rect 11428 28364 11480 28373
rect 15108 28364 15160 28416
rect 16028 28407 16080 28416
rect 16028 28373 16037 28407
rect 16037 28373 16071 28407
rect 16071 28373 16080 28407
rect 16028 28364 16080 28373
rect 16120 28364 16172 28416
rect 19984 28364 20036 28416
rect 37096 28432 37148 28484
rect 37924 28364 37976 28416
rect 39028 28500 39080 28552
rect 45468 28568 45520 28620
rect 43536 28500 43588 28552
rect 45100 28500 45152 28552
rect 46020 28543 46072 28552
rect 46020 28509 46029 28543
rect 46029 28509 46063 28543
rect 46063 28509 46072 28543
rect 46020 28500 46072 28509
rect 46572 28636 46624 28688
rect 47492 28611 47544 28620
rect 47492 28577 47501 28611
rect 47501 28577 47535 28611
rect 47535 28577 47544 28611
rect 47492 28568 47544 28577
rect 49240 28611 49292 28620
rect 49240 28577 49249 28611
rect 49249 28577 49283 28611
rect 49283 28577 49292 28611
rect 49240 28568 49292 28577
rect 46480 28543 46532 28552
rect 46480 28509 46489 28543
rect 46489 28509 46523 28543
rect 46523 28509 46532 28543
rect 46480 28500 46532 28509
rect 49516 28543 49568 28552
rect 49516 28509 49525 28543
rect 49525 28509 49559 28543
rect 49559 28509 49568 28543
rect 49516 28500 49568 28509
rect 40224 28364 40276 28416
rect 43996 28432 44048 28484
rect 46204 28432 46256 28484
rect 41420 28364 41472 28416
rect 42892 28364 42944 28416
rect 43168 28407 43220 28416
rect 43168 28373 43177 28407
rect 43177 28373 43211 28407
rect 43211 28373 43220 28407
rect 43168 28364 43220 28373
rect 45284 28364 45336 28416
rect 45468 28364 45520 28416
rect 46664 28475 46716 28484
rect 46664 28441 46673 28475
rect 46673 28441 46707 28475
rect 46707 28441 46716 28475
rect 46664 28432 46716 28441
rect 48228 28364 48280 28416
rect 55956 28364 56008 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 66314 28262 66366 28314
rect 66378 28262 66430 28314
rect 66442 28262 66494 28314
rect 66506 28262 66558 28314
rect 66570 28262 66622 28314
rect 9496 28160 9548 28212
rect 10692 28160 10744 28212
rect 14740 28160 14792 28212
rect 17960 28160 18012 28212
rect 20352 28160 20404 28212
rect 20536 28160 20588 28212
rect 10508 28067 10560 28076
rect 10508 28033 10517 28067
rect 10517 28033 10551 28067
rect 10551 28033 10560 28067
rect 10508 28024 10560 28033
rect 10600 28067 10652 28076
rect 10600 28033 10609 28067
rect 10609 28033 10643 28067
rect 10643 28033 10652 28067
rect 10600 28024 10652 28033
rect 10784 28024 10836 28076
rect 10968 28067 11020 28076
rect 10968 28033 10977 28067
rect 10977 28033 11011 28067
rect 11011 28033 11020 28067
rect 10968 28024 11020 28033
rect 13268 28092 13320 28144
rect 15016 28092 15068 28144
rect 16028 28092 16080 28144
rect 18604 28092 18656 28144
rect 19984 28135 20036 28144
rect 19984 28101 19993 28135
rect 19993 28101 20027 28135
rect 20027 28101 20036 28135
rect 19984 28092 20036 28101
rect 20076 28092 20128 28144
rect 42800 28160 42852 28212
rect 45928 28160 45980 28212
rect 15476 28067 15528 28076
rect 15476 28033 15485 28067
rect 15485 28033 15519 28067
rect 15519 28033 15528 28067
rect 15476 28024 15528 28033
rect 15660 28067 15712 28076
rect 15660 28033 15669 28067
rect 15669 28033 15703 28067
rect 15703 28033 15712 28067
rect 15660 28024 15712 28033
rect 15752 28067 15804 28076
rect 15752 28033 15761 28067
rect 15761 28033 15795 28067
rect 15795 28033 15804 28067
rect 15752 28024 15804 28033
rect 16120 28024 16172 28076
rect 20168 28067 20220 28076
rect 20168 28033 20177 28067
rect 20177 28033 20211 28067
rect 20211 28033 20220 28067
rect 20168 28024 20220 28033
rect 37096 28092 37148 28144
rect 42892 28092 42944 28144
rect 45468 28135 45520 28144
rect 10232 27956 10284 28008
rect 13360 27999 13412 28008
rect 13360 27965 13369 27999
rect 13369 27965 13403 27999
rect 13403 27965 13412 27999
rect 13360 27956 13412 27965
rect 14740 27956 14792 28008
rect 32036 27956 32088 28008
rect 33232 27999 33284 28008
rect 33232 27965 33241 27999
rect 33241 27965 33275 27999
rect 33275 27965 33284 27999
rect 33232 27956 33284 27965
rect 40868 28024 40920 28076
rect 42800 28024 42852 28076
rect 35348 27956 35400 28008
rect 41236 27999 41288 28008
rect 41236 27965 41245 27999
rect 41245 27965 41279 27999
rect 41279 27965 41288 27999
rect 41236 27956 41288 27965
rect 42984 27956 43036 28008
rect 45468 28101 45477 28135
rect 45477 28101 45511 28135
rect 45511 28101 45520 28135
rect 47492 28160 47544 28212
rect 48504 28160 48556 28212
rect 45468 28092 45520 28101
rect 46664 28092 46716 28144
rect 43536 28024 43588 28076
rect 43720 28024 43772 28076
rect 44180 28067 44232 28076
rect 44180 28033 44190 28067
rect 44190 28033 44224 28067
rect 44224 28033 44232 28067
rect 44180 28024 44232 28033
rect 44732 28024 44784 28076
rect 45100 28024 45152 28076
rect 46572 28024 46624 28076
rect 48320 28024 48372 28076
rect 940 27888 992 27940
rect 14648 27820 14700 27872
rect 16120 27863 16172 27872
rect 16120 27829 16129 27863
rect 16129 27829 16163 27863
rect 16163 27829 16172 27863
rect 16120 27820 16172 27829
rect 18604 27863 18656 27872
rect 18604 27829 18613 27863
rect 18613 27829 18647 27863
rect 18647 27829 18656 27863
rect 18604 27820 18656 27829
rect 19432 27820 19484 27872
rect 34520 27820 34572 27872
rect 36544 27820 36596 27872
rect 42984 27820 43036 27872
rect 46112 27956 46164 28008
rect 44732 27888 44784 27940
rect 43628 27820 43680 27872
rect 45836 27820 45888 27872
rect 46020 27863 46072 27872
rect 46020 27829 46029 27863
rect 46029 27829 46063 27863
rect 46063 27829 46072 27863
rect 46020 27820 46072 27829
rect 46112 27863 46164 27872
rect 46112 27829 46121 27863
rect 46121 27829 46155 27863
rect 46155 27829 46164 27863
rect 46112 27820 46164 27829
rect 47676 27820 47728 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 10600 27616 10652 27668
rect 16120 27659 16172 27668
rect 16120 27625 16150 27659
rect 16150 27625 16172 27659
rect 16120 27616 16172 27625
rect 17592 27659 17644 27668
rect 17592 27625 17601 27659
rect 17601 27625 17635 27659
rect 17635 27625 17644 27659
rect 17592 27616 17644 27625
rect 33232 27616 33284 27668
rect 35348 27616 35400 27668
rect 36728 27616 36780 27668
rect 42708 27616 42760 27668
rect 13360 27548 13412 27600
rect 34428 27548 34480 27600
rect 12440 27523 12492 27532
rect 12440 27489 12449 27523
rect 12449 27489 12483 27523
rect 12483 27489 12492 27523
rect 12440 27480 12492 27489
rect 14740 27480 14792 27532
rect 20168 27480 20220 27532
rect 31668 27480 31720 27532
rect 10968 27455 11020 27464
rect 10968 27421 10977 27455
rect 10977 27421 11011 27455
rect 11011 27421 11020 27455
rect 10968 27412 11020 27421
rect 11336 27412 11388 27464
rect 14648 27455 14700 27464
rect 14648 27421 14657 27455
rect 14657 27421 14691 27455
rect 14691 27421 14700 27455
rect 14648 27412 14700 27421
rect 19432 27455 19484 27464
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 15016 27344 15068 27396
rect 23572 27412 23624 27464
rect 34060 27455 34112 27464
rect 34060 27421 34069 27455
rect 34069 27421 34103 27455
rect 34103 27421 34112 27455
rect 34060 27412 34112 27421
rect 34152 27455 34204 27464
rect 34152 27421 34161 27455
rect 34161 27421 34195 27455
rect 34195 27421 34204 27455
rect 34152 27412 34204 27421
rect 34520 27412 34572 27464
rect 940 27276 992 27328
rect 20628 27344 20680 27396
rect 17960 27276 18012 27328
rect 18512 27276 18564 27328
rect 20352 27276 20404 27328
rect 21916 27344 21968 27396
rect 32588 27344 32640 27396
rect 35440 27455 35492 27464
rect 35440 27421 35449 27455
rect 35449 27421 35483 27455
rect 35483 27421 35492 27455
rect 35440 27412 35492 27421
rect 36544 27412 36596 27464
rect 36912 27455 36964 27464
rect 36912 27421 36921 27455
rect 36921 27421 36955 27455
rect 36955 27421 36964 27455
rect 36912 27412 36964 27421
rect 22836 27276 22888 27328
rect 36360 27276 36412 27328
rect 37832 27523 37884 27532
rect 37832 27489 37841 27523
rect 37841 27489 37875 27523
rect 37875 27489 37884 27523
rect 37832 27480 37884 27489
rect 38752 27480 38804 27532
rect 42892 27548 42944 27600
rect 43536 27616 43588 27668
rect 37924 27412 37976 27464
rect 38108 27412 38160 27464
rect 44180 27480 44232 27532
rect 39212 27344 39264 27396
rect 41236 27344 41288 27396
rect 42984 27412 43036 27464
rect 43352 27455 43404 27464
rect 43352 27421 43361 27455
rect 43361 27421 43395 27455
rect 43395 27421 43404 27455
rect 43352 27412 43404 27421
rect 43628 27455 43680 27464
rect 43628 27421 43637 27455
rect 43637 27421 43671 27455
rect 43671 27421 43680 27455
rect 43628 27412 43680 27421
rect 43720 27455 43772 27464
rect 43720 27421 43730 27455
rect 43730 27421 43764 27455
rect 43764 27421 43772 27455
rect 43720 27412 43772 27421
rect 45836 27455 45888 27464
rect 45836 27421 45845 27455
rect 45845 27421 45879 27455
rect 45879 27421 45888 27455
rect 45836 27412 45888 27421
rect 38660 27276 38712 27328
rect 43260 27319 43312 27328
rect 43260 27285 43269 27319
rect 43269 27285 43303 27319
rect 43303 27285 43312 27319
rect 43260 27276 43312 27285
rect 45928 27319 45980 27328
rect 45928 27285 45937 27319
rect 45937 27285 45971 27319
rect 45971 27285 45980 27319
rect 45928 27276 45980 27285
rect 49332 27276 49384 27328
rect 51264 27276 51316 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 66314 27174 66366 27226
rect 66378 27174 66430 27226
rect 66442 27174 66494 27226
rect 66506 27174 66558 27226
rect 66570 27174 66622 27226
rect 10784 27072 10836 27124
rect 12072 27072 12124 27124
rect 10048 27004 10100 27056
rect 10600 26936 10652 26988
rect 11336 26936 11388 26988
rect 12072 26936 12124 26988
rect 12440 26979 12492 26988
rect 12440 26945 12449 26979
rect 12449 26945 12483 26979
rect 12483 26945 12492 26979
rect 12440 26936 12492 26945
rect 18144 27072 18196 27124
rect 18604 27072 18656 27124
rect 20168 27072 20220 27124
rect 21916 27072 21968 27124
rect 31392 27072 31444 27124
rect 18512 27047 18564 27056
rect 18512 27013 18521 27047
rect 18521 27013 18555 27047
rect 18555 27013 18564 27047
rect 18512 27004 18564 27013
rect 35440 27072 35492 27124
rect 34520 27004 34572 27056
rect 12992 26936 13044 26988
rect 13360 26936 13412 26988
rect 14740 26979 14792 26988
rect 14740 26945 14749 26979
rect 14749 26945 14783 26979
rect 14783 26945 14792 26979
rect 14740 26936 14792 26945
rect 20444 26979 20496 26988
rect 20444 26945 20453 26979
rect 20453 26945 20487 26979
rect 20487 26945 20496 26979
rect 20444 26936 20496 26945
rect 20628 26979 20680 26988
rect 20628 26945 20637 26979
rect 20637 26945 20671 26979
rect 20671 26945 20680 26979
rect 20628 26936 20680 26945
rect 2044 26911 2096 26920
rect 2044 26877 2053 26911
rect 2053 26877 2087 26911
rect 2087 26877 2096 26911
rect 2044 26868 2096 26877
rect 10140 26775 10192 26784
rect 10140 26741 10149 26775
rect 10149 26741 10183 26775
rect 10183 26741 10192 26775
rect 10140 26732 10192 26741
rect 12164 26800 12216 26852
rect 18236 26911 18288 26920
rect 18236 26877 18245 26911
rect 18245 26877 18279 26911
rect 18279 26877 18288 26911
rect 18236 26868 18288 26877
rect 32036 26868 32088 26920
rect 32496 26911 32548 26920
rect 32496 26877 32505 26911
rect 32505 26877 32539 26911
rect 32539 26877 32548 26911
rect 32496 26868 32548 26877
rect 12532 26800 12584 26852
rect 11980 26732 12032 26784
rect 12992 26775 13044 26784
rect 12992 26741 13001 26775
rect 13001 26741 13035 26775
rect 13035 26741 13044 26775
rect 12992 26732 13044 26741
rect 14648 26732 14700 26784
rect 18144 26775 18196 26784
rect 18144 26741 18153 26775
rect 18153 26741 18187 26775
rect 18187 26741 18196 26775
rect 18144 26732 18196 26741
rect 33968 26732 34020 26784
rect 34612 26732 34664 26784
rect 35532 26979 35584 26988
rect 35532 26945 35541 26979
rect 35541 26945 35575 26979
rect 35575 26945 35584 26979
rect 35532 26936 35584 26945
rect 35624 26979 35676 26988
rect 35624 26945 35633 26979
rect 35633 26945 35667 26979
rect 35667 26945 35676 26979
rect 35624 26936 35676 26945
rect 36728 27072 36780 27124
rect 36912 27115 36964 27124
rect 36912 27081 36921 27115
rect 36921 27081 36955 27115
rect 36955 27081 36964 27115
rect 36912 27072 36964 27081
rect 38108 27115 38160 27124
rect 38108 27081 38117 27115
rect 38117 27081 38151 27115
rect 38151 27081 38160 27115
rect 38108 27072 38160 27081
rect 37004 27004 37056 27056
rect 39212 27004 39264 27056
rect 36544 26868 36596 26920
rect 36728 26979 36780 26988
rect 36728 26945 36737 26979
rect 36737 26945 36771 26979
rect 36771 26945 36780 26979
rect 36728 26936 36780 26945
rect 37280 26936 37332 26988
rect 37372 26936 37424 26988
rect 38384 26979 38436 26988
rect 38384 26945 38393 26979
rect 38393 26945 38427 26979
rect 38427 26945 38436 26979
rect 38384 26936 38436 26945
rect 38660 26979 38712 26988
rect 38660 26945 38669 26979
rect 38669 26945 38703 26979
rect 38703 26945 38712 26979
rect 38660 26936 38712 26945
rect 38752 26936 38804 26988
rect 42800 26936 42852 26988
rect 43720 27072 43772 27124
rect 46020 27115 46072 27124
rect 46020 27081 46029 27115
rect 46029 27081 46063 27115
rect 46063 27081 46072 27115
rect 46020 27072 46072 27081
rect 48412 27072 48464 27124
rect 43536 26936 43588 26988
rect 40408 26868 40460 26920
rect 41236 26868 41288 26920
rect 43260 26868 43312 26920
rect 43352 26911 43404 26920
rect 43352 26877 43361 26911
rect 43361 26877 43395 26911
rect 43395 26877 43404 26911
rect 53932 27004 53984 27056
rect 43352 26868 43404 26877
rect 44272 26868 44324 26920
rect 37188 26800 37240 26852
rect 43628 26800 43680 26852
rect 44180 26843 44232 26852
rect 44180 26809 44189 26843
rect 44189 26809 44223 26843
rect 44223 26809 44232 26843
rect 44180 26800 44232 26809
rect 38108 26732 38160 26784
rect 38936 26732 38988 26784
rect 42708 26732 42760 26784
rect 43720 26732 43772 26784
rect 44824 26911 44876 26920
rect 44824 26877 44833 26911
rect 44833 26877 44867 26911
rect 44867 26877 44876 26911
rect 44824 26868 44876 26877
rect 45284 26936 45336 26988
rect 48504 26911 48556 26920
rect 48504 26877 48513 26911
rect 48513 26877 48547 26911
rect 48547 26877 48556 26911
rect 48504 26868 48556 26877
rect 49148 26868 49200 26920
rect 45928 26800 45980 26852
rect 49976 26732 50028 26784
rect 51172 26868 51224 26920
rect 51264 26868 51316 26920
rect 52368 26868 52420 26920
rect 54208 26911 54260 26920
rect 54208 26877 54217 26911
rect 54217 26877 54251 26911
rect 54251 26877 54260 26911
rect 54208 26868 54260 26877
rect 54484 26911 54536 26920
rect 54484 26877 54493 26911
rect 54493 26877 54527 26911
rect 54527 26877 54536 26911
rect 54484 26868 54536 26877
rect 51080 26732 51132 26784
rect 52092 26775 52144 26784
rect 52092 26741 52101 26775
rect 52101 26741 52135 26775
rect 52135 26741 52144 26775
rect 52092 26732 52144 26741
rect 52736 26775 52788 26784
rect 52736 26741 52745 26775
rect 52745 26741 52779 26775
rect 52779 26741 52788 26775
rect 52736 26732 52788 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 1308 26528 1360 26580
rect 10968 26528 11020 26580
rect 11980 26571 12032 26580
rect 11980 26537 11989 26571
rect 11989 26537 12023 26571
rect 12023 26537 12032 26571
rect 11980 26528 12032 26537
rect 12440 26528 12492 26580
rect 20352 26571 20404 26580
rect 20352 26537 20361 26571
rect 20361 26537 20395 26571
rect 20395 26537 20404 26571
rect 20352 26528 20404 26537
rect 31116 26528 31168 26580
rect 31668 26528 31720 26580
rect 32496 26528 32548 26580
rect 34152 26528 34204 26580
rect 40408 26571 40460 26580
rect 40408 26537 40417 26571
rect 40417 26537 40451 26571
rect 40451 26537 40460 26571
rect 40408 26528 40460 26537
rect 41144 26528 41196 26580
rect 42800 26528 42852 26580
rect 49148 26571 49200 26580
rect 49148 26537 49157 26571
rect 49157 26537 49191 26571
rect 49191 26537 49200 26571
rect 49148 26528 49200 26537
rect 51540 26528 51592 26580
rect 54208 26528 54260 26580
rect 10232 26392 10284 26444
rect 10692 26392 10744 26444
rect 13360 26460 13412 26512
rect 2044 26367 2096 26376
rect 2044 26333 2053 26367
rect 2053 26333 2087 26367
rect 2087 26333 2096 26367
rect 2044 26324 2096 26333
rect 10140 26256 10192 26308
rect 10324 26256 10376 26308
rect 10692 26256 10744 26308
rect 12532 26392 12584 26444
rect 12900 26392 12952 26444
rect 20628 26392 20680 26444
rect 12072 26324 12124 26376
rect 12440 26367 12492 26376
rect 12440 26333 12449 26367
rect 12449 26333 12483 26367
rect 12483 26333 12492 26367
rect 12440 26324 12492 26333
rect 12992 26324 13044 26376
rect 20168 26324 20220 26376
rect 12164 26299 12216 26308
rect 12164 26265 12173 26299
rect 12173 26265 12207 26299
rect 12207 26265 12216 26299
rect 12164 26256 12216 26265
rect 20720 26256 20772 26308
rect 30380 26324 30432 26376
rect 30840 26367 30892 26376
rect 30840 26333 30849 26367
rect 30849 26333 30883 26367
rect 30883 26333 30892 26367
rect 30840 26324 30892 26333
rect 31576 26324 31628 26376
rect 32128 26367 32180 26376
rect 32128 26333 32159 26367
rect 32159 26333 32180 26367
rect 32128 26324 32180 26333
rect 32404 26367 32456 26376
rect 32404 26333 32413 26367
rect 32413 26333 32447 26367
rect 32447 26333 32456 26367
rect 32404 26324 32456 26333
rect 32588 26324 32640 26376
rect 34612 26324 34664 26376
rect 44088 26460 44140 26512
rect 46020 26460 46072 26512
rect 36544 26324 36596 26376
rect 41236 26324 41288 26376
rect 43628 26324 43680 26376
rect 44732 26324 44784 26376
rect 45008 26324 45060 26376
rect 34520 26256 34572 26308
rect 35072 26299 35124 26308
rect 35072 26265 35081 26299
rect 35081 26265 35115 26299
rect 35115 26265 35124 26299
rect 35072 26256 35124 26265
rect 35624 26256 35676 26308
rect 44456 26299 44508 26308
rect 44456 26265 44465 26299
rect 44465 26265 44499 26299
rect 44499 26265 44508 26299
rect 44456 26256 44508 26265
rect 45468 26324 45520 26376
rect 45836 26392 45888 26444
rect 48504 26392 48556 26444
rect 49516 26460 49568 26512
rect 51080 26460 51132 26512
rect 49976 26392 50028 26444
rect 46112 26299 46164 26308
rect 46112 26265 46129 26299
rect 46129 26265 46164 26299
rect 46112 26256 46164 26265
rect 19432 26188 19484 26240
rect 21364 26231 21416 26240
rect 21364 26197 21373 26231
rect 21373 26197 21407 26231
rect 21407 26197 21416 26231
rect 21364 26188 21416 26197
rect 30564 26231 30616 26240
rect 30564 26197 30573 26231
rect 30573 26197 30607 26231
rect 30607 26197 30616 26231
rect 30564 26188 30616 26197
rect 40868 26231 40920 26240
rect 40868 26197 40877 26231
rect 40877 26197 40911 26231
rect 40911 26197 40920 26231
rect 40868 26188 40920 26197
rect 44824 26188 44876 26240
rect 45284 26188 45336 26240
rect 46480 26367 46532 26376
rect 46480 26333 46489 26367
rect 46489 26333 46523 26367
rect 46523 26333 46532 26367
rect 46480 26324 46532 26333
rect 49332 26367 49384 26376
rect 49332 26333 49341 26367
rect 49341 26333 49375 26367
rect 49375 26333 49384 26367
rect 49332 26324 49384 26333
rect 52276 26392 52328 26444
rect 54484 26460 54536 26512
rect 52460 26392 52512 26444
rect 46756 26299 46808 26308
rect 46756 26265 46765 26299
rect 46765 26265 46799 26299
rect 46799 26265 46808 26299
rect 46756 26256 46808 26265
rect 48412 26256 48464 26308
rect 48504 26299 48556 26308
rect 48504 26265 48513 26299
rect 48513 26265 48547 26299
rect 48547 26265 48556 26299
rect 48504 26256 48556 26265
rect 51356 26324 51408 26376
rect 52736 26367 52788 26376
rect 49884 26256 49936 26308
rect 50804 26256 50856 26308
rect 52736 26333 52745 26367
rect 52745 26333 52779 26367
rect 52779 26333 52788 26367
rect 52736 26324 52788 26333
rect 53748 26367 53800 26376
rect 53748 26333 53757 26367
rect 53757 26333 53791 26367
rect 53791 26333 53800 26367
rect 53748 26324 53800 26333
rect 51816 26256 51868 26308
rect 52460 26256 52512 26308
rect 53012 26256 53064 26308
rect 51448 26231 51500 26240
rect 51448 26197 51457 26231
rect 51457 26197 51491 26231
rect 51491 26197 51500 26231
rect 51448 26188 51500 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 66314 26086 66366 26138
rect 66378 26086 66430 26138
rect 66442 26086 66494 26138
rect 66506 26086 66558 26138
rect 66570 26086 66622 26138
rect 940 25984 992 26036
rect 10048 25984 10100 26036
rect 12992 25984 13044 26036
rect 15476 25984 15528 26036
rect 16948 25984 17000 26036
rect 17960 25984 18012 26036
rect 29184 25984 29236 26036
rect 15108 25959 15160 25968
rect 15108 25925 15117 25959
rect 15117 25925 15151 25959
rect 15151 25925 15160 25959
rect 15108 25916 15160 25925
rect 19432 25916 19484 25968
rect 17592 25848 17644 25900
rect 17960 25848 18012 25900
rect 19524 25848 19576 25900
rect 17316 25780 17368 25832
rect 20628 25848 20680 25900
rect 21364 25916 21416 25968
rect 22836 25916 22888 25968
rect 31392 25984 31444 26036
rect 32404 26027 32456 26036
rect 32404 25993 32413 26027
rect 32413 25993 32447 26027
rect 32447 25993 32456 26027
rect 32404 25984 32456 25993
rect 37280 25984 37332 26036
rect 37740 25984 37792 26036
rect 38384 25984 38436 26036
rect 40868 26027 40920 26036
rect 40868 25993 40877 26027
rect 40877 25993 40911 26027
rect 40911 25993 40920 26027
rect 40868 25984 40920 25993
rect 43076 25984 43128 26036
rect 46480 25984 46532 26036
rect 46756 25984 46808 26036
rect 48504 25984 48556 26036
rect 49884 26027 49936 26036
rect 49884 25993 49893 26027
rect 49893 25993 49927 26027
rect 49927 25993 49936 26027
rect 49884 25984 49936 25993
rect 51080 26027 51132 26036
rect 51080 25993 51089 26027
rect 51089 25993 51123 26027
rect 51123 25993 51132 26027
rect 51080 25984 51132 25993
rect 51356 25984 51408 26036
rect 53748 25984 53800 26036
rect 20076 25780 20128 25832
rect 23572 25823 23624 25832
rect 23572 25789 23581 25823
rect 23581 25789 23615 25823
rect 23615 25789 23624 25823
rect 23572 25780 23624 25789
rect 20720 25712 20772 25764
rect 31576 25916 31628 25968
rect 32588 25891 32640 25900
rect 32588 25857 32597 25891
rect 32597 25857 32631 25891
rect 32631 25857 32640 25891
rect 32588 25848 32640 25857
rect 34796 25916 34848 25968
rect 35072 25916 35124 25968
rect 28448 25780 28500 25832
rect 30564 25780 30616 25832
rect 31392 25780 31444 25832
rect 29184 25712 29236 25764
rect 14556 25644 14608 25696
rect 17684 25687 17736 25696
rect 17684 25653 17693 25687
rect 17693 25653 17727 25687
rect 17727 25653 17736 25687
rect 17684 25644 17736 25653
rect 19064 25644 19116 25696
rect 34060 25848 34112 25900
rect 36636 25848 36688 25900
rect 37372 25848 37424 25900
rect 34244 25823 34296 25832
rect 34244 25789 34253 25823
rect 34253 25789 34287 25823
rect 34287 25789 34296 25823
rect 34244 25780 34296 25789
rect 37740 25891 37792 25900
rect 37740 25857 37749 25891
rect 37749 25857 37783 25891
rect 37783 25857 37792 25891
rect 37740 25848 37792 25857
rect 38108 25848 38160 25900
rect 43168 25916 43220 25968
rect 37648 25712 37700 25764
rect 37924 25780 37976 25832
rect 42800 25848 42852 25900
rect 44548 25891 44600 25900
rect 44548 25857 44557 25891
rect 44557 25857 44591 25891
rect 44591 25857 44600 25891
rect 44548 25848 44600 25857
rect 45008 25916 45060 25968
rect 45468 25916 45520 25968
rect 44824 25891 44876 25900
rect 44824 25857 44833 25891
rect 44833 25857 44867 25891
rect 44867 25857 44876 25891
rect 44824 25848 44876 25857
rect 45284 25848 45336 25900
rect 49148 25848 49200 25900
rect 49424 25848 49476 25900
rect 52552 25916 52604 25968
rect 41236 25780 41288 25832
rect 38752 25712 38804 25764
rect 47676 25823 47728 25832
rect 47676 25789 47685 25823
rect 47685 25789 47719 25823
rect 47719 25789 47728 25823
rect 47676 25780 47728 25789
rect 47952 25780 48004 25832
rect 51172 25848 51224 25900
rect 51448 25848 51500 25900
rect 51540 25823 51592 25832
rect 51540 25789 51549 25823
rect 51549 25789 51583 25823
rect 51583 25789 51592 25823
rect 51540 25780 51592 25789
rect 44180 25712 44232 25764
rect 44732 25712 44784 25764
rect 46756 25712 46808 25764
rect 51172 25712 51224 25764
rect 52092 25848 52144 25900
rect 53012 25780 53064 25832
rect 34704 25644 34756 25696
rect 37280 25687 37332 25696
rect 37280 25653 37289 25687
rect 37289 25653 37323 25687
rect 37323 25653 37332 25687
rect 37280 25644 37332 25653
rect 44364 25687 44416 25696
rect 44364 25653 44373 25687
rect 44373 25653 44407 25687
rect 44407 25653 44416 25687
rect 44364 25644 44416 25653
rect 50528 25644 50580 25696
rect 51816 25687 51868 25696
rect 51816 25653 51825 25687
rect 51825 25653 51859 25687
rect 51859 25653 51868 25687
rect 51816 25644 51868 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 13820 25440 13872 25492
rect 12440 25304 12492 25356
rect 12900 25279 12952 25288
rect 12900 25245 12909 25279
rect 12909 25245 12943 25279
rect 12943 25245 12952 25279
rect 12900 25236 12952 25245
rect 13452 25236 13504 25288
rect 13728 25236 13780 25288
rect 14556 25483 14608 25492
rect 14556 25449 14565 25483
rect 14565 25449 14599 25483
rect 14599 25449 14608 25483
rect 14556 25440 14608 25449
rect 20628 25440 20680 25492
rect 17684 25372 17736 25424
rect 16580 25304 16632 25356
rect 18236 25304 18288 25356
rect 23572 25304 23624 25356
rect 14372 25279 14424 25288
rect 14372 25245 14381 25279
rect 14381 25245 14415 25279
rect 14415 25245 14424 25279
rect 14372 25236 14424 25245
rect 14464 25236 14516 25288
rect 15016 25236 15068 25288
rect 16948 25236 17000 25288
rect 13176 25168 13228 25220
rect 17684 25279 17736 25288
rect 17684 25245 17693 25279
rect 17693 25245 17727 25279
rect 17727 25245 17736 25279
rect 17684 25236 17736 25245
rect 17960 25279 18012 25288
rect 17960 25245 17969 25279
rect 17969 25245 18003 25279
rect 18003 25245 18012 25279
rect 17960 25236 18012 25245
rect 18328 25236 18380 25288
rect 19064 25279 19116 25288
rect 19064 25245 19073 25279
rect 19073 25245 19107 25279
rect 19107 25245 19116 25279
rect 19064 25236 19116 25245
rect 940 25100 992 25152
rect 14740 25143 14792 25152
rect 14740 25109 14749 25143
rect 14749 25109 14783 25143
rect 14783 25109 14792 25143
rect 14740 25100 14792 25109
rect 17868 25168 17920 25220
rect 27712 25440 27764 25492
rect 29368 25440 29420 25492
rect 30840 25440 30892 25492
rect 42432 25440 42484 25492
rect 51540 25440 51592 25492
rect 51908 25483 51960 25492
rect 51908 25449 51917 25483
rect 51917 25449 51951 25483
rect 51951 25449 51960 25483
rect 51908 25440 51960 25449
rect 53656 25483 53708 25492
rect 53656 25449 53665 25483
rect 53665 25449 53699 25483
rect 53699 25449 53708 25483
rect 53656 25440 53708 25449
rect 31300 25304 31352 25356
rect 32588 25304 32640 25356
rect 34428 25347 34480 25356
rect 34428 25313 34437 25347
rect 34437 25313 34471 25347
rect 34471 25313 34480 25347
rect 34428 25304 34480 25313
rect 34796 25304 34848 25356
rect 31392 25279 31444 25288
rect 31392 25245 31401 25279
rect 31401 25245 31435 25279
rect 31435 25245 31444 25279
rect 31392 25236 31444 25245
rect 32128 25236 32180 25288
rect 33968 25236 34020 25288
rect 34060 25236 34112 25288
rect 16856 25100 16908 25152
rect 17316 25143 17368 25152
rect 17316 25109 17325 25143
rect 17325 25109 17359 25143
rect 17359 25109 17368 25143
rect 17316 25100 17368 25109
rect 17408 25143 17460 25152
rect 17408 25109 17417 25143
rect 17417 25109 17451 25143
rect 17451 25109 17460 25143
rect 17408 25100 17460 25109
rect 17776 25143 17828 25152
rect 17776 25109 17785 25143
rect 17785 25109 17819 25143
rect 17819 25109 17828 25143
rect 17776 25100 17828 25109
rect 18144 25143 18196 25152
rect 18144 25109 18153 25143
rect 18153 25109 18187 25143
rect 18187 25109 18196 25143
rect 18144 25100 18196 25109
rect 18328 25143 18380 25152
rect 18328 25109 18337 25143
rect 18337 25109 18371 25143
rect 18371 25109 18380 25143
rect 18328 25100 18380 25109
rect 18512 25143 18564 25152
rect 18512 25109 18521 25143
rect 18521 25109 18555 25143
rect 18555 25109 18564 25143
rect 18512 25100 18564 25109
rect 18604 25100 18656 25152
rect 28448 25168 28500 25220
rect 30932 25168 30984 25220
rect 34520 25279 34572 25288
rect 34520 25245 34529 25279
rect 34529 25245 34563 25279
rect 34563 25245 34572 25279
rect 34520 25236 34572 25245
rect 34888 25279 34940 25288
rect 34888 25245 34897 25279
rect 34897 25245 34931 25279
rect 34931 25245 34940 25279
rect 34888 25236 34940 25245
rect 37832 25347 37884 25356
rect 37832 25313 37841 25347
rect 37841 25313 37875 25347
rect 37875 25313 37884 25347
rect 37832 25304 37884 25313
rect 35440 25236 35492 25288
rect 33784 25100 33836 25152
rect 34796 25168 34848 25220
rect 34888 25100 34940 25152
rect 36084 25279 36136 25288
rect 36084 25245 36093 25279
rect 36093 25245 36127 25279
rect 36127 25245 36136 25279
rect 36084 25236 36136 25245
rect 38200 25279 38252 25288
rect 38200 25245 38209 25279
rect 38209 25245 38243 25279
rect 38243 25245 38252 25279
rect 38200 25236 38252 25245
rect 42524 25372 42576 25424
rect 42800 25372 42852 25424
rect 40868 25304 40920 25356
rect 41420 25279 41472 25288
rect 41420 25245 41429 25279
rect 41429 25245 41463 25279
rect 41463 25245 41472 25279
rect 41420 25236 41472 25245
rect 37096 25168 37148 25220
rect 39212 25168 39264 25220
rect 42156 25236 42208 25288
rect 42616 25236 42668 25288
rect 41696 25211 41748 25220
rect 41696 25177 41705 25211
rect 41705 25177 41739 25211
rect 41739 25177 41748 25211
rect 41696 25168 41748 25177
rect 37556 25100 37608 25152
rect 39764 25100 39816 25152
rect 41236 25100 41288 25152
rect 43168 25304 43220 25356
rect 52368 25372 52420 25424
rect 54484 25372 54536 25424
rect 46572 25236 46624 25288
rect 51264 25236 51316 25288
rect 43352 25168 43404 25220
rect 51724 25279 51776 25288
rect 51724 25245 51733 25279
rect 51733 25245 51767 25279
rect 51767 25245 51776 25279
rect 51724 25236 51776 25245
rect 52000 25279 52052 25288
rect 52000 25245 52009 25279
rect 52009 25245 52043 25279
rect 52043 25245 52052 25279
rect 52000 25236 52052 25245
rect 53380 25279 53432 25288
rect 53380 25245 53389 25279
rect 53389 25245 53423 25279
rect 53423 25245 53432 25279
rect 53380 25236 53432 25245
rect 53472 25279 53524 25288
rect 53472 25245 53481 25279
rect 53481 25245 53515 25279
rect 53515 25245 53524 25279
rect 53472 25236 53524 25245
rect 53564 25236 53616 25288
rect 52276 25168 52328 25220
rect 55588 25211 55640 25220
rect 55588 25177 55597 25211
rect 55597 25177 55631 25211
rect 55631 25177 55640 25211
rect 55588 25168 55640 25177
rect 43720 25100 43772 25152
rect 51080 25100 51132 25152
rect 53196 25143 53248 25152
rect 53196 25109 53205 25143
rect 53205 25109 53239 25143
rect 53239 25109 53248 25143
rect 53196 25100 53248 25109
rect 53932 25100 53984 25152
rect 54484 25100 54536 25152
rect 55772 25100 55824 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 66314 24998 66366 25050
rect 66378 24998 66430 25050
rect 66442 24998 66494 25050
rect 66506 24998 66558 25050
rect 66570 24998 66622 25050
rect 12900 24896 12952 24948
rect 13728 24896 13780 24948
rect 14372 24896 14424 24948
rect 13820 24828 13872 24880
rect 17408 24896 17460 24948
rect 17868 24896 17920 24948
rect 18052 24896 18104 24948
rect 18604 24896 18656 24948
rect 20076 24939 20128 24948
rect 20076 24905 20103 24939
rect 20103 24905 20128 24939
rect 20076 24896 20128 24905
rect 7748 24735 7800 24744
rect 7748 24701 7757 24735
rect 7757 24701 7791 24735
rect 7791 24701 7800 24735
rect 7748 24692 7800 24701
rect 9036 24692 9088 24744
rect 10876 24760 10928 24812
rect 10416 24624 10468 24676
rect 11060 24735 11112 24744
rect 11060 24701 11069 24735
rect 11069 24701 11103 24735
rect 11103 24701 11112 24735
rect 11060 24692 11112 24701
rect 11152 24692 11204 24744
rect 12532 24803 12584 24812
rect 12532 24769 12541 24803
rect 12541 24769 12575 24803
rect 12575 24769 12584 24803
rect 12532 24760 12584 24769
rect 13728 24760 13780 24812
rect 13452 24735 13504 24744
rect 13452 24701 13461 24735
rect 13461 24701 13495 24735
rect 13495 24701 13504 24735
rect 13452 24692 13504 24701
rect 14280 24803 14332 24812
rect 14280 24769 14289 24803
rect 14289 24769 14323 24803
rect 14323 24769 14332 24803
rect 14280 24760 14332 24769
rect 15108 24760 15160 24812
rect 20628 24828 20680 24880
rect 30840 24896 30892 24948
rect 34520 24896 34572 24948
rect 35348 24896 35400 24948
rect 36084 24896 36136 24948
rect 29184 24828 29236 24880
rect 16856 24760 16908 24812
rect 17316 24760 17368 24812
rect 17776 24760 17828 24812
rect 18512 24760 18564 24812
rect 28448 24803 28500 24812
rect 28448 24769 28457 24803
rect 28457 24769 28491 24803
rect 28491 24769 28500 24803
rect 28448 24760 28500 24769
rect 30472 24760 30524 24812
rect 30656 24803 30708 24812
rect 30656 24769 30665 24803
rect 30665 24769 30699 24803
rect 30699 24769 30708 24803
rect 30656 24760 30708 24769
rect 30932 24803 30984 24812
rect 30932 24769 30941 24803
rect 30941 24769 30975 24803
rect 30975 24769 30984 24803
rect 30932 24760 30984 24769
rect 33784 24803 33836 24812
rect 33784 24769 33793 24803
rect 33793 24769 33827 24803
rect 33827 24769 33836 24803
rect 33784 24760 33836 24769
rect 940 24556 992 24608
rect 9588 24599 9640 24608
rect 9588 24565 9597 24599
rect 9597 24565 9631 24599
rect 9631 24565 9640 24599
rect 9588 24556 9640 24565
rect 11244 24624 11296 24676
rect 13176 24624 13228 24676
rect 14372 24624 14424 24676
rect 14464 24667 14516 24676
rect 14464 24633 14473 24667
rect 14473 24633 14507 24667
rect 14507 24633 14516 24667
rect 14464 24624 14516 24633
rect 11888 24556 11940 24608
rect 13636 24556 13688 24608
rect 15016 24556 15068 24608
rect 17868 24692 17920 24744
rect 31116 24692 31168 24744
rect 33416 24735 33468 24744
rect 33416 24701 33425 24735
rect 33425 24701 33459 24735
rect 33459 24701 33468 24735
rect 33416 24692 33468 24701
rect 34888 24692 34940 24744
rect 18144 24624 18196 24676
rect 30932 24624 30984 24676
rect 18328 24556 18380 24608
rect 19248 24556 19300 24608
rect 20720 24556 20772 24608
rect 34152 24556 34204 24608
rect 36176 24828 36228 24880
rect 37096 24896 37148 24948
rect 38200 24939 38252 24948
rect 38200 24905 38209 24939
rect 38209 24905 38243 24939
rect 38243 24905 38252 24939
rect 38200 24896 38252 24905
rect 43076 24896 43128 24948
rect 44364 24896 44416 24948
rect 46388 24896 46440 24948
rect 51724 24896 51776 24948
rect 52000 24896 52052 24948
rect 36636 24803 36688 24812
rect 36636 24769 36645 24803
rect 36645 24769 36679 24803
rect 36679 24769 36688 24803
rect 36636 24760 36688 24769
rect 37556 24803 37608 24812
rect 37556 24769 37565 24803
rect 37565 24769 37599 24803
rect 37599 24769 37608 24803
rect 37556 24760 37608 24769
rect 37648 24760 37700 24812
rect 37280 24692 37332 24744
rect 37188 24624 37240 24676
rect 37924 24803 37976 24812
rect 37924 24769 37933 24803
rect 37933 24769 37967 24803
rect 37967 24769 37976 24803
rect 37924 24760 37976 24769
rect 41696 24828 41748 24880
rect 38752 24803 38804 24812
rect 38752 24769 38761 24803
rect 38761 24769 38795 24803
rect 38795 24769 38804 24803
rect 38752 24760 38804 24769
rect 39764 24760 39816 24812
rect 42616 24760 42668 24812
rect 42800 24803 42852 24812
rect 42800 24769 42809 24803
rect 42809 24769 42843 24803
rect 42843 24769 42852 24803
rect 42800 24760 42852 24769
rect 42892 24803 42944 24812
rect 42892 24769 42901 24803
rect 42901 24769 42935 24803
rect 42935 24769 42944 24803
rect 42892 24760 42944 24769
rect 43168 24760 43220 24812
rect 44088 24760 44140 24812
rect 43904 24692 43956 24744
rect 48412 24828 48464 24880
rect 50896 24828 50948 24880
rect 53564 24896 53616 24948
rect 54760 24939 54812 24948
rect 54760 24905 54769 24939
rect 54769 24905 54803 24939
rect 54803 24905 54812 24939
rect 54760 24896 54812 24905
rect 55588 24896 55640 24948
rect 53196 24828 53248 24880
rect 55772 24828 55824 24880
rect 44456 24760 44508 24812
rect 44824 24760 44876 24812
rect 45284 24760 45336 24812
rect 49424 24760 49476 24812
rect 43352 24624 43404 24676
rect 45468 24692 45520 24744
rect 48412 24692 48464 24744
rect 38936 24556 38988 24608
rect 42156 24556 42208 24608
rect 43444 24556 43496 24608
rect 43720 24556 43772 24608
rect 44088 24599 44140 24608
rect 44088 24565 44097 24599
rect 44097 24565 44131 24599
rect 44131 24565 44140 24599
rect 44088 24556 44140 24565
rect 49148 24556 49200 24608
rect 50804 24803 50856 24812
rect 50804 24769 50813 24803
rect 50813 24769 50847 24803
rect 50847 24769 50856 24803
rect 50804 24760 50856 24769
rect 51356 24760 51408 24812
rect 52092 24760 52144 24812
rect 52368 24760 52420 24812
rect 52552 24735 52604 24744
rect 52552 24701 52561 24735
rect 52561 24701 52595 24735
rect 52595 24701 52604 24735
rect 52552 24692 52604 24701
rect 53380 24692 53432 24744
rect 55312 24760 55364 24812
rect 55404 24803 55456 24812
rect 55404 24769 55413 24803
rect 55413 24769 55447 24803
rect 55447 24769 55456 24803
rect 55404 24760 55456 24769
rect 53012 24624 53064 24676
rect 54484 24692 54536 24744
rect 49516 24599 49568 24608
rect 49516 24565 49525 24599
rect 49525 24565 49559 24599
rect 49559 24565 49568 24599
rect 49516 24556 49568 24565
rect 55220 24599 55272 24608
rect 55220 24565 55229 24599
rect 55229 24565 55263 24599
rect 55263 24565 55272 24599
rect 55220 24556 55272 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 9036 24395 9088 24404
rect 9036 24361 9045 24395
rect 9045 24361 9079 24395
rect 9079 24361 9088 24395
rect 9036 24352 9088 24361
rect 13452 24352 13504 24404
rect 13820 24395 13872 24404
rect 13820 24361 13829 24395
rect 13829 24361 13863 24395
rect 13863 24361 13872 24395
rect 13820 24352 13872 24361
rect 14924 24352 14976 24404
rect 15108 24352 15160 24404
rect 30656 24352 30708 24404
rect 39672 24352 39724 24404
rect 43076 24352 43128 24404
rect 43904 24395 43956 24404
rect 43904 24361 43913 24395
rect 43913 24361 43947 24395
rect 43947 24361 43956 24395
rect 43904 24352 43956 24361
rect 48412 24395 48464 24404
rect 48412 24361 48421 24395
rect 48421 24361 48455 24395
rect 48455 24361 48464 24395
rect 48412 24352 48464 24361
rect 49424 24352 49476 24404
rect 11336 24284 11388 24336
rect 34796 24284 34848 24336
rect 37832 24284 37884 24336
rect 38200 24284 38252 24336
rect 42064 24284 42116 24336
rect 9588 24148 9640 24200
rect 10600 24148 10652 24200
rect 11060 24216 11112 24268
rect 11888 24259 11940 24268
rect 11888 24225 11897 24259
rect 11897 24225 11931 24259
rect 11931 24225 11940 24259
rect 11888 24216 11940 24225
rect 12532 24216 12584 24268
rect 14740 24259 14792 24268
rect 14740 24225 14749 24259
rect 14749 24225 14783 24259
rect 14783 24225 14792 24259
rect 14740 24216 14792 24225
rect 31392 24216 31444 24268
rect 10876 24191 10928 24200
rect 10876 24157 10885 24191
rect 10885 24157 10919 24191
rect 10919 24157 10928 24191
rect 10876 24148 10928 24157
rect 10968 24148 11020 24200
rect 10048 24123 10100 24132
rect 10048 24089 10057 24123
rect 10057 24089 10091 24123
rect 10091 24089 10100 24123
rect 10048 24080 10100 24089
rect 10416 24123 10468 24132
rect 10416 24089 10425 24123
rect 10425 24089 10459 24123
rect 10459 24089 10468 24123
rect 10416 24080 10468 24089
rect 2044 24055 2096 24064
rect 2044 24021 2053 24055
rect 2053 24021 2087 24055
rect 2087 24021 2096 24055
rect 2044 24012 2096 24021
rect 9036 24012 9088 24064
rect 11152 24080 11204 24132
rect 11244 24080 11296 24132
rect 13636 24191 13688 24200
rect 13636 24157 13645 24191
rect 13645 24157 13679 24191
rect 13679 24157 13688 24191
rect 13636 24148 13688 24157
rect 14372 24148 14424 24200
rect 17224 24148 17276 24200
rect 17500 24148 17552 24200
rect 18512 24148 18564 24200
rect 21088 24191 21140 24200
rect 21088 24157 21097 24191
rect 21097 24157 21131 24191
rect 21131 24157 21140 24191
rect 21088 24148 21140 24157
rect 31300 24191 31352 24200
rect 31300 24157 31309 24191
rect 31309 24157 31343 24191
rect 31343 24157 31352 24191
rect 31300 24148 31352 24157
rect 37096 24216 37148 24268
rect 31576 24148 31628 24200
rect 38844 24148 38896 24200
rect 42248 24148 42300 24200
rect 15016 24080 15068 24132
rect 13820 24012 13872 24064
rect 14924 24012 14976 24064
rect 17592 24012 17644 24064
rect 19524 24012 19576 24064
rect 31300 24012 31352 24064
rect 32772 24080 32824 24132
rect 33416 24080 33468 24132
rect 35992 24080 36044 24132
rect 37464 24080 37516 24132
rect 40040 24123 40092 24132
rect 40040 24089 40049 24123
rect 40049 24089 40083 24123
rect 40083 24089 40092 24123
rect 40040 24080 40092 24089
rect 35440 24012 35492 24064
rect 36452 24012 36504 24064
rect 36912 24012 36964 24064
rect 38200 24012 38252 24064
rect 39120 24012 39172 24064
rect 40408 24055 40460 24064
rect 40408 24021 40417 24055
rect 40417 24021 40451 24055
rect 40451 24021 40460 24055
rect 40408 24012 40460 24021
rect 42340 24055 42392 24064
rect 42340 24021 42349 24055
rect 42349 24021 42383 24055
rect 42383 24021 42392 24055
rect 42340 24012 42392 24021
rect 42616 24284 42668 24336
rect 45284 24284 45336 24336
rect 43260 24216 43312 24268
rect 45468 24259 45520 24268
rect 45468 24225 45477 24259
rect 45477 24225 45511 24259
rect 45511 24225 45520 24259
rect 45468 24216 45520 24225
rect 53288 24352 53340 24404
rect 53472 24352 53524 24404
rect 55404 24352 55456 24404
rect 52092 24284 52144 24336
rect 48504 24216 48556 24268
rect 42708 24191 42760 24200
rect 42708 24157 42717 24191
rect 42717 24157 42751 24191
rect 42751 24157 42760 24191
rect 42708 24148 42760 24157
rect 44364 24148 44416 24200
rect 44180 24080 44232 24132
rect 48412 24148 48464 24200
rect 49516 24216 49568 24268
rect 52368 24216 52420 24268
rect 45744 24123 45796 24132
rect 45744 24089 45753 24123
rect 45753 24089 45787 24123
rect 45787 24089 45796 24123
rect 45744 24080 45796 24089
rect 42892 24012 42944 24064
rect 44364 24012 44416 24064
rect 48596 24012 48648 24064
rect 49240 24191 49292 24200
rect 49240 24157 49249 24191
rect 49249 24157 49283 24191
rect 49283 24157 49292 24191
rect 49240 24148 49292 24157
rect 49424 24191 49476 24200
rect 49424 24157 49433 24191
rect 49433 24157 49467 24191
rect 49467 24157 49476 24191
rect 49424 24148 49476 24157
rect 49608 24191 49660 24200
rect 49608 24157 49617 24191
rect 49617 24157 49651 24191
rect 49651 24157 49660 24191
rect 49608 24148 49660 24157
rect 50068 24148 50120 24200
rect 48780 24080 48832 24132
rect 49884 24080 49936 24132
rect 51080 24123 51132 24132
rect 51080 24089 51089 24123
rect 51089 24089 51123 24123
rect 51123 24089 51132 24123
rect 51080 24080 51132 24089
rect 52920 24148 52972 24200
rect 54944 24216 54996 24268
rect 53012 24123 53064 24132
rect 53012 24089 53021 24123
rect 53021 24089 53055 24123
rect 53055 24089 53064 24123
rect 53012 24080 53064 24089
rect 54760 24148 54812 24200
rect 54944 24080 54996 24132
rect 52552 24055 52604 24064
rect 52552 24021 52561 24055
rect 52561 24021 52595 24055
rect 52595 24021 52604 24055
rect 52552 24012 52604 24021
rect 53748 24012 53800 24064
rect 55588 24123 55640 24132
rect 55588 24089 55597 24123
rect 55597 24089 55631 24123
rect 55631 24089 55640 24123
rect 55588 24080 55640 24089
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 66314 23910 66366 23962
rect 66378 23910 66430 23962
rect 66442 23910 66494 23962
rect 66506 23910 66558 23962
rect 66570 23910 66622 23962
rect 1308 23808 1360 23860
rect 2044 23715 2096 23724
rect 2044 23681 2053 23715
rect 2053 23681 2087 23715
rect 2087 23681 2096 23715
rect 2044 23672 2096 23681
rect 7748 23672 7800 23724
rect 9680 23808 9732 23860
rect 10968 23808 11020 23860
rect 14280 23808 14332 23860
rect 9036 23783 9088 23792
rect 9036 23749 9045 23783
rect 9045 23749 9079 23783
rect 9079 23749 9088 23783
rect 9036 23740 9088 23749
rect 10324 23740 10376 23792
rect 10600 23783 10652 23792
rect 10600 23749 10609 23783
rect 10609 23749 10643 23783
rect 10643 23749 10652 23783
rect 10600 23740 10652 23749
rect 17684 23808 17736 23860
rect 21088 23808 21140 23860
rect 17592 23783 17644 23792
rect 17592 23749 17601 23783
rect 17601 23749 17635 23783
rect 17635 23749 17644 23783
rect 17592 23740 17644 23749
rect 18052 23740 18104 23792
rect 2136 23647 2188 23656
rect 2136 23613 2145 23647
rect 2145 23613 2179 23647
rect 2179 23613 2188 23647
rect 2136 23604 2188 23613
rect 10876 23672 10928 23724
rect 11152 23672 11204 23724
rect 16948 23715 17000 23724
rect 16948 23681 16957 23715
rect 16957 23681 16991 23715
rect 16991 23681 17000 23715
rect 16948 23672 17000 23681
rect 17040 23715 17092 23724
rect 17040 23681 17049 23715
rect 17049 23681 17083 23715
rect 17083 23681 17092 23715
rect 17040 23672 17092 23681
rect 19524 23672 19576 23724
rect 11060 23536 11112 23588
rect 10876 23468 10928 23520
rect 14464 23604 14516 23656
rect 16672 23604 16724 23656
rect 17224 23579 17276 23588
rect 17224 23545 17233 23579
rect 17233 23545 17267 23579
rect 17267 23545 17276 23579
rect 17224 23536 17276 23545
rect 17592 23604 17644 23656
rect 19248 23604 19300 23656
rect 22836 23808 22888 23860
rect 30104 23808 30156 23860
rect 30932 23808 30984 23860
rect 30840 23740 30892 23792
rect 34152 23740 34204 23792
rect 34704 23740 34756 23792
rect 35440 23740 35492 23792
rect 37096 23851 37148 23860
rect 28448 23672 28500 23724
rect 31300 23672 31352 23724
rect 30472 23647 30524 23656
rect 30472 23613 30481 23647
rect 30481 23613 30515 23647
rect 30515 23613 30524 23647
rect 30472 23604 30524 23613
rect 30840 23604 30892 23656
rect 32128 23604 32180 23656
rect 32772 23647 32824 23656
rect 32772 23613 32781 23647
rect 32781 23613 32815 23647
rect 32815 23613 32824 23647
rect 32772 23604 32824 23613
rect 33140 23647 33192 23656
rect 33140 23613 33149 23647
rect 33149 23613 33183 23647
rect 33183 23613 33192 23647
rect 33140 23604 33192 23613
rect 34796 23672 34848 23724
rect 33324 23604 33376 23656
rect 30380 23468 30432 23520
rect 31024 23468 31076 23520
rect 32956 23468 33008 23520
rect 33968 23536 34020 23588
rect 35256 23715 35308 23724
rect 35256 23681 35265 23715
rect 35265 23681 35299 23715
rect 35299 23681 35308 23715
rect 35256 23672 35308 23681
rect 35348 23715 35400 23724
rect 35348 23681 35357 23715
rect 35357 23681 35391 23715
rect 35391 23681 35400 23715
rect 35348 23672 35400 23681
rect 35992 23740 36044 23792
rect 37096 23817 37105 23851
rect 37105 23817 37139 23851
rect 37139 23817 37148 23851
rect 37096 23808 37148 23817
rect 38200 23851 38252 23860
rect 37188 23740 37240 23792
rect 37556 23783 37608 23792
rect 37556 23749 37565 23783
rect 37565 23749 37599 23783
rect 37599 23749 37608 23783
rect 37556 23740 37608 23749
rect 38200 23817 38209 23851
rect 38209 23817 38243 23851
rect 38243 23817 38252 23851
rect 38200 23808 38252 23817
rect 39212 23808 39264 23860
rect 40040 23808 40092 23860
rect 43812 23808 43864 23860
rect 45744 23808 45796 23860
rect 49332 23808 49384 23860
rect 52092 23808 52144 23860
rect 36084 23536 36136 23588
rect 37832 23715 37884 23724
rect 37832 23681 37841 23715
rect 37841 23681 37875 23715
rect 37875 23681 37884 23715
rect 37832 23672 37884 23681
rect 39488 23740 39540 23792
rect 42064 23740 42116 23792
rect 42708 23740 42760 23792
rect 39120 23715 39172 23724
rect 39120 23681 39129 23715
rect 39129 23681 39163 23715
rect 39163 23681 39172 23715
rect 39120 23672 39172 23681
rect 37372 23604 37424 23656
rect 40316 23672 40368 23724
rect 39672 23647 39724 23656
rect 39672 23613 39681 23647
rect 39681 23613 39715 23647
rect 39715 23613 39724 23647
rect 39672 23604 39724 23613
rect 43720 23672 43772 23724
rect 44180 23672 44232 23724
rect 44640 23740 44692 23792
rect 45284 23740 45336 23792
rect 44364 23715 44416 23724
rect 44364 23681 44373 23715
rect 44373 23681 44407 23715
rect 44407 23681 44416 23715
rect 44364 23672 44416 23681
rect 44456 23715 44508 23724
rect 44456 23681 44465 23715
rect 44465 23681 44499 23715
rect 44499 23681 44508 23715
rect 44456 23672 44508 23681
rect 46388 23715 46440 23724
rect 46388 23681 46397 23715
rect 46397 23681 46431 23715
rect 46431 23681 46440 23715
rect 46388 23672 46440 23681
rect 48412 23740 48464 23792
rect 52552 23740 52604 23792
rect 48320 23715 48372 23724
rect 48320 23681 48329 23715
rect 48329 23681 48363 23715
rect 48363 23681 48372 23715
rect 48320 23672 48372 23681
rect 48964 23672 49016 23724
rect 50528 23672 50580 23724
rect 50712 23672 50764 23724
rect 43628 23604 43680 23656
rect 45836 23647 45888 23656
rect 45836 23613 45845 23647
rect 45845 23613 45879 23647
rect 45879 23613 45888 23647
rect 45836 23604 45888 23613
rect 38476 23536 38528 23588
rect 42248 23536 42300 23588
rect 34704 23511 34756 23520
rect 34704 23477 34713 23511
rect 34713 23477 34747 23511
rect 34747 23477 34756 23511
rect 34704 23468 34756 23477
rect 36728 23511 36780 23520
rect 36728 23477 36737 23511
rect 36737 23477 36771 23511
rect 36771 23477 36780 23511
rect 36728 23468 36780 23477
rect 37280 23511 37332 23520
rect 37280 23477 37289 23511
rect 37289 23477 37323 23511
rect 37323 23477 37332 23511
rect 37280 23468 37332 23477
rect 41696 23468 41748 23520
rect 44180 23468 44232 23520
rect 44456 23468 44508 23520
rect 48044 23511 48096 23520
rect 48044 23477 48053 23511
rect 48053 23477 48087 23511
rect 48087 23477 48096 23511
rect 48044 23468 48096 23477
rect 48504 23647 48556 23656
rect 48504 23613 48513 23647
rect 48513 23613 48547 23647
rect 48547 23613 48556 23647
rect 48504 23604 48556 23613
rect 49240 23604 49292 23656
rect 49424 23647 49476 23656
rect 49424 23613 49433 23647
rect 49433 23613 49467 23647
rect 49467 23613 49476 23647
rect 49424 23604 49476 23613
rect 50252 23647 50304 23656
rect 50252 23613 50261 23647
rect 50261 23613 50295 23647
rect 50295 23613 50304 23647
rect 52920 23672 52972 23724
rect 55312 23740 55364 23792
rect 50252 23604 50304 23613
rect 49056 23536 49108 23588
rect 50528 23579 50580 23588
rect 50528 23545 50537 23579
rect 50537 23545 50571 23579
rect 50571 23545 50580 23579
rect 53748 23604 53800 23656
rect 54576 23715 54628 23724
rect 54576 23681 54585 23715
rect 54585 23681 54619 23715
rect 54619 23681 54628 23715
rect 54576 23672 54628 23681
rect 54944 23672 54996 23724
rect 58532 23672 58584 23724
rect 50528 23536 50580 23545
rect 56048 23536 56100 23588
rect 51080 23468 51132 23520
rect 55128 23468 55180 23520
rect 78220 23511 78272 23520
rect 78220 23477 78229 23511
rect 78229 23477 78263 23511
rect 78263 23477 78272 23511
rect 78220 23468 78272 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 17500 23264 17552 23316
rect 1216 23196 1268 23248
rect 17040 23196 17092 23248
rect 17776 23264 17828 23316
rect 10876 23171 10928 23180
rect 10876 23137 10885 23171
rect 10885 23137 10919 23171
rect 10919 23137 10928 23171
rect 10876 23128 10928 23137
rect 11152 23171 11204 23180
rect 11152 23137 11161 23171
rect 11161 23137 11195 23171
rect 11195 23137 11204 23171
rect 11152 23128 11204 23137
rect 15476 23128 15528 23180
rect 18236 23128 18288 23180
rect 2136 23103 2188 23112
rect 2136 23069 2145 23103
rect 2145 23069 2179 23103
rect 2179 23069 2188 23103
rect 2136 23060 2188 23069
rect 10692 23060 10744 23112
rect 14464 23060 14516 23112
rect 19340 23264 19392 23316
rect 30012 23264 30064 23316
rect 30380 23264 30432 23316
rect 30472 23264 30524 23316
rect 31116 23264 31168 23316
rect 32588 23264 32640 23316
rect 33140 23264 33192 23316
rect 35992 23264 36044 23316
rect 36176 23264 36228 23316
rect 40316 23264 40368 23316
rect 42340 23264 42392 23316
rect 13728 22992 13780 23044
rect 16672 22992 16724 23044
rect 17684 22992 17736 23044
rect 19156 22992 19208 23044
rect 30288 23128 30340 23180
rect 29828 23060 29880 23112
rect 29920 23060 29972 23112
rect 30104 23103 30156 23112
rect 30104 23069 30113 23103
rect 30113 23069 30147 23103
rect 30147 23069 30156 23103
rect 30104 23060 30156 23069
rect 31392 23196 31444 23248
rect 32864 23196 32916 23248
rect 31208 23128 31260 23180
rect 32588 23128 32640 23180
rect 30380 23035 30432 23044
rect 30380 23001 30389 23035
rect 30389 23001 30423 23035
rect 30423 23001 30432 23035
rect 30380 22992 30432 23001
rect 940 22924 992 22976
rect 13084 22924 13136 22976
rect 16948 22924 17000 22976
rect 17592 22967 17644 22976
rect 17592 22933 17609 22967
rect 17609 22933 17644 22967
rect 17592 22924 17644 22933
rect 18604 22924 18656 22976
rect 19248 22924 19300 22976
rect 30104 22924 30156 22976
rect 30656 23060 30708 23112
rect 31300 23103 31352 23112
rect 31300 23069 31309 23103
rect 31309 23069 31343 23103
rect 31343 23069 31352 23103
rect 31300 23060 31352 23069
rect 31852 23060 31904 23112
rect 32312 23060 32364 23112
rect 31760 22992 31812 23044
rect 33232 22992 33284 23044
rect 34796 23060 34848 23112
rect 35348 23060 35400 23112
rect 36176 23128 36228 23180
rect 39948 23196 40000 23248
rect 48228 23264 48280 23316
rect 48320 23264 48372 23316
rect 50896 23264 50948 23316
rect 51540 23264 51592 23316
rect 51908 23264 51960 23316
rect 55220 23264 55272 23316
rect 55312 23307 55364 23316
rect 55312 23273 55321 23307
rect 55321 23273 55355 23307
rect 55355 23273 55364 23307
rect 55312 23264 55364 23273
rect 55588 23264 55640 23316
rect 58532 23307 58584 23316
rect 58532 23273 58541 23307
rect 58541 23273 58575 23307
rect 58575 23273 58584 23307
rect 58532 23264 58584 23273
rect 37280 23128 37332 23180
rect 39764 23128 39816 23180
rect 42708 23196 42760 23248
rect 34704 22992 34756 23044
rect 36544 23103 36596 23112
rect 36544 23069 36553 23103
rect 36553 23069 36587 23103
rect 36587 23069 36596 23103
rect 36544 23060 36596 23069
rect 36820 23060 36872 23112
rect 39120 23060 39172 23112
rect 42524 23128 42576 23180
rect 43076 23171 43128 23180
rect 43076 23137 43085 23171
rect 43085 23137 43119 23171
rect 43119 23137 43128 23171
rect 43076 23128 43128 23137
rect 44088 23128 44140 23180
rect 44272 23171 44324 23180
rect 44272 23137 44281 23171
rect 44281 23137 44315 23171
rect 44315 23137 44324 23171
rect 44272 23128 44324 23137
rect 44732 23128 44784 23180
rect 31576 22924 31628 22976
rect 37188 22992 37240 23044
rect 39580 22992 39632 23044
rect 36176 22967 36228 22976
rect 36176 22933 36185 22967
rect 36185 22933 36219 22967
rect 36219 22933 36228 22967
rect 36176 22924 36228 22933
rect 36544 22924 36596 22976
rect 40224 23035 40276 23044
rect 40224 23001 40233 23035
rect 40233 23001 40267 23035
rect 40267 23001 40276 23035
rect 40224 22992 40276 23001
rect 40500 22924 40552 22976
rect 42248 23103 42300 23112
rect 42248 23069 42257 23103
rect 42257 23069 42291 23103
rect 42291 23069 42300 23103
rect 42248 23060 42300 23069
rect 42984 23060 43036 23112
rect 43628 23060 43680 23112
rect 43812 23103 43864 23112
rect 43812 23069 43821 23103
rect 43821 23069 43855 23103
rect 43855 23069 43864 23103
rect 43812 23060 43864 23069
rect 43904 23103 43956 23112
rect 43904 23069 43913 23103
rect 43913 23069 43947 23103
rect 43947 23069 43956 23103
rect 43904 23060 43956 23069
rect 45192 23171 45244 23180
rect 45192 23137 45201 23171
rect 45201 23137 45235 23171
rect 45235 23137 45244 23171
rect 45192 23128 45244 23137
rect 45376 23196 45428 23248
rect 49056 23196 49108 23248
rect 48044 23128 48096 23180
rect 48596 23128 48648 23180
rect 49148 23128 49200 23180
rect 42524 22992 42576 23044
rect 42892 22992 42944 23044
rect 42616 22924 42668 22976
rect 43444 22924 43496 22976
rect 45376 23103 45428 23112
rect 45376 23069 45385 23103
rect 45385 23069 45419 23103
rect 45419 23069 45428 23103
rect 45376 23060 45428 23069
rect 46020 23060 46072 23112
rect 46388 23103 46440 23112
rect 46388 23069 46397 23103
rect 46397 23069 46431 23103
rect 46431 23069 46440 23103
rect 46388 23060 46440 23069
rect 47308 23103 47360 23112
rect 47308 23069 47317 23103
rect 47317 23069 47351 23103
rect 47351 23069 47360 23103
rect 47308 23060 47360 23069
rect 48688 23060 48740 23112
rect 49332 23103 49384 23112
rect 49332 23069 49341 23103
rect 49341 23069 49375 23103
rect 49375 23069 49384 23103
rect 49332 23060 49384 23069
rect 44732 22992 44784 23044
rect 45192 22992 45244 23044
rect 46664 22992 46716 23044
rect 50620 23060 50672 23112
rect 51080 23103 51132 23112
rect 51080 23069 51089 23103
rect 51089 23069 51123 23103
rect 51123 23069 51132 23103
rect 51080 23060 51132 23069
rect 52920 23128 52972 23180
rect 51540 23103 51592 23112
rect 51540 23069 51554 23103
rect 51554 23069 51588 23103
rect 51588 23069 51592 23103
rect 51540 23060 51592 23069
rect 52276 23060 52328 23112
rect 53196 23103 53248 23112
rect 53196 23069 53205 23103
rect 53205 23069 53239 23103
rect 53239 23069 53248 23103
rect 53196 23060 53248 23069
rect 44640 22967 44692 22976
rect 44640 22933 44649 22967
rect 44649 22933 44683 22967
rect 44683 22933 44692 22967
rect 44640 22924 44692 22933
rect 45008 22967 45060 22976
rect 45008 22933 45017 22967
rect 45017 22933 45051 22967
rect 45051 22933 45060 22967
rect 45008 22924 45060 22933
rect 45100 22924 45152 22976
rect 49884 22992 49936 23044
rect 50896 23035 50948 23044
rect 50896 23001 50905 23035
rect 50905 23001 50939 23035
rect 50939 23001 50948 23035
rect 50896 22992 50948 23001
rect 49240 22924 49292 22976
rect 49700 22967 49752 22976
rect 49700 22933 49709 22967
rect 49709 22933 49743 22967
rect 49743 22933 49752 22967
rect 49700 22924 49752 22933
rect 50160 22924 50212 22976
rect 50712 22967 50764 22976
rect 50712 22933 50721 22967
rect 50721 22933 50755 22967
rect 50755 22933 50764 22967
rect 52552 22992 52604 23044
rect 54484 23128 54536 23180
rect 56232 23128 56284 23180
rect 54576 23103 54628 23112
rect 54576 23069 54585 23103
rect 54585 23069 54619 23103
rect 54619 23069 54628 23103
rect 54576 23060 54628 23069
rect 57060 23103 57112 23112
rect 57060 23069 57069 23103
rect 57069 23069 57103 23103
rect 57103 23069 57112 23103
rect 57060 23060 57112 23069
rect 56232 22992 56284 23044
rect 50712 22924 50764 22933
rect 51540 22924 51592 22976
rect 53012 22924 53064 22976
rect 54852 22924 54904 22976
rect 55312 22924 55364 22976
rect 55404 22924 55456 22976
rect 56876 22992 56928 23044
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 66314 22822 66366 22874
rect 66378 22822 66430 22874
rect 66442 22822 66494 22874
rect 66506 22822 66558 22874
rect 66570 22822 66622 22874
rect 10692 22763 10744 22772
rect 10692 22729 10701 22763
rect 10701 22729 10735 22763
rect 10735 22729 10744 22763
rect 10692 22720 10744 22729
rect 14464 22720 14516 22772
rect 17132 22720 17184 22772
rect 17868 22720 17920 22772
rect 19248 22720 19300 22772
rect 9680 22695 9732 22704
rect 9680 22661 9689 22695
rect 9689 22661 9723 22695
rect 9723 22661 9732 22695
rect 9680 22652 9732 22661
rect 13728 22652 13780 22704
rect 15476 22695 15528 22704
rect 15476 22661 15485 22695
rect 15485 22661 15519 22695
rect 15519 22661 15528 22695
rect 15476 22652 15528 22661
rect 18236 22652 18288 22704
rect 30472 22720 30524 22772
rect 30840 22720 30892 22772
rect 32036 22720 32088 22772
rect 32680 22720 32732 22772
rect 13084 22627 13136 22636
rect 13084 22593 13093 22627
rect 13093 22593 13127 22627
rect 13127 22593 13136 22627
rect 13084 22584 13136 22593
rect 18052 22584 18104 22636
rect 18604 22584 18656 22636
rect 28448 22584 28500 22636
rect 30104 22627 30156 22636
rect 30104 22593 30113 22627
rect 30113 22593 30147 22627
rect 30147 22593 30156 22627
rect 30104 22584 30156 22593
rect 30196 22627 30248 22636
rect 30196 22593 30205 22627
rect 30205 22593 30239 22627
rect 30239 22593 30248 22627
rect 30196 22584 30248 22593
rect 11060 22516 11112 22568
rect 12440 22516 12492 22568
rect 12900 22516 12952 22568
rect 15108 22559 15160 22568
rect 15108 22525 15117 22559
rect 15117 22525 15151 22559
rect 15151 22525 15160 22559
rect 15108 22516 15160 22525
rect 16672 22559 16724 22568
rect 14096 22448 14148 22500
rect 14372 22380 14424 22432
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 16948 22559 17000 22568
rect 16948 22525 16957 22559
rect 16957 22525 16991 22559
rect 16991 22525 17000 22559
rect 16948 22516 17000 22525
rect 17960 22516 18012 22568
rect 29552 22516 29604 22568
rect 29920 22516 29972 22568
rect 30380 22584 30432 22636
rect 30656 22584 30708 22636
rect 31852 22584 31904 22636
rect 32312 22627 32364 22636
rect 32312 22593 32321 22627
rect 32321 22593 32355 22627
rect 32355 22593 32364 22627
rect 32312 22584 32364 22593
rect 32864 22652 32916 22704
rect 32680 22627 32732 22636
rect 32680 22593 32689 22627
rect 32689 22593 32723 22627
rect 32723 22593 32732 22627
rect 32680 22584 32732 22593
rect 32956 22627 33008 22636
rect 32956 22593 32965 22627
rect 32965 22593 32999 22627
rect 32999 22593 33008 22627
rect 32956 22584 33008 22593
rect 33048 22627 33100 22636
rect 33048 22593 33057 22627
rect 33057 22593 33091 22627
rect 33091 22593 33100 22627
rect 33324 22627 33376 22636
rect 33048 22584 33100 22593
rect 33324 22593 33347 22627
rect 33347 22593 33376 22627
rect 33324 22584 33376 22593
rect 33784 22584 33836 22636
rect 32036 22516 32088 22568
rect 35624 22584 35676 22636
rect 36544 22627 36596 22636
rect 36544 22593 36553 22627
rect 36553 22593 36587 22627
rect 36587 22593 36596 22627
rect 36544 22584 36596 22593
rect 38384 22720 38436 22772
rect 37740 22695 37792 22704
rect 37740 22661 37749 22695
rect 37749 22661 37783 22695
rect 37783 22661 37792 22695
rect 37740 22652 37792 22661
rect 38108 22652 38160 22704
rect 38200 22652 38252 22704
rect 39120 22763 39172 22772
rect 39120 22729 39129 22763
rect 39129 22729 39163 22763
rect 39163 22729 39172 22763
rect 39120 22720 39172 22729
rect 39948 22763 40000 22772
rect 39948 22729 39957 22763
rect 39957 22729 39991 22763
rect 39991 22729 40000 22763
rect 39948 22720 40000 22729
rect 40224 22720 40276 22772
rect 41236 22720 41288 22772
rect 39212 22695 39264 22704
rect 39212 22661 39221 22695
rect 39221 22661 39255 22695
rect 39255 22661 39264 22695
rect 39212 22652 39264 22661
rect 41512 22720 41564 22772
rect 42064 22720 42116 22772
rect 44180 22720 44232 22772
rect 45192 22720 45244 22772
rect 48228 22720 48280 22772
rect 38292 22584 38344 22636
rect 38752 22584 38804 22636
rect 39580 22627 39632 22636
rect 39580 22593 39589 22627
rect 39589 22593 39623 22627
rect 39623 22593 39632 22627
rect 39580 22584 39632 22593
rect 42340 22584 42392 22636
rect 42616 22627 42668 22636
rect 42616 22593 42625 22627
rect 42625 22593 42659 22627
rect 42659 22593 42668 22627
rect 42616 22584 42668 22593
rect 42708 22627 42760 22636
rect 42708 22593 42717 22627
rect 42717 22593 42751 22627
rect 42751 22593 42760 22627
rect 42708 22584 42760 22593
rect 44364 22652 44416 22704
rect 44640 22652 44692 22704
rect 48136 22652 48188 22704
rect 45008 22584 45060 22636
rect 45744 22584 45796 22636
rect 48320 22584 48372 22636
rect 48596 22627 48648 22636
rect 48596 22593 48603 22627
rect 48603 22593 48648 22627
rect 48596 22584 48648 22593
rect 50620 22720 50672 22772
rect 30104 22448 30156 22500
rect 33048 22448 33100 22500
rect 38660 22516 38712 22568
rect 43168 22559 43220 22568
rect 43168 22525 43177 22559
rect 43177 22525 43211 22559
rect 43211 22525 43220 22559
rect 43168 22516 43220 22525
rect 43536 22559 43588 22568
rect 43536 22525 43545 22559
rect 43545 22525 43579 22559
rect 43579 22525 43588 22559
rect 43536 22516 43588 22525
rect 44272 22516 44324 22568
rect 47216 22516 47268 22568
rect 47952 22516 48004 22568
rect 37372 22448 37424 22500
rect 37832 22448 37884 22500
rect 29920 22423 29972 22432
rect 29920 22389 29929 22423
rect 29929 22389 29963 22423
rect 29963 22389 29972 22423
rect 29920 22380 29972 22389
rect 30196 22380 30248 22432
rect 31116 22380 31168 22432
rect 32404 22380 32456 22432
rect 32588 22423 32640 22432
rect 32588 22389 32597 22423
rect 32597 22389 32631 22423
rect 32631 22389 32640 22423
rect 32588 22380 32640 22389
rect 32680 22380 32732 22432
rect 33784 22380 33836 22432
rect 35624 22423 35676 22432
rect 35624 22389 35633 22423
rect 35633 22389 35667 22423
rect 35667 22389 35676 22423
rect 35624 22380 35676 22389
rect 36728 22423 36780 22432
rect 36728 22389 36737 22423
rect 36737 22389 36771 22423
rect 36771 22389 36780 22423
rect 36728 22380 36780 22389
rect 40224 22423 40276 22432
rect 40224 22389 40233 22423
rect 40233 22389 40267 22423
rect 40267 22389 40276 22423
rect 40224 22380 40276 22389
rect 40500 22380 40552 22432
rect 44916 22380 44968 22432
rect 49516 22516 49568 22568
rect 49700 22627 49752 22636
rect 49700 22593 49709 22627
rect 49709 22593 49743 22627
rect 49743 22593 49752 22627
rect 49700 22584 49752 22593
rect 49792 22627 49844 22636
rect 49792 22593 49802 22627
rect 49802 22593 49836 22627
rect 49836 22593 49844 22627
rect 49792 22584 49844 22593
rect 48596 22380 48648 22432
rect 49792 22448 49844 22500
rect 49516 22380 49568 22432
rect 49976 22448 50028 22500
rect 50160 22627 50212 22636
rect 53012 22695 53064 22704
rect 53012 22661 53021 22695
rect 53021 22661 53055 22695
rect 53055 22661 53064 22695
rect 53012 22652 53064 22661
rect 54484 22652 54536 22704
rect 55404 22695 55456 22704
rect 55404 22661 55413 22695
rect 55413 22661 55447 22695
rect 55447 22661 55456 22695
rect 55404 22652 55456 22661
rect 56048 22695 56100 22704
rect 56048 22661 56057 22695
rect 56057 22661 56091 22695
rect 56091 22661 56100 22695
rect 56048 22652 56100 22661
rect 50160 22593 50174 22627
rect 50174 22593 50208 22627
rect 50208 22593 50212 22627
rect 50160 22584 50212 22593
rect 50988 22627 51040 22636
rect 50988 22593 51002 22627
rect 51002 22593 51036 22627
rect 51036 22593 51040 22627
rect 50988 22584 51040 22593
rect 51172 22584 51224 22636
rect 51356 22559 51408 22568
rect 51356 22525 51365 22559
rect 51365 22525 51399 22559
rect 51399 22525 51408 22559
rect 51356 22516 51408 22525
rect 51540 22627 51592 22636
rect 51540 22593 51549 22627
rect 51549 22593 51583 22627
rect 51583 22593 51592 22627
rect 51540 22584 51592 22593
rect 54852 22627 54904 22636
rect 54852 22593 54861 22627
rect 54861 22593 54895 22627
rect 54895 22593 54904 22627
rect 54852 22584 54904 22593
rect 55128 22627 55180 22636
rect 55128 22593 55137 22627
rect 55137 22593 55171 22627
rect 55171 22593 55180 22627
rect 55128 22584 55180 22593
rect 52644 22516 52696 22568
rect 52736 22559 52788 22568
rect 52736 22525 52745 22559
rect 52745 22525 52779 22559
rect 52779 22525 52788 22559
rect 52736 22516 52788 22525
rect 56876 22763 56928 22772
rect 56876 22729 56885 22763
rect 56885 22729 56919 22763
rect 56919 22729 56928 22763
rect 56876 22720 56928 22729
rect 58532 22720 58584 22772
rect 56324 22584 56376 22636
rect 50160 22380 50212 22432
rect 54116 22448 54168 22500
rect 55220 22448 55272 22500
rect 54484 22423 54536 22432
rect 54484 22389 54493 22423
rect 54493 22389 54527 22423
rect 54527 22389 54536 22423
rect 54484 22380 54536 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 11152 22176 11204 22228
rect 15108 22176 15160 22228
rect 16948 22176 17000 22228
rect 29828 22176 29880 22228
rect 30012 22219 30064 22228
rect 30012 22185 30021 22219
rect 30021 22185 30055 22219
rect 30055 22185 30064 22219
rect 30012 22176 30064 22185
rect 31116 22176 31168 22228
rect 38200 22176 38252 22228
rect 12992 22151 13044 22160
rect 12992 22117 13001 22151
rect 13001 22117 13035 22151
rect 13035 22117 13044 22151
rect 12992 22108 13044 22117
rect 30196 22108 30248 22160
rect 30472 22151 30524 22160
rect 30472 22117 30481 22151
rect 30481 22117 30515 22151
rect 30515 22117 30524 22151
rect 30472 22108 30524 22117
rect 30564 22108 30616 22160
rect 31208 22108 31260 22160
rect 35624 22108 35676 22160
rect 40592 22176 40644 22228
rect 44272 22176 44324 22228
rect 45284 22176 45336 22228
rect 9680 22040 9732 22092
rect 12440 22040 12492 22092
rect 14096 22040 14148 22092
rect 17500 22040 17552 22092
rect 18604 22083 18656 22092
rect 18604 22049 18613 22083
rect 18613 22049 18647 22083
rect 18647 22049 18656 22083
rect 18604 22040 18656 22049
rect 29552 22083 29604 22092
rect 29552 22049 29561 22083
rect 29561 22049 29595 22083
rect 29595 22049 29604 22083
rect 29552 22040 29604 22049
rect 7012 21972 7064 22024
rect 17132 21972 17184 22024
rect 10048 21904 10100 21956
rect 29920 21972 29972 22024
rect 30104 22015 30156 22024
rect 30104 21981 30113 22015
rect 30113 21981 30147 22015
rect 30147 21981 30156 22015
rect 30104 21972 30156 21981
rect 30288 22015 30340 22024
rect 30288 21981 30297 22015
rect 30297 21981 30331 22015
rect 30331 21981 30340 22015
rect 31116 22015 31168 22024
rect 30288 21972 30340 21981
rect 31116 21981 31125 22015
rect 31125 21981 31159 22015
rect 31159 21981 31168 22015
rect 31116 21972 31168 21981
rect 30656 21904 30708 21956
rect 30748 21904 30800 21956
rect 32128 21972 32180 22024
rect 32404 22083 32456 22092
rect 32404 22049 32413 22083
rect 32413 22049 32447 22083
rect 32447 22049 32456 22083
rect 32404 22040 32456 22049
rect 33784 22040 33836 22092
rect 37188 22040 37240 22092
rect 43996 22108 44048 22160
rect 45192 22108 45244 22160
rect 47216 22176 47268 22228
rect 47400 22176 47452 22228
rect 46756 22108 46808 22160
rect 49700 22176 49752 22228
rect 49976 22176 50028 22228
rect 50160 22176 50212 22228
rect 53196 22176 53248 22228
rect 34612 21972 34664 22024
rect 31944 21904 31996 21956
rect 33416 21904 33468 21956
rect 35992 21904 36044 21956
rect 41604 21904 41656 21956
rect 41788 21947 41840 21956
rect 41788 21913 41797 21947
rect 41797 21913 41831 21947
rect 41831 21913 41840 21947
rect 41788 21904 41840 21913
rect 41972 21904 42024 21956
rect 42156 21947 42208 21956
rect 42156 21913 42165 21947
rect 42165 21913 42199 21947
rect 42199 21913 42208 21947
rect 42156 21904 42208 21913
rect 42524 22040 42576 22092
rect 43076 22040 43128 22092
rect 43904 22040 43956 22092
rect 42616 22015 42668 22024
rect 42616 21981 42625 22015
rect 42625 21981 42659 22015
rect 42659 21981 42668 22015
rect 42616 21972 42668 21981
rect 42800 21904 42852 21956
rect 848 21836 900 21888
rect 11060 21836 11112 21888
rect 13912 21836 13964 21888
rect 29736 21836 29788 21888
rect 34244 21836 34296 21888
rect 37464 21836 37516 21888
rect 37924 21836 37976 21888
rect 38292 21879 38344 21888
rect 38292 21845 38301 21879
rect 38301 21845 38335 21879
rect 38335 21845 38344 21879
rect 38292 21836 38344 21845
rect 38660 21836 38712 21888
rect 39856 21836 39908 21888
rect 42984 21947 43036 21956
rect 42984 21913 42993 21947
rect 42993 21913 43027 21947
rect 43027 21913 43036 21947
rect 42984 21904 43036 21913
rect 43076 21947 43128 21956
rect 43076 21913 43085 21947
rect 43085 21913 43119 21947
rect 43119 21913 43128 21947
rect 43076 21904 43128 21913
rect 47400 22083 47452 22092
rect 47400 22049 47409 22083
rect 47409 22049 47443 22083
rect 47443 22049 47452 22083
rect 47400 22040 47452 22049
rect 49700 22040 49752 22092
rect 49792 22040 49844 22092
rect 50988 22040 51040 22092
rect 52552 22040 52604 22092
rect 43352 21947 43404 21956
rect 43352 21913 43361 21947
rect 43361 21913 43395 21947
rect 43395 21913 43404 21947
rect 43352 21904 43404 21913
rect 43536 21904 43588 21956
rect 43904 21904 43956 21956
rect 45100 21904 45152 21956
rect 45560 21904 45612 21956
rect 45744 21947 45796 21956
rect 45744 21913 45753 21947
rect 45753 21913 45787 21947
rect 45787 21913 45796 21947
rect 45744 21904 45796 21913
rect 44272 21836 44324 21888
rect 46388 21972 46440 22024
rect 47032 21972 47084 22024
rect 49240 22015 49292 22024
rect 49240 21981 49249 22015
rect 49249 21981 49283 22015
rect 49283 21981 49292 22015
rect 49240 21972 49292 21981
rect 49608 22015 49660 22024
rect 49608 21981 49617 22015
rect 49617 21981 49651 22015
rect 49651 21981 49660 22015
rect 49608 21972 49660 21981
rect 52644 21972 52696 22024
rect 52920 22040 52972 22092
rect 56968 22040 57020 22092
rect 53012 22015 53064 22024
rect 53012 21981 53021 22015
rect 53021 21981 53055 22015
rect 53055 21981 53064 22015
rect 53012 21972 53064 21981
rect 54944 21972 54996 22024
rect 47768 21904 47820 21956
rect 48872 21904 48924 21956
rect 49332 21904 49384 21956
rect 52828 21904 52880 21956
rect 46940 21836 46992 21888
rect 48136 21836 48188 21888
rect 49884 21836 49936 21888
rect 50160 21879 50212 21888
rect 50160 21845 50169 21879
rect 50169 21845 50203 21879
rect 50203 21845 50212 21879
rect 50160 21836 50212 21845
rect 50620 21836 50672 21888
rect 53380 21947 53432 21956
rect 53380 21913 53389 21947
rect 53389 21913 53423 21947
rect 53423 21913 53432 21947
rect 53380 21904 53432 21913
rect 53748 21836 53800 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 66314 21734 66366 21786
rect 66378 21734 66430 21786
rect 66442 21734 66494 21786
rect 66506 21734 66558 21786
rect 66570 21734 66622 21786
rect 12440 21675 12492 21684
rect 12440 21641 12449 21675
rect 12449 21641 12483 21675
rect 12483 21641 12492 21675
rect 12440 21632 12492 21641
rect 7380 21496 7432 21548
rect 7748 21564 7800 21616
rect 9680 21564 9732 21616
rect 10048 21564 10100 21616
rect 13452 21564 13504 21616
rect 29828 21632 29880 21684
rect 13912 21607 13964 21616
rect 13912 21573 13921 21607
rect 13921 21573 13955 21607
rect 13955 21573 13964 21607
rect 13912 21564 13964 21573
rect 30104 21607 30156 21616
rect 30104 21573 30113 21607
rect 30113 21573 30147 21607
rect 30147 21573 30156 21607
rect 30104 21564 30156 21573
rect 31116 21632 31168 21684
rect 38752 21632 38804 21684
rect 33416 21564 33468 21616
rect 29736 21539 29788 21548
rect 29736 21505 29745 21539
rect 29745 21505 29779 21539
rect 29779 21505 29788 21539
rect 29736 21496 29788 21505
rect 29920 21496 29972 21548
rect 30564 21496 30616 21548
rect 30656 21539 30708 21548
rect 30656 21505 30665 21539
rect 30665 21505 30699 21539
rect 30699 21505 30708 21539
rect 30656 21496 30708 21505
rect 14280 21428 14332 21480
rect 30472 21471 30524 21480
rect 30472 21437 30481 21471
rect 30481 21437 30515 21471
rect 30515 21437 30524 21471
rect 30472 21428 30524 21437
rect 7564 21360 7616 21412
rect 848 21292 900 21344
rect 8208 21292 8260 21344
rect 31024 21539 31076 21548
rect 31024 21505 31033 21539
rect 31033 21505 31067 21539
rect 31067 21505 31076 21539
rect 31024 21496 31076 21505
rect 31392 21539 31444 21548
rect 31392 21505 31401 21539
rect 31401 21505 31435 21539
rect 31435 21505 31444 21539
rect 31392 21496 31444 21505
rect 32128 21496 32180 21548
rect 37464 21539 37516 21548
rect 37464 21505 37473 21539
rect 37473 21505 37507 21539
rect 37507 21505 37516 21539
rect 37464 21496 37516 21505
rect 37648 21539 37700 21548
rect 37648 21505 37657 21539
rect 37657 21505 37691 21539
rect 37691 21505 37700 21539
rect 37648 21496 37700 21505
rect 34704 21428 34756 21480
rect 35440 21428 35492 21480
rect 30840 21292 30892 21344
rect 31392 21292 31444 21344
rect 35348 21360 35400 21412
rect 34336 21292 34388 21344
rect 37280 21335 37332 21344
rect 37280 21301 37289 21335
rect 37289 21301 37323 21335
rect 37323 21301 37332 21335
rect 37280 21292 37332 21301
rect 37556 21292 37608 21344
rect 37832 21292 37884 21344
rect 39488 21564 39540 21616
rect 39672 21564 39724 21616
rect 42156 21564 42208 21616
rect 49792 21632 49844 21684
rect 50068 21632 50120 21684
rect 50344 21632 50396 21684
rect 51356 21632 51408 21684
rect 53380 21632 53432 21684
rect 45376 21564 45428 21616
rect 46664 21564 46716 21616
rect 45100 21539 45152 21548
rect 45100 21505 45109 21539
rect 45109 21505 45143 21539
rect 45143 21505 45152 21539
rect 45100 21496 45152 21505
rect 45284 21539 45336 21548
rect 45284 21505 45293 21539
rect 45293 21505 45327 21539
rect 45327 21505 45336 21539
rect 45284 21496 45336 21505
rect 46940 21496 46992 21548
rect 47768 21539 47820 21548
rect 47768 21505 47777 21539
rect 47777 21505 47811 21539
rect 47811 21505 47820 21539
rect 47768 21496 47820 21505
rect 50804 21564 50856 21616
rect 52828 21564 52880 21616
rect 54484 21632 54536 21684
rect 53748 21564 53800 21616
rect 55312 21564 55364 21616
rect 49976 21539 50028 21548
rect 49976 21505 49985 21539
rect 49985 21505 50019 21539
rect 50019 21505 50028 21539
rect 49976 21496 50028 21505
rect 50068 21496 50120 21548
rect 39764 21471 39816 21480
rect 39764 21437 39773 21471
rect 39773 21437 39807 21471
rect 39807 21437 39816 21471
rect 39764 21428 39816 21437
rect 44916 21428 44968 21480
rect 40592 21360 40644 21412
rect 42616 21360 42668 21412
rect 46112 21360 46164 21412
rect 38660 21292 38712 21344
rect 46204 21335 46256 21344
rect 46204 21301 46213 21335
rect 46213 21301 46247 21335
rect 46247 21301 46256 21335
rect 46204 21292 46256 21301
rect 47400 21292 47452 21344
rect 48044 21335 48096 21344
rect 48044 21301 48053 21335
rect 48053 21301 48087 21335
rect 48087 21301 48096 21335
rect 48044 21292 48096 21301
rect 49700 21403 49752 21412
rect 49700 21369 49709 21403
rect 49709 21369 49743 21403
rect 49743 21369 49752 21403
rect 49700 21360 49752 21369
rect 50068 21360 50120 21412
rect 50436 21292 50488 21344
rect 50896 21539 50948 21548
rect 50896 21505 50905 21539
rect 50905 21505 50939 21539
rect 50939 21505 50948 21539
rect 50896 21496 50948 21505
rect 51172 21496 51224 21548
rect 54484 21496 54536 21548
rect 54852 21539 54904 21548
rect 54852 21505 54861 21539
rect 54861 21505 54895 21539
rect 54895 21505 54904 21539
rect 54852 21496 54904 21505
rect 54944 21539 54996 21548
rect 54944 21505 54953 21539
rect 54953 21505 54987 21539
rect 54987 21505 54996 21539
rect 54944 21496 54996 21505
rect 52184 21428 52236 21480
rect 56968 21539 57020 21548
rect 56968 21505 56977 21539
rect 56977 21505 57011 21539
rect 57011 21505 57020 21539
rect 56968 21496 57020 21505
rect 56232 21428 56284 21480
rect 56600 21428 56652 21480
rect 51632 21360 51684 21412
rect 52368 21360 52420 21412
rect 52920 21360 52972 21412
rect 55496 21360 55548 21412
rect 54208 21292 54260 21344
rect 55128 21335 55180 21344
rect 55128 21301 55137 21335
rect 55137 21301 55171 21335
rect 55171 21301 55180 21335
rect 55128 21292 55180 21301
rect 55220 21335 55272 21344
rect 55220 21301 55229 21335
rect 55229 21301 55263 21335
rect 55263 21301 55272 21335
rect 55220 21292 55272 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 7564 21131 7616 21140
rect 7564 21097 7573 21131
rect 7573 21097 7607 21131
rect 7607 21097 7616 21131
rect 7564 21088 7616 21097
rect 7932 21020 7984 21072
rect 7012 20995 7064 21004
rect 7012 20961 7021 20995
rect 7021 20961 7055 20995
rect 7055 20961 7064 20995
rect 7012 20952 7064 20961
rect 8208 20952 8260 21004
rect 7104 20927 7156 20936
rect 7104 20893 7113 20927
rect 7113 20893 7147 20927
rect 7147 20893 7156 20927
rect 7104 20884 7156 20893
rect 12992 20952 13044 21004
rect 11520 20927 11572 20936
rect 11520 20893 11529 20927
rect 11529 20893 11563 20927
rect 11563 20893 11572 20927
rect 11520 20884 11572 20893
rect 14924 21088 14976 21140
rect 31944 21088 31996 21140
rect 34520 21088 34572 21140
rect 34796 21088 34848 21140
rect 37372 21088 37424 21140
rect 39764 21088 39816 21140
rect 39856 21088 39908 21140
rect 38292 21020 38344 21072
rect 30472 20952 30524 21004
rect 29552 20927 29604 20936
rect 29552 20893 29561 20927
rect 29561 20893 29595 20927
rect 29595 20893 29604 20927
rect 29552 20884 29604 20893
rect 34520 20884 34572 20936
rect 37464 20952 37516 21004
rect 38568 20952 38620 21004
rect 39212 20995 39264 21004
rect 39212 20961 39221 20995
rect 39221 20961 39255 20995
rect 39255 20961 39264 20995
rect 39212 20952 39264 20961
rect 39488 21020 39540 21072
rect 41788 21088 41840 21140
rect 35992 20884 36044 20936
rect 38660 20884 38712 20936
rect 38936 20884 38988 20936
rect 39396 20927 39448 20936
rect 39396 20893 39405 20927
rect 39405 20893 39439 20927
rect 39439 20893 39448 20927
rect 39396 20884 39448 20893
rect 8576 20859 8628 20868
rect 8576 20825 8585 20859
rect 8585 20825 8619 20859
rect 8619 20825 8628 20859
rect 8576 20816 8628 20825
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 7472 20791 7524 20800
rect 7472 20757 7481 20791
rect 7481 20757 7515 20791
rect 7515 20757 7524 20791
rect 7472 20748 7524 20757
rect 7748 20748 7800 20800
rect 10600 20748 10652 20800
rect 10692 20748 10744 20800
rect 13544 20748 13596 20800
rect 30288 20816 30340 20868
rect 34612 20816 34664 20868
rect 31116 20748 31168 20800
rect 34980 20748 35032 20800
rect 37464 20859 37516 20868
rect 37464 20825 37473 20859
rect 37473 20825 37507 20859
rect 37507 20825 37516 20859
rect 37464 20816 37516 20825
rect 36176 20748 36228 20800
rect 36636 20748 36688 20800
rect 39672 20952 39724 21004
rect 45560 21020 45612 21072
rect 41972 20884 42024 20936
rect 42984 20884 43036 20936
rect 45376 20952 45428 21004
rect 46112 21088 46164 21140
rect 50804 21088 50856 21140
rect 53656 21088 53708 21140
rect 54944 21088 54996 21140
rect 56600 21131 56652 21140
rect 56600 21097 56609 21131
rect 56609 21097 56643 21131
rect 56643 21097 56652 21131
rect 56600 21088 56652 21097
rect 47124 21020 47176 21072
rect 50252 21020 50304 21072
rect 50896 21020 50948 21072
rect 51540 21020 51592 21072
rect 53012 21020 53064 21072
rect 48412 20952 48464 21004
rect 48596 20952 48648 21004
rect 40132 20859 40184 20868
rect 40132 20825 40141 20859
rect 40141 20825 40175 20859
rect 40175 20825 40184 20859
rect 40132 20816 40184 20825
rect 41144 20816 41196 20868
rect 42156 20859 42208 20868
rect 42156 20825 42165 20859
rect 42165 20825 42199 20859
rect 42199 20825 42208 20859
rect 42156 20816 42208 20825
rect 42524 20859 42576 20868
rect 42524 20825 42533 20859
rect 42533 20825 42567 20859
rect 42567 20825 42576 20859
rect 42524 20816 42576 20825
rect 42800 20816 42852 20868
rect 43352 20816 43404 20868
rect 44088 20859 44140 20868
rect 44088 20825 44097 20859
rect 44097 20825 44131 20859
rect 44131 20825 44140 20859
rect 44088 20816 44140 20825
rect 45192 20884 45244 20936
rect 45560 20884 45612 20936
rect 46756 20884 46808 20936
rect 50528 20952 50580 21004
rect 44548 20816 44600 20868
rect 44732 20816 44784 20868
rect 47124 20816 47176 20868
rect 41512 20748 41564 20800
rect 42708 20791 42760 20800
rect 42708 20757 42717 20791
rect 42717 20757 42751 20791
rect 42751 20757 42760 20791
rect 44272 20791 44324 20800
rect 42708 20748 42760 20757
rect 44272 20757 44281 20791
rect 44281 20757 44315 20791
rect 44315 20757 44324 20791
rect 45192 20791 45244 20800
rect 44272 20748 44324 20757
rect 45192 20757 45201 20791
rect 45201 20757 45235 20791
rect 45235 20757 45244 20791
rect 45192 20748 45244 20757
rect 48596 20791 48648 20800
rect 48596 20757 48605 20791
rect 48605 20757 48639 20791
rect 48639 20757 48648 20791
rect 48596 20748 48648 20757
rect 48872 20748 48924 20800
rect 49976 20884 50028 20936
rect 51632 20952 51684 21004
rect 52276 20995 52328 21004
rect 50896 20927 50948 20936
rect 50896 20893 50905 20927
rect 50905 20893 50939 20927
rect 50939 20893 50948 20927
rect 50896 20884 50948 20893
rect 52276 20961 52285 20995
rect 52285 20961 52319 20995
rect 52319 20961 52328 20995
rect 52276 20952 52328 20961
rect 52920 20927 52972 20936
rect 52920 20893 52929 20927
rect 52929 20893 52963 20927
rect 52963 20893 52972 20927
rect 52920 20884 52972 20893
rect 54208 20995 54260 21004
rect 54208 20961 54217 20995
rect 54217 20961 54251 20995
rect 54251 20961 54260 20995
rect 55128 21020 55180 21072
rect 54208 20952 54260 20961
rect 55220 20952 55272 21004
rect 52828 20816 52880 20868
rect 54576 20859 54628 20868
rect 54576 20825 54585 20859
rect 54585 20825 54619 20859
rect 54619 20825 54628 20859
rect 54576 20816 54628 20825
rect 50252 20748 50304 20800
rect 50804 20748 50856 20800
rect 53012 20748 53064 20800
rect 53104 20748 53156 20800
rect 55496 20816 55548 20868
rect 55128 20748 55180 20800
rect 55956 20748 56008 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 66314 20646 66366 20698
rect 66378 20646 66430 20698
rect 66442 20646 66494 20698
rect 66506 20646 66558 20698
rect 66570 20646 66622 20698
rect 7104 20544 7156 20596
rect 7932 20544 7984 20596
rect 7472 20476 7524 20528
rect 9680 20476 9732 20528
rect 34704 20587 34756 20596
rect 34704 20553 34713 20587
rect 34713 20553 34747 20587
rect 34747 20553 34756 20587
rect 34704 20544 34756 20553
rect 37280 20544 37332 20596
rect 37556 20544 37608 20596
rect 7380 20408 7432 20460
rect 7656 20408 7708 20460
rect 7840 20451 7892 20460
rect 7840 20417 7849 20451
rect 7849 20417 7883 20451
rect 7883 20417 7892 20451
rect 7840 20408 7892 20417
rect 8576 20340 8628 20392
rect 9496 20340 9548 20392
rect 10140 20476 10192 20528
rect 11520 20476 11572 20528
rect 12072 20476 12124 20528
rect 13544 20476 13596 20528
rect 19340 20476 19392 20528
rect 10140 20383 10192 20392
rect 10140 20349 10149 20383
rect 10149 20349 10183 20383
rect 10183 20349 10192 20383
rect 10140 20340 10192 20349
rect 10692 20340 10744 20392
rect 10968 20340 11020 20392
rect 9864 20247 9916 20256
rect 9864 20213 9873 20247
rect 9873 20213 9907 20247
rect 9907 20213 9916 20247
rect 9864 20204 9916 20213
rect 10416 20204 10468 20256
rect 14556 20204 14608 20256
rect 33416 20476 33468 20528
rect 27896 20451 27948 20460
rect 27896 20417 27905 20451
rect 27905 20417 27939 20451
rect 27939 20417 27948 20451
rect 27896 20408 27948 20417
rect 32128 20451 32180 20460
rect 32128 20417 32137 20451
rect 32137 20417 32171 20451
rect 32171 20417 32180 20451
rect 32128 20408 32180 20417
rect 33692 20408 33744 20460
rect 34980 20451 35032 20460
rect 34980 20417 34989 20451
rect 34989 20417 35023 20451
rect 35023 20417 35032 20451
rect 34980 20408 35032 20417
rect 35348 20408 35400 20460
rect 36636 20451 36688 20460
rect 36636 20417 36645 20451
rect 36645 20417 36679 20451
rect 36679 20417 36688 20451
rect 36636 20408 36688 20417
rect 37648 20476 37700 20528
rect 38200 20519 38252 20528
rect 38200 20485 38209 20519
rect 38209 20485 38243 20519
rect 38243 20485 38252 20519
rect 38200 20476 38252 20485
rect 39396 20544 39448 20596
rect 40132 20544 40184 20596
rect 41144 20544 41196 20596
rect 43904 20587 43956 20596
rect 43904 20553 43913 20587
rect 43913 20553 43947 20587
rect 43947 20553 43956 20587
rect 43904 20544 43956 20553
rect 44088 20476 44140 20528
rect 44364 20476 44416 20528
rect 46020 20476 46072 20528
rect 26608 20340 26660 20392
rect 29552 20340 29604 20392
rect 32404 20383 32456 20392
rect 32404 20349 32413 20383
rect 32413 20349 32447 20383
rect 32447 20349 32456 20383
rect 32404 20340 32456 20349
rect 34520 20340 34572 20392
rect 37464 20340 37516 20392
rect 39764 20408 39816 20460
rect 39856 20451 39908 20460
rect 39856 20417 39865 20451
rect 39865 20417 39899 20451
rect 39899 20417 39908 20451
rect 39856 20408 39908 20417
rect 40040 20408 40092 20460
rect 41604 20451 41656 20460
rect 41604 20417 41613 20451
rect 41613 20417 41647 20451
rect 41647 20417 41656 20451
rect 41604 20408 41656 20417
rect 31760 20272 31812 20324
rect 36176 20272 36228 20324
rect 25412 20204 25464 20256
rect 27896 20204 27948 20256
rect 33968 20247 34020 20256
rect 33968 20213 33977 20247
rect 33977 20213 34011 20247
rect 34011 20213 34020 20247
rect 33968 20204 34020 20213
rect 34428 20204 34480 20256
rect 36912 20247 36964 20256
rect 36912 20213 36921 20247
rect 36921 20213 36955 20247
rect 36955 20213 36964 20247
rect 36912 20204 36964 20213
rect 37004 20204 37056 20256
rect 41052 20340 41104 20392
rect 41512 20340 41564 20392
rect 39488 20247 39540 20256
rect 39488 20213 39497 20247
rect 39497 20213 39531 20247
rect 39531 20213 39540 20247
rect 39488 20204 39540 20213
rect 39856 20204 39908 20256
rect 39948 20204 40000 20256
rect 46664 20451 46716 20460
rect 46664 20417 46673 20451
rect 46673 20417 46707 20451
rect 46707 20417 46716 20451
rect 46664 20408 46716 20417
rect 47032 20544 47084 20596
rect 47216 20519 47268 20528
rect 47216 20485 47225 20519
rect 47225 20485 47259 20519
rect 47259 20485 47268 20519
rect 47216 20476 47268 20485
rect 47308 20408 47360 20460
rect 48688 20476 48740 20528
rect 52736 20544 52788 20596
rect 50804 20519 50856 20528
rect 50804 20485 50813 20519
rect 50813 20485 50847 20519
rect 50847 20485 50856 20519
rect 50804 20476 50856 20485
rect 53012 20519 53064 20528
rect 53012 20485 53021 20519
rect 53021 20485 53055 20519
rect 53055 20485 53064 20519
rect 53012 20476 53064 20485
rect 55220 20544 55272 20596
rect 55956 20587 56008 20596
rect 55956 20553 55965 20587
rect 55965 20553 55999 20587
rect 55999 20553 56008 20587
rect 55956 20544 56008 20553
rect 52736 20451 52788 20460
rect 52736 20417 52745 20451
rect 52745 20417 52779 20451
rect 52779 20417 52788 20451
rect 52736 20408 52788 20417
rect 54852 20451 54904 20460
rect 54852 20417 54861 20451
rect 54861 20417 54895 20451
rect 54895 20417 54904 20451
rect 54852 20408 54904 20417
rect 55128 20451 55180 20460
rect 55128 20417 55137 20451
rect 55137 20417 55171 20451
rect 55171 20417 55180 20451
rect 55128 20408 55180 20417
rect 55496 20408 55548 20460
rect 45192 20340 45244 20392
rect 47400 20340 47452 20392
rect 48412 20383 48464 20392
rect 48412 20349 48421 20383
rect 48421 20349 48455 20383
rect 48455 20349 48464 20383
rect 48412 20340 48464 20349
rect 52276 20383 52328 20392
rect 52276 20349 52285 20383
rect 52285 20349 52319 20383
rect 52319 20349 52328 20383
rect 52276 20340 52328 20349
rect 42524 20272 42576 20324
rect 44180 20272 44232 20324
rect 52184 20272 52236 20324
rect 54208 20272 54260 20324
rect 55128 20272 55180 20324
rect 44364 20204 44416 20256
rect 47860 20204 47912 20256
rect 48964 20204 49016 20256
rect 49516 20204 49568 20256
rect 53656 20204 53708 20256
rect 54944 20247 54996 20256
rect 54944 20213 54953 20247
rect 54953 20213 54987 20247
rect 54987 20213 54996 20247
rect 54944 20204 54996 20213
rect 55404 20247 55456 20256
rect 55404 20213 55413 20247
rect 55413 20213 55447 20247
rect 55447 20213 55456 20247
rect 55404 20204 55456 20213
rect 56048 20204 56100 20256
rect 56324 20204 56376 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 7380 19932 7432 19984
rect 7012 19864 7064 19916
rect 7656 20000 7708 20052
rect 7932 20000 7984 20052
rect 9864 20043 9916 20052
rect 9864 20009 9873 20043
rect 9873 20009 9907 20043
rect 9907 20009 9916 20043
rect 9864 20000 9916 20009
rect 10048 20043 10100 20052
rect 10048 20009 10057 20043
rect 10057 20009 10091 20043
rect 10091 20009 10100 20043
rect 10048 20000 10100 20009
rect 10140 20000 10192 20052
rect 7840 19864 7892 19916
rect 10968 19864 11020 19916
rect 27252 20000 27304 20052
rect 30104 20000 30156 20052
rect 31760 20043 31812 20052
rect 31760 20009 31769 20043
rect 31769 20009 31803 20043
rect 31803 20009 31812 20043
rect 31760 20000 31812 20009
rect 32404 20000 32456 20052
rect 34060 20043 34112 20052
rect 34060 20009 34069 20043
rect 34069 20009 34103 20043
rect 34103 20009 34112 20043
rect 34060 20000 34112 20009
rect 36268 20000 36320 20052
rect 36820 20000 36872 20052
rect 36912 20000 36964 20052
rect 39212 20000 39264 20052
rect 39948 20000 40000 20052
rect 47400 20000 47452 20052
rect 8208 19796 8260 19848
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 7840 19728 7892 19780
rect 12624 19796 12676 19848
rect 14280 19907 14332 19916
rect 14280 19873 14289 19907
rect 14289 19873 14323 19907
rect 14323 19873 14332 19907
rect 14280 19864 14332 19873
rect 14556 19907 14608 19916
rect 14556 19873 14565 19907
rect 14565 19873 14599 19907
rect 14599 19873 14608 19907
rect 14556 19864 14608 19873
rect 18512 19839 18564 19848
rect 18512 19805 18521 19839
rect 18521 19805 18555 19839
rect 18555 19805 18564 19839
rect 18512 19796 18564 19805
rect 24584 19796 24636 19848
rect 26608 19839 26660 19848
rect 26608 19805 26617 19839
rect 26617 19805 26651 19839
rect 26651 19805 26660 19839
rect 26608 19796 26660 19805
rect 26884 19796 26936 19848
rect 44548 19932 44600 19984
rect 46020 19932 46072 19984
rect 46848 19932 46900 19984
rect 48412 20000 48464 20052
rect 49148 20000 49200 20052
rect 48504 19975 48556 19984
rect 48504 19941 48513 19975
rect 48513 19941 48547 19975
rect 48547 19941 48556 19975
rect 50804 20000 50856 20052
rect 50896 20043 50948 20052
rect 50896 20009 50905 20043
rect 50905 20009 50939 20043
rect 50939 20009 50948 20043
rect 50896 20000 50948 20009
rect 51632 20000 51684 20052
rect 52828 20043 52880 20052
rect 52828 20009 52837 20043
rect 52837 20009 52871 20043
rect 52871 20009 52880 20043
rect 52828 20000 52880 20009
rect 54852 20000 54904 20052
rect 48504 19932 48556 19941
rect 33692 19864 33744 19916
rect 34428 19864 34480 19916
rect 10416 19771 10468 19780
rect 10416 19737 10425 19771
rect 10425 19737 10459 19771
rect 10459 19737 10468 19771
rect 10416 19728 10468 19737
rect 848 19660 900 19712
rect 7472 19703 7524 19712
rect 7472 19669 7481 19703
rect 7481 19669 7515 19703
rect 7515 19669 7524 19703
rect 7472 19660 7524 19669
rect 7748 19703 7800 19712
rect 7748 19669 7775 19703
rect 7775 19669 7800 19703
rect 7748 19660 7800 19669
rect 9680 19660 9732 19712
rect 30288 19728 30340 19780
rect 33968 19796 34020 19848
rect 34612 19796 34664 19848
rect 34888 19839 34940 19848
rect 34888 19805 34897 19839
rect 34897 19805 34931 19839
rect 34931 19805 34940 19839
rect 34888 19796 34940 19805
rect 35440 19864 35492 19916
rect 38936 19864 38988 19916
rect 39580 19864 39632 19916
rect 40684 19864 40736 19916
rect 35348 19796 35400 19848
rect 42984 19864 43036 19916
rect 42708 19796 42760 19848
rect 46664 19839 46716 19848
rect 46664 19805 46673 19839
rect 46673 19805 46707 19839
rect 46707 19805 46716 19839
rect 46664 19796 46716 19805
rect 46940 19796 46992 19848
rect 47768 19796 47820 19848
rect 50252 19864 50304 19916
rect 48780 19839 48832 19848
rect 48780 19805 48789 19839
rect 48789 19805 48823 19839
rect 48823 19805 48832 19839
rect 48780 19796 48832 19805
rect 48872 19839 48924 19848
rect 48872 19805 48881 19839
rect 48881 19805 48915 19839
rect 48915 19805 48924 19839
rect 48872 19796 48924 19805
rect 49056 19796 49108 19848
rect 49516 19796 49568 19848
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 14924 19660 14976 19712
rect 17868 19660 17920 19712
rect 17960 19703 18012 19712
rect 17960 19669 17969 19703
rect 17969 19669 18003 19703
rect 18003 19669 18012 19703
rect 17960 19660 18012 19669
rect 28816 19660 28868 19712
rect 30932 19660 30984 19712
rect 35164 19728 35216 19780
rect 37924 19728 37976 19780
rect 40868 19728 40920 19780
rect 44088 19728 44140 19780
rect 44548 19728 44600 19780
rect 47216 19771 47268 19780
rect 47216 19737 47225 19771
rect 47225 19737 47259 19771
rect 47259 19737 47268 19771
rect 47216 19728 47268 19737
rect 47400 19728 47452 19780
rect 35992 19660 36044 19712
rect 36728 19660 36780 19712
rect 36912 19660 36964 19712
rect 38200 19660 38252 19712
rect 38476 19660 38528 19712
rect 38844 19660 38896 19712
rect 44272 19660 44324 19712
rect 47032 19660 47084 19712
rect 48596 19728 48648 19780
rect 50436 19796 50488 19848
rect 50528 19839 50580 19848
rect 50528 19805 50537 19839
rect 50537 19805 50571 19839
rect 50571 19805 50580 19839
rect 50528 19796 50580 19805
rect 51080 19864 51132 19916
rect 50804 19796 50856 19848
rect 52184 19796 52236 19848
rect 52368 19796 52420 19848
rect 55404 19864 55456 19916
rect 57060 19907 57112 19916
rect 57060 19873 57069 19907
rect 57069 19873 57103 19907
rect 57103 19873 57112 19907
rect 57060 19864 57112 19873
rect 53104 19796 53156 19848
rect 54576 19728 54628 19780
rect 55220 19728 55272 19780
rect 50528 19660 50580 19712
rect 52368 19660 52420 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 66314 19558 66366 19610
rect 66378 19558 66430 19610
rect 66442 19558 66494 19610
rect 66506 19558 66558 19610
rect 66570 19558 66622 19610
rect 12072 19499 12124 19508
rect 12072 19465 12081 19499
rect 12081 19465 12115 19499
rect 12115 19465 12124 19499
rect 12072 19456 12124 19465
rect 15476 19456 15528 19508
rect 12992 19431 13044 19440
rect 12992 19397 13001 19431
rect 13001 19397 13035 19431
rect 13035 19397 13044 19431
rect 12992 19388 13044 19397
rect 14004 19388 14056 19440
rect 17960 19388 18012 19440
rect 24952 19388 25004 19440
rect 26608 19388 26660 19440
rect 7472 19320 7524 19372
rect 7748 19363 7800 19372
rect 7748 19329 7757 19363
rect 7757 19329 7791 19363
rect 7791 19329 7800 19363
rect 7748 19320 7800 19329
rect 7840 19363 7892 19372
rect 7840 19329 7849 19363
rect 7849 19329 7883 19363
rect 7883 19329 7892 19363
rect 7840 19320 7892 19329
rect 10600 19363 10652 19372
rect 10600 19329 10609 19363
rect 10609 19329 10643 19363
rect 10643 19329 10652 19363
rect 10600 19320 10652 19329
rect 9496 19252 9548 19304
rect 10048 19252 10100 19304
rect 12624 19320 12676 19372
rect 12716 19363 12768 19372
rect 12716 19329 12725 19363
rect 12725 19329 12759 19363
rect 12759 19329 12768 19363
rect 12716 19320 12768 19329
rect 16580 19320 16632 19372
rect 24584 19363 24636 19372
rect 24584 19329 24593 19363
rect 24593 19329 24627 19363
rect 24627 19329 24636 19363
rect 24584 19320 24636 19329
rect 26884 19320 26936 19372
rect 26976 19320 27028 19372
rect 27252 19363 27304 19372
rect 27252 19329 27261 19363
rect 27261 19329 27295 19363
rect 27295 19329 27304 19363
rect 27252 19320 27304 19329
rect 27344 19363 27396 19372
rect 27344 19329 27353 19363
rect 27353 19329 27387 19363
rect 27387 19329 27396 19363
rect 27344 19320 27396 19329
rect 27528 19363 27580 19372
rect 27528 19329 27537 19363
rect 27537 19329 27571 19363
rect 27571 19329 27580 19363
rect 27528 19320 27580 19329
rect 28816 19388 28868 19440
rect 30932 19388 30984 19440
rect 29644 19320 29696 19372
rect 35164 19388 35216 19440
rect 35440 19388 35492 19440
rect 19248 19252 19300 19304
rect 24860 19295 24912 19304
rect 24860 19261 24869 19295
rect 24869 19261 24903 19295
rect 24903 19261 24912 19295
rect 24860 19252 24912 19261
rect 28356 19295 28408 19304
rect 28356 19261 28365 19295
rect 28365 19261 28399 19295
rect 28399 19261 28408 19295
rect 28356 19252 28408 19261
rect 29828 19295 29880 19304
rect 29828 19261 29837 19295
rect 29837 19261 29871 19295
rect 29871 19261 29880 19295
rect 29828 19252 29880 19261
rect 31116 19252 31168 19304
rect 32956 19320 33008 19372
rect 34888 19320 34940 19372
rect 35348 19320 35400 19372
rect 35992 19320 36044 19372
rect 36176 19363 36228 19372
rect 36176 19329 36185 19363
rect 36185 19329 36219 19363
rect 36219 19329 36228 19363
rect 36176 19320 36228 19329
rect 36268 19363 36320 19372
rect 36268 19329 36277 19363
rect 36277 19329 36311 19363
rect 36311 19329 36320 19363
rect 36268 19320 36320 19329
rect 36728 19363 36780 19372
rect 36728 19329 36737 19363
rect 36737 19329 36771 19363
rect 36771 19329 36780 19363
rect 36728 19320 36780 19329
rect 36820 19363 36872 19372
rect 36820 19329 36829 19363
rect 36829 19329 36863 19363
rect 36863 19329 36872 19363
rect 36820 19320 36872 19329
rect 37188 19320 37240 19372
rect 37648 19456 37700 19508
rect 38016 19456 38068 19508
rect 38292 19456 38344 19508
rect 38384 19499 38436 19508
rect 38384 19465 38393 19499
rect 38393 19465 38427 19499
rect 38427 19465 38436 19499
rect 38384 19456 38436 19465
rect 38476 19456 38528 19508
rect 37924 19431 37976 19440
rect 37924 19397 37933 19431
rect 37933 19397 37967 19431
rect 37967 19397 37976 19431
rect 37924 19388 37976 19397
rect 40040 19499 40092 19508
rect 40040 19465 40049 19499
rect 40049 19465 40083 19499
rect 40083 19465 40092 19499
rect 40040 19456 40092 19465
rect 42616 19456 42668 19508
rect 43444 19456 43496 19508
rect 43628 19456 43680 19508
rect 44272 19499 44324 19508
rect 44272 19465 44281 19499
rect 44281 19465 44315 19499
rect 44315 19465 44324 19499
rect 44272 19456 44324 19465
rect 45192 19456 45244 19508
rect 47124 19456 47176 19508
rect 48504 19456 48556 19508
rect 32680 19252 32732 19304
rect 37372 19295 37424 19304
rect 7288 19116 7340 19168
rect 10232 19116 10284 19168
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 19064 19159 19116 19168
rect 19064 19125 19073 19159
rect 19073 19125 19107 19159
rect 19107 19125 19116 19159
rect 19064 19116 19116 19125
rect 26240 19116 26292 19168
rect 36544 19184 36596 19236
rect 37372 19261 37381 19295
rect 37381 19261 37415 19295
rect 37415 19261 37424 19295
rect 37372 19252 37424 19261
rect 38016 19363 38068 19372
rect 38016 19329 38030 19363
rect 38030 19329 38064 19363
rect 38064 19329 38068 19363
rect 38016 19320 38068 19329
rect 38936 19320 38988 19372
rect 39580 19320 39632 19372
rect 42340 19388 42392 19440
rect 42892 19388 42944 19440
rect 46848 19388 46900 19440
rect 47952 19431 48004 19440
rect 47952 19397 47961 19431
rect 47961 19397 47995 19431
rect 47995 19397 48004 19431
rect 47952 19388 48004 19397
rect 48688 19388 48740 19440
rect 56048 19388 56100 19440
rect 38292 19252 38344 19304
rect 38752 19252 38804 19304
rect 39028 19252 39080 19304
rect 39396 19252 39448 19304
rect 39856 19363 39908 19372
rect 39856 19329 39865 19363
rect 39865 19329 39899 19363
rect 39899 19329 39908 19363
rect 39856 19320 39908 19329
rect 40224 19320 40276 19372
rect 40316 19363 40368 19372
rect 40316 19329 40325 19363
rect 40325 19329 40359 19363
rect 40359 19329 40368 19363
rect 40316 19320 40368 19329
rect 40040 19252 40092 19304
rect 40684 19363 40736 19372
rect 40684 19329 40693 19363
rect 40693 19329 40727 19363
rect 40727 19329 40736 19363
rect 40684 19320 40736 19329
rect 40776 19320 40828 19372
rect 40960 19320 41012 19372
rect 39120 19184 39172 19236
rect 40316 19184 40368 19236
rect 32128 19159 32180 19168
rect 32128 19125 32137 19159
rect 32137 19125 32171 19159
rect 32171 19125 32180 19159
rect 32128 19116 32180 19125
rect 32864 19159 32916 19168
rect 32864 19125 32873 19159
rect 32873 19125 32907 19159
rect 32907 19125 32916 19159
rect 32864 19116 32916 19125
rect 32956 19116 33008 19168
rect 33416 19116 33468 19168
rect 34612 19116 34664 19168
rect 37188 19116 37240 19168
rect 38200 19159 38252 19168
rect 38200 19125 38209 19159
rect 38209 19125 38243 19159
rect 38243 19125 38252 19159
rect 38200 19116 38252 19125
rect 38384 19116 38436 19168
rect 39856 19116 39908 19168
rect 40132 19159 40184 19168
rect 40132 19125 40141 19159
rect 40141 19125 40175 19159
rect 40175 19125 40184 19159
rect 40132 19116 40184 19125
rect 41512 19116 41564 19168
rect 43720 19363 43772 19372
rect 43720 19329 43729 19363
rect 43729 19329 43763 19363
rect 43763 19329 43772 19363
rect 43720 19320 43772 19329
rect 44180 19363 44232 19372
rect 44180 19329 44189 19363
rect 44189 19329 44223 19363
rect 44223 19329 44232 19363
rect 44180 19320 44232 19329
rect 44548 19363 44600 19372
rect 44548 19329 44557 19363
rect 44557 19329 44591 19363
rect 44591 19329 44600 19363
rect 44548 19320 44600 19329
rect 47768 19363 47820 19372
rect 47768 19329 47777 19363
rect 47777 19329 47811 19363
rect 47811 19329 47820 19363
rect 47768 19320 47820 19329
rect 43260 19252 43312 19304
rect 44640 19295 44692 19304
rect 44640 19261 44649 19295
rect 44649 19261 44683 19295
rect 44683 19261 44692 19295
rect 44640 19252 44692 19261
rect 47124 19252 47176 19304
rect 49148 19320 49200 19372
rect 48228 19295 48280 19304
rect 48228 19261 48237 19295
rect 48237 19261 48271 19295
rect 48271 19261 48280 19295
rect 48228 19252 48280 19261
rect 48136 19184 48188 19236
rect 48872 19184 48924 19236
rect 43812 19116 43864 19168
rect 44824 19159 44876 19168
rect 44824 19125 44833 19159
rect 44833 19125 44867 19159
rect 44867 19125 44876 19159
rect 44824 19116 44876 19125
rect 51356 19116 51408 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 7840 18912 7892 18964
rect 9496 18776 9548 18828
rect 10784 18912 10836 18964
rect 18512 18912 18564 18964
rect 28356 18955 28408 18964
rect 28356 18921 28365 18955
rect 28365 18921 28399 18955
rect 28399 18921 28408 18955
rect 28356 18912 28408 18921
rect 29828 18955 29880 18964
rect 29828 18921 29837 18955
rect 29837 18921 29871 18955
rect 29871 18921 29880 18955
rect 29828 18912 29880 18921
rect 31116 18955 31168 18964
rect 31116 18921 31125 18955
rect 31125 18921 31159 18955
rect 31159 18921 31168 18955
rect 31116 18912 31168 18921
rect 32404 18912 32456 18964
rect 16488 18776 16540 18828
rect 17868 18776 17920 18828
rect 18604 18819 18656 18828
rect 18604 18785 18613 18819
rect 18613 18785 18647 18819
rect 18647 18785 18656 18819
rect 18604 18776 18656 18785
rect 19248 18819 19300 18828
rect 19248 18785 19257 18819
rect 19257 18785 19291 18819
rect 19291 18785 19300 18819
rect 19248 18776 19300 18785
rect 32864 18844 32916 18896
rect 35440 18912 35492 18964
rect 37280 18955 37332 18964
rect 37280 18921 37289 18955
rect 37289 18921 37323 18955
rect 37323 18921 37332 18955
rect 37280 18912 37332 18921
rect 37740 18912 37792 18964
rect 38108 18912 38160 18964
rect 38200 18955 38252 18964
rect 38200 18921 38209 18955
rect 38209 18921 38243 18955
rect 38243 18921 38252 18955
rect 38200 18912 38252 18921
rect 38752 18912 38804 18964
rect 33508 18844 33560 18896
rect 34520 18844 34572 18896
rect 9772 18708 9824 18760
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 10232 18751 10284 18760
rect 10232 18717 10241 18751
rect 10241 18717 10275 18751
rect 10275 18717 10284 18751
rect 10232 18708 10284 18717
rect 19064 18708 19116 18760
rect 23848 18708 23900 18760
rect 27344 18708 27396 18760
rect 7288 18683 7340 18692
rect 7288 18649 7297 18683
rect 7297 18649 7331 18683
rect 7331 18649 7340 18683
rect 7288 18640 7340 18649
rect 9312 18640 9364 18692
rect 14924 18640 14976 18692
rect 9864 18572 9916 18624
rect 10692 18572 10744 18624
rect 17960 18640 18012 18692
rect 18604 18640 18656 18692
rect 28080 18640 28132 18692
rect 28632 18640 28684 18692
rect 29184 18683 29236 18692
rect 29184 18649 29193 18683
rect 29193 18649 29227 18683
rect 29227 18649 29236 18683
rect 29184 18640 29236 18649
rect 29552 18751 29604 18760
rect 29552 18717 29561 18751
rect 29561 18717 29595 18751
rect 29595 18717 29604 18751
rect 29552 18708 29604 18717
rect 32128 18751 32180 18760
rect 32128 18717 32137 18751
rect 32137 18717 32171 18751
rect 32171 18717 32180 18751
rect 32128 18708 32180 18717
rect 32588 18708 32640 18760
rect 32772 18708 32824 18760
rect 34336 18819 34388 18828
rect 34336 18785 34345 18819
rect 34345 18785 34379 18819
rect 34379 18785 34388 18819
rect 34336 18776 34388 18785
rect 33324 18708 33376 18760
rect 33416 18751 33468 18760
rect 33416 18717 33425 18751
rect 33425 18717 33459 18751
rect 33459 18717 33468 18751
rect 33416 18708 33468 18717
rect 33508 18751 33560 18760
rect 33508 18717 33517 18751
rect 33517 18717 33551 18751
rect 33551 18717 33560 18751
rect 33508 18708 33560 18717
rect 33600 18751 33652 18760
rect 33600 18717 33633 18751
rect 33633 18717 33652 18751
rect 33600 18708 33652 18717
rect 33784 18708 33836 18760
rect 34060 18751 34112 18760
rect 34060 18717 34069 18751
rect 34069 18717 34103 18751
rect 34103 18717 34112 18751
rect 34060 18708 34112 18717
rect 18052 18572 18104 18624
rect 19800 18572 19852 18624
rect 21272 18572 21324 18624
rect 28356 18572 28408 18624
rect 29276 18615 29328 18624
rect 29276 18581 29285 18615
rect 29285 18581 29319 18615
rect 29319 18581 29328 18615
rect 29276 18572 29328 18581
rect 32036 18640 32088 18692
rect 32956 18640 33008 18692
rect 35348 18708 35400 18760
rect 36176 18751 36228 18760
rect 36176 18717 36185 18751
rect 36185 18717 36219 18751
rect 36219 18717 36228 18751
rect 36176 18708 36228 18717
rect 36912 18844 36964 18896
rect 38292 18844 38344 18896
rect 36452 18751 36504 18760
rect 36452 18717 36461 18751
rect 36461 18717 36495 18751
rect 36495 18717 36504 18751
rect 36452 18708 36504 18717
rect 36544 18751 36596 18760
rect 36544 18717 36553 18751
rect 36553 18717 36587 18751
rect 36587 18717 36596 18751
rect 36544 18708 36596 18717
rect 37004 18683 37056 18692
rect 30288 18572 30340 18624
rect 32496 18572 32548 18624
rect 37004 18649 37013 18683
rect 37013 18649 37047 18683
rect 37047 18649 37056 18683
rect 37004 18640 37056 18649
rect 37188 18708 37240 18760
rect 37464 18751 37516 18760
rect 37464 18717 37474 18751
rect 37474 18717 37508 18751
rect 37508 18717 37516 18751
rect 37464 18708 37516 18717
rect 37648 18751 37700 18760
rect 37648 18717 37657 18751
rect 37657 18717 37691 18751
rect 37691 18717 37700 18751
rect 37648 18708 37700 18717
rect 37832 18751 37884 18760
rect 37832 18717 37846 18751
rect 37846 18717 37880 18751
rect 37880 18717 37884 18751
rect 37832 18708 37884 18717
rect 40132 18955 40184 18964
rect 40132 18921 40141 18955
rect 40141 18921 40175 18955
rect 40175 18921 40184 18955
rect 40132 18912 40184 18921
rect 40500 18912 40552 18964
rect 41052 18955 41104 18964
rect 41052 18921 41061 18955
rect 41061 18921 41095 18955
rect 41095 18921 41104 18955
rect 41052 18912 41104 18921
rect 48228 18912 48280 18964
rect 52460 18912 52512 18964
rect 40684 18844 40736 18896
rect 47216 18844 47268 18896
rect 47308 18844 47360 18896
rect 49148 18844 49200 18896
rect 38844 18751 38896 18760
rect 38844 18717 38853 18751
rect 38853 18717 38887 18751
rect 38887 18717 38896 18751
rect 38844 18708 38896 18717
rect 39028 18751 39080 18760
rect 39028 18717 39035 18751
rect 39035 18717 39080 18751
rect 39028 18708 39080 18717
rect 39580 18751 39632 18760
rect 39580 18717 39589 18751
rect 39589 18717 39623 18751
rect 39623 18717 39632 18751
rect 39580 18708 39632 18717
rect 33876 18615 33928 18624
rect 33876 18581 33885 18615
rect 33885 18581 33919 18615
rect 33919 18581 33928 18615
rect 33876 18572 33928 18581
rect 36728 18572 36780 18624
rect 37280 18572 37332 18624
rect 37372 18572 37424 18624
rect 39212 18683 39264 18692
rect 39212 18649 39221 18683
rect 39221 18649 39255 18683
rect 39255 18649 39264 18683
rect 39212 18640 39264 18649
rect 39396 18572 39448 18624
rect 49700 18776 49752 18828
rect 51264 18776 51316 18828
rect 52092 18844 52144 18896
rect 55864 18912 55916 18964
rect 41052 18708 41104 18760
rect 40868 18683 40920 18692
rect 40868 18649 40877 18683
rect 40877 18649 40911 18683
rect 40911 18649 40920 18683
rect 40868 18640 40920 18649
rect 43260 18683 43312 18692
rect 43260 18649 43269 18683
rect 43269 18649 43303 18683
rect 43303 18649 43312 18683
rect 43260 18640 43312 18649
rect 43536 18751 43588 18760
rect 43536 18717 43545 18751
rect 43545 18717 43579 18751
rect 43579 18717 43588 18751
rect 43536 18708 43588 18717
rect 43720 18708 43772 18760
rect 45192 18708 45244 18760
rect 48412 18751 48464 18760
rect 48412 18717 48421 18751
rect 48421 18717 48455 18751
rect 48455 18717 48464 18751
rect 48412 18708 48464 18717
rect 49976 18751 50028 18760
rect 49976 18717 49985 18751
rect 49985 18717 50019 18751
rect 50019 18717 50028 18751
rect 49976 18708 50028 18717
rect 54484 18887 54536 18896
rect 54484 18853 54493 18887
rect 54493 18853 54527 18887
rect 54527 18853 54536 18887
rect 54484 18844 54536 18853
rect 54944 18844 54996 18896
rect 52276 18776 52328 18828
rect 56416 18776 56468 18828
rect 54392 18751 54444 18760
rect 54392 18717 54401 18751
rect 54401 18717 54435 18751
rect 54435 18717 54444 18751
rect 54392 18708 54444 18717
rect 54668 18751 54720 18760
rect 54668 18717 54677 18751
rect 54677 18717 54711 18751
rect 54711 18717 54720 18751
rect 54668 18708 54720 18717
rect 44640 18640 44692 18692
rect 50528 18683 50580 18692
rect 50528 18649 50537 18683
rect 50537 18649 50571 18683
rect 50571 18649 50580 18683
rect 50528 18640 50580 18649
rect 51908 18640 51960 18692
rect 54024 18683 54076 18692
rect 54024 18649 54033 18683
rect 54033 18649 54067 18683
rect 54067 18649 54076 18683
rect 54024 18640 54076 18649
rect 41696 18572 41748 18624
rect 42248 18572 42300 18624
rect 43168 18615 43220 18624
rect 43168 18581 43177 18615
rect 43177 18581 43211 18615
rect 43211 18581 43220 18615
rect 43168 18572 43220 18581
rect 43352 18572 43404 18624
rect 48136 18572 48188 18624
rect 48320 18572 48372 18624
rect 51448 18572 51500 18624
rect 53012 18572 53064 18624
rect 56140 18572 56192 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 66314 18470 66366 18522
rect 66378 18470 66430 18522
rect 66442 18470 66494 18522
rect 66506 18470 66558 18522
rect 66570 18470 66622 18522
rect 20352 18368 20404 18420
rect 23848 18411 23900 18420
rect 23848 18377 23857 18411
rect 23857 18377 23891 18411
rect 23891 18377 23900 18411
rect 23848 18368 23900 18377
rect 24860 18368 24912 18420
rect 9772 18232 9824 18284
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 17868 18232 17920 18284
rect 19248 18232 19300 18284
rect 20076 18275 20128 18284
rect 20076 18241 20085 18275
rect 20085 18241 20119 18275
rect 20119 18241 20128 18275
rect 20076 18232 20128 18241
rect 20444 18232 20496 18284
rect 20536 18232 20588 18284
rect 21272 18275 21324 18284
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 21272 18232 21324 18241
rect 27528 18368 27580 18420
rect 28356 18411 28408 18420
rect 28356 18377 28365 18411
rect 28365 18377 28399 18411
rect 28399 18377 28408 18411
rect 28356 18368 28408 18377
rect 28632 18368 28684 18420
rect 30748 18368 30800 18420
rect 33324 18368 33376 18420
rect 34796 18368 34848 18420
rect 34888 18368 34940 18420
rect 14280 18207 14332 18216
rect 14280 18173 14289 18207
rect 14289 18173 14323 18207
rect 14323 18173 14332 18207
rect 14280 18164 14332 18173
rect 21456 18164 21508 18216
rect 22100 18207 22152 18216
rect 22100 18173 22109 18207
rect 22109 18173 22143 18207
rect 22143 18173 22152 18207
rect 22100 18164 22152 18173
rect 18604 18139 18656 18148
rect 18604 18105 18613 18139
rect 18613 18105 18647 18139
rect 18647 18105 18656 18139
rect 18604 18096 18656 18105
rect 24492 18275 24544 18284
rect 24492 18241 24501 18275
rect 24501 18241 24535 18275
rect 24535 18241 24544 18275
rect 24492 18232 24544 18241
rect 25596 18232 25648 18284
rect 25688 18275 25740 18284
rect 25688 18241 25697 18275
rect 25697 18241 25731 18275
rect 25731 18241 25740 18275
rect 25688 18232 25740 18241
rect 27436 18300 27488 18352
rect 29276 18343 29328 18352
rect 25964 18275 26016 18284
rect 25964 18241 25973 18275
rect 25973 18241 26007 18275
rect 26007 18241 26016 18275
rect 25964 18232 26016 18241
rect 27804 18232 27856 18284
rect 28080 18275 28132 18284
rect 28080 18241 28089 18275
rect 28089 18241 28123 18275
rect 28123 18241 28132 18275
rect 28080 18232 28132 18241
rect 28172 18275 28224 18284
rect 28172 18241 28181 18275
rect 28181 18241 28215 18275
rect 28215 18241 28224 18275
rect 28172 18232 28224 18241
rect 26332 18207 26384 18216
rect 26332 18173 26341 18207
rect 26341 18173 26375 18207
rect 26375 18173 26384 18207
rect 26332 18164 26384 18173
rect 26516 18207 26568 18216
rect 26516 18173 26525 18207
rect 26525 18173 26559 18207
rect 26559 18173 26568 18207
rect 26516 18164 26568 18173
rect 27620 18164 27672 18216
rect 28632 18275 28684 18284
rect 28632 18241 28641 18275
rect 28641 18241 28675 18275
rect 28675 18241 28684 18275
rect 28632 18232 28684 18241
rect 29276 18309 29285 18343
rect 29285 18309 29319 18343
rect 29319 18309 29328 18343
rect 29276 18300 29328 18309
rect 32220 18300 32272 18352
rect 30748 18232 30800 18284
rect 32036 18232 32088 18284
rect 33784 18300 33836 18352
rect 33876 18343 33928 18352
rect 33876 18309 33885 18343
rect 33885 18309 33919 18343
rect 33919 18309 33928 18343
rect 33876 18300 33928 18309
rect 35440 18300 35492 18352
rect 36176 18368 36228 18420
rect 36452 18368 36504 18420
rect 36728 18368 36780 18420
rect 37280 18368 37332 18420
rect 37556 18368 37608 18420
rect 39396 18368 39448 18420
rect 32496 18232 32548 18284
rect 32680 18275 32732 18284
rect 32680 18241 32689 18275
rect 32689 18241 32723 18275
rect 32723 18241 32732 18275
rect 32680 18232 32732 18241
rect 35532 18232 35584 18284
rect 29460 18207 29512 18216
rect 29460 18173 29469 18207
rect 29469 18173 29503 18207
rect 29503 18173 29512 18207
rect 29460 18164 29512 18173
rect 33876 18164 33928 18216
rect 34888 18164 34940 18216
rect 36084 18275 36136 18284
rect 36084 18241 36093 18275
rect 36093 18241 36127 18275
rect 36127 18241 36136 18275
rect 36084 18232 36136 18241
rect 36268 18164 36320 18216
rect 36452 18164 36504 18216
rect 24860 18096 24912 18148
rect 24952 18096 25004 18148
rect 25504 18096 25556 18148
rect 27344 18096 27396 18148
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 13268 18028 13320 18080
rect 19984 18028 20036 18080
rect 23020 18028 23072 18080
rect 25688 18028 25740 18080
rect 28264 18028 28316 18080
rect 30656 18028 30708 18080
rect 30748 18071 30800 18080
rect 30748 18037 30757 18071
rect 30757 18037 30791 18071
rect 30791 18037 30800 18071
rect 30748 18028 30800 18037
rect 32128 18071 32180 18080
rect 32128 18037 32137 18071
rect 32137 18037 32171 18071
rect 32171 18037 32180 18071
rect 32128 18028 32180 18037
rect 32404 18028 32456 18080
rect 33416 18028 33468 18080
rect 34520 18028 34572 18080
rect 36820 18232 36872 18284
rect 37832 18300 37884 18352
rect 38108 18343 38160 18352
rect 38108 18309 38117 18343
rect 38117 18309 38151 18343
rect 38151 18309 38160 18343
rect 38108 18300 38160 18309
rect 41512 18300 41564 18352
rect 42984 18368 43036 18420
rect 43352 18300 43404 18352
rect 44364 18300 44416 18352
rect 46848 18368 46900 18420
rect 37004 18164 37056 18216
rect 37740 18232 37792 18284
rect 40684 18232 40736 18284
rect 42708 18232 42760 18284
rect 49976 18368 50028 18420
rect 48320 18343 48372 18352
rect 48320 18309 48329 18343
rect 48329 18309 48363 18343
rect 48363 18309 48372 18343
rect 48320 18300 48372 18309
rect 37464 18164 37516 18216
rect 40224 18164 40276 18216
rect 37372 18096 37424 18148
rect 38292 18096 38344 18148
rect 39304 18096 39356 18148
rect 35348 18071 35400 18080
rect 35348 18037 35357 18071
rect 35357 18037 35391 18071
rect 35391 18037 35400 18071
rect 35348 18028 35400 18037
rect 36084 18028 36136 18080
rect 38384 18028 38436 18080
rect 38752 18028 38804 18080
rect 42248 18207 42300 18216
rect 42248 18173 42257 18207
rect 42257 18173 42291 18207
rect 42291 18173 42300 18207
rect 42800 18207 42852 18216
rect 42248 18164 42300 18173
rect 42800 18173 42809 18207
rect 42809 18173 42843 18207
rect 42843 18173 42852 18207
rect 42800 18164 42852 18173
rect 43076 18207 43128 18216
rect 43076 18173 43085 18207
rect 43085 18173 43119 18207
rect 43119 18173 43128 18207
rect 43076 18164 43128 18173
rect 45560 18207 45612 18216
rect 45560 18173 45569 18207
rect 45569 18173 45603 18207
rect 45603 18173 45612 18207
rect 45560 18164 45612 18173
rect 48320 18164 48372 18216
rect 50252 18275 50304 18284
rect 50252 18241 50261 18275
rect 50261 18241 50295 18275
rect 50295 18241 50304 18275
rect 50252 18232 50304 18241
rect 50528 18368 50580 18420
rect 54024 18368 54076 18420
rect 51448 18300 51500 18352
rect 54116 18300 54168 18352
rect 55864 18300 55916 18352
rect 56140 18343 56192 18352
rect 56140 18309 56149 18343
rect 56149 18309 56183 18343
rect 56183 18309 56192 18343
rect 56140 18300 56192 18309
rect 50436 18232 50488 18284
rect 50804 18232 50856 18284
rect 42892 18028 42944 18080
rect 44548 18071 44600 18080
rect 44548 18037 44557 18071
rect 44557 18037 44591 18071
rect 44591 18037 44600 18071
rect 44548 18028 44600 18037
rect 47032 18071 47084 18080
rect 47032 18037 47041 18071
rect 47041 18037 47075 18071
rect 47075 18037 47084 18071
rect 47032 18028 47084 18037
rect 50620 18164 50672 18216
rect 52460 18275 52512 18284
rect 52460 18241 52469 18275
rect 52469 18241 52503 18275
rect 52503 18241 52512 18275
rect 52460 18232 52512 18241
rect 53012 18275 53064 18284
rect 53012 18241 53021 18275
rect 53021 18241 53055 18275
rect 53055 18241 53064 18275
rect 53012 18232 53064 18241
rect 54024 18275 54076 18284
rect 54024 18241 54033 18275
rect 54033 18241 54067 18275
rect 54067 18241 54076 18275
rect 54024 18232 54076 18241
rect 56416 18275 56468 18284
rect 56416 18241 56425 18275
rect 56425 18241 56459 18275
rect 56459 18241 56468 18275
rect 56416 18232 56468 18241
rect 51908 18096 51960 18148
rect 51356 18071 51408 18080
rect 51356 18037 51365 18071
rect 51365 18037 51399 18071
rect 51399 18037 51408 18071
rect 54484 18164 54536 18216
rect 51356 18028 51408 18037
rect 53932 18028 53984 18080
rect 54392 18028 54444 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 16212 17799 16264 17808
rect 16212 17765 16221 17799
rect 16221 17765 16255 17799
rect 16255 17765 16264 17799
rect 16212 17756 16264 17765
rect 10692 17731 10744 17740
rect 10692 17697 10701 17731
rect 10701 17697 10735 17731
rect 10735 17697 10744 17731
rect 10692 17688 10744 17697
rect 13268 17731 13320 17740
rect 13268 17697 13277 17731
rect 13277 17697 13311 17731
rect 13311 17697 13320 17731
rect 13268 17688 13320 17697
rect 15108 17688 15160 17740
rect 9496 17620 9548 17672
rect 12716 17620 12768 17672
rect 16488 17688 16540 17740
rect 22100 17824 22152 17876
rect 26516 17824 26568 17876
rect 29736 17824 29788 17876
rect 30748 17824 30800 17876
rect 31392 17824 31444 17876
rect 32680 17824 32732 17876
rect 32956 17824 33008 17876
rect 33048 17824 33100 17876
rect 19340 17799 19392 17808
rect 17500 17663 17552 17672
rect 17500 17629 17509 17663
rect 17509 17629 17543 17663
rect 17543 17629 17552 17663
rect 19340 17765 19349 17799
rect 19349 17765 19383 17799
rect 19383 17765 19392 17799
rect 19340 17756 19392 17765
rect 20536 17799 20588 17808
rect 20536 17765 20545 17799
rect 20545 17765 20579 17799
rect 20579 17765 20588 17799
rect 20536 17756 20588 17765
rect 18420 17688 18472 17740
rect 19984 17688 20036 17740
rect 21456 17799 21508 17808
rect 21456 17765 21465 17799
rect 21465 17765 21499 17799
rect 21499 17765 21508 17799
rect 21456 17756 21508 17765
rect 25596 17756 25648 17808
rect 17500 17620 17552 17629
rect 11152 17552 11204 17604
rect 14188 17552 14240 17604
rect 14740 17595 14792 17604
rect 14740 17561 14749 17595
rect 14749 17561 14783 17595
rect 14783 17561 14792 17595
rect 14740 17552 14792 17561
rect 18144 17552 18196 17604
rect 18604 17620 18656 17672
rect 20076 17620 20128 17672
rect 20628 17620 20680 17672
rect 20444 17552 20496 17604
rect 22100 17620 22152 17672
rect 25964 17663 26016 17672
rect 25964 17629 25972 17663
rect 25972 17629 26006 17663
rect 26006 17629 26016 17663
rect 25964 17620 26016 17629
rect 26240 17620 26292 17672
rect 27252 17663 27304 17672
rect 27252 17629 27261 17663
rect 27261 17629 27295 17663
rect 27295 17629 27304 17663
rect 27252 17620 27304 17629
rect 12440 17484 12492 17536
rect 14924 17484 14976 17536
rect 15568 17484 15620 17536
rect 20996 17527 21048 17536
rect 20996 17493 21005 17527
rect 21005 17493 21039 17527
rect 21039 17493 21048 17527
rect 26976 17552 27028 17604
rect 27436 17620 27488 17672
rect 31024 17756 31076 17808
rect 27712 17552 27764 17604
rect 28540 17688 28592 17740
rect 28264 17663 28316 17672
rect 28264 17629 28273 17663
rect 28273 17629 28307 17663
rect 28307 17629 28316 17663
rect 28264 17620 28316 17629
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 30656 17688 30708 17740
rect 31116 17731 31168 17740
rect 31116 17697 31125 17731
rect 31125 17697 31159 17731
rect 31159 17697 31168 17731
rect 31116 17688 31168 17697
rect 32128 17688 32180 17740
rect 28908 17552 28960 17604
rect 20996 17484 21048 17493
rect 27252 17484 27304 17536
rect 30932 17620 30984 17672
rect 31024 17552 31076 17604
rect 31116 17552 31168 17604
rect 29828 17484 29880 17536
rect 30748 17484 30800 17536
rect 33140 17527 33192 17536
rect 33140 17493 33149 17527
rect 33149 17493 33183 17527
rect 33183 17493 33192 17527
rect 33140 17484 33192 17493
rect 33324 17484 33376 17536
rect 33784 17867 33836 17876
rect 33784 17833 33793 17867
rect 33793 17833 33827 17867
rect 33827 17833 33836 17867
rect 33784 17824 33836 17833
rect 34428 17824 34480 17876
rect 36452 17799 36504 17808
rect 36452 17765 36461 17799
rect 36461 17765 36495 17799
rect 36495 17765 36504 17799
rect 36452 17756 36504 17765
rect 33600 17620 33652 17672
rect 35348 17688 35400 17740
rect 35440 17620 35492 17672
rect 37556 17824 37608 17876
rect 38844 17824 38896 17876
rect 40868 17824 40920 17876
rect 41328 17824 41380 17876
rect 42248 17824 42300 17876
rect 43444 17824 43496 17876
rect 45560 17824 45612 17876
rect 37280 17756 37332 17808
rect 38476 17756 38528 17808
rect 39396 17756 39448 17808
rect 37464 17688 37516 17740
rect 38568 17688 38620 17740
rect 40868 17688 40920 17740
rect 41328 17731 41380 17740
rect 41328 17697 41337 17731
rect 41337 17697 41371 17731
rect 41371 17697 41380 17731
rect 41328 17688 41380 17697
rect 36544 17552 36596 17604
rect 33784 17484 33836 17536
rect 34520 17484 34572 17536
rect 35348 17484 35400 17536
rect 35532 17484 35584 17536
rect 36360 17484 36412 17536
rect 37372 17620 37424 17672
rect 39028 17620 39080 17672
rect 40040 17663 40092 17672
rect 40040 17629 40047 17663
rect 40047 17629 40092 17663
rect 38200 17595 38252 17604
rect 38200 17561 38209 17595
rect 38209 17561 38243 17595
rect 38243 17561 38252 17595
rect 38200 17552 38252 17561
rect 39672 17552 39724 17604
rect 37280 17527 37332 17536
rect 37280 17493 37289 17527
rect 37289 17493 37323 17527
rect 37323 17493 37332 17527
rect 37280 17484 37332 17493
rect 37372 17484 37424 17536
rect 39028 17484 39080 17536
rect 40040 17620 40092 17629
rect 40224 17663 40276 17672
rect 40224 17629 40233 17663
rect 40233 17629 40267 17663
rect 40267 17629 40276 17663
rect 40224 17620 40276 17629
rect 40316 17663 40368 17672
rect 40316 17629 40330 17663
rect 40330 17629 40364 17663
rect 40364 17629 40368 17663
rect 40316 17620 40368 17629
rect 40960 17620 41012 17672
rect 42432 17731 42484 17740
rect 42432 17697 42441 17731
rect 42441 17697 42475 17731
rect 42475 17697 42484 17731
rect 42432 17688 42484 17697
rect 42524 17688 42576 17740
rect 40592 17595 40644 17604
rect 40592 17561 40601 17595
rect 40601 17561 40635 17595
rect 40635 17561 40644 17595
rect 40592 17552 40644 17561
rect 41420 17552 41472 17604
rect 42616 17663 42668 17672
rect 42616 17629 42625 17663
rect 42625 17629 42659 17663
rect 42659 17629 42668 17663
rect 42616 17620 42668 17629
rect 42892 17731 42944 17740
rect 42892 17697 42901 17731
rect 42901 17697 42935 17731
rect 42935 17697 42944 17731
rect 42892 17688 42944 17697
rect 44548 17688 44600 17740
rect 46296 17799 46348 17808
rect 46296 17765 46305 17799
rect 46305 17765 46339 17799
rect 46339 17765 46348 17799
rect 46296 17756 46348 17765
rect 47308 17756 47360 17808
rect 47584 17824 47636 17876
rect 47860 17824 47912 17876
rect 48412 17867 48464 17876
rect 48412 17833 48421 17867
rect 48421 17833 48455 17867
rect 48455 17833 48464 17867
rect 48412 17824 48464 17833
rect 50804 17824 50856 17876
rect 51080 17824 51132 17876
rect 52552 17824 52604 17876
rect 53196 17824 53248 17876
rect 54024 17824 54076 17876
rect 54668 17824 54720 17876
rect 48780 17756 48832 17808
rect 50252 17756 50304 17808
rect 47032 17688 47084 17740
rect 47952 17688 48004 17740
rect 43168 17663 43220 17672
rect 43168 17629 43177 17663
rect 43177 17629 43211 17663
rect 43211 17629 43220 17663
rect 43168 17620 43220 17629
rect 43352 17663 43404 17672
rect 43352 17629 43361 17663
rect 43361 17629 43395 17663
rect 43395 17629 43404 17663
rect 43352 17620 43404 17629
rect 46020 17663 46072 17672
rect 46020 17629 46029 17663
rect 46029 17629 46063 17663
rect 46063 17629 46072 17663
rect 46020 17620 46072 17629
rect 46112 17663 46164 17672
rect 46112 17629 46121 17663
rect 46121 17629 46155 17663
rect 46155 17629 46164 17663
rect 46112 17620 46164 17629
rect 47768 17663 47820 17672
rect 47768 17629 47777 17663
rect 47777 17629 47811 17663
rect 47811 17629 47820 17663
rect 47768 17620 47820 17629
rect 47860 17663 47912 17672
rect 47860 17629 47870 17663
rect 47870 17629 47904 17663
rect 47904 17629 47912 17663
rect 47860 17620 47912 17629
rect 48136 17663 48188 17672
rect 48136 17629 48145 17663
rect 48145 17629 48179 17663
rect 48179 17629 48188 17663
rect 48136 17620 48188 17629
rect 49516 17688 49568 17740
rect 50988 17688 51040 17740
rect 51908 17620 51960 17672
rect 52460 17688 52512 17740
rect 41328 17484 41380 17536
rect 43168 17484 43220 17536
rect 43444 17484 43496 17536
rect 43720 17484 43772 17536
rect 45928 17552 45980 17604
rect 50344 17552 50396 17604
rect 51080 17552 51132 17604
rect 53196 17663 53248 17672
rect 54116 17756 54168 17808
rect 53196 17629 53210 17663
rect 53210 17629 53244 17663
rect 53244 17629 53248 17663
rect 53196 17620 53248 17629
rect 54116 17620 54168 17672
rect 54576 17620 54628 17672
rect 46204 17484 46256 17536
rect 47584 17527 47636 17536
rect 47584 17493 47593 17527
rect 47593 17493 47627 17527
rect 47627 17493 47636 17527
rect 47584 17484 47636 17493
rect 47768 17484 47820 17536
rect 50252 17484 50304 17536
rect 53012 17595 53064 17604
rect 53012 17561 53021 17595
rect 53021 17561 53055 17595
rect 53055 17561 53064 17595
rect 53012 17552 53064 17561
rect 55036 17552 55088 17604
rect 53932 17484 53984 17536
rect 54116 17484 54168 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 66314 17382 66366 17434
rect 66378 17382 66430 17434
rect 66442 17382 66494 17434
rect 66506 17382 66558 17434
rect 66570 17382 66622 17434
rect 9496 17280 9548 17332
rect 9680 17212 9732 17264
rect 14740 17280 14792 17332
rect 15476 17323 15528 17332
rect 15476 17289 15485 17323
rect 15485 17289 15519 17323
rect 15519 17289 15528 17323
rect 15476 17280 15528 17289
rect 15568 17323 15620 17332
rect 15568 17289 15577 17323
rect 15577 17289 15611 17323
rect 15611 17289 15620 17323
rect 15568 17280 15620 17289
rect 9496 17187 9548 17196
rect 9496 17153 9505 17187
rect 9505 17153 9539 17187
rect 9539 17153 9548 17187
rect 9496 17144 9548 17153
rect 9312 17076 9364 17128
rect 10784 17076 10836 17128
rect 11152 17144 11204 17196
rect 12716 17212 12768 17264
rect 14004 17212 14056 17264
rect 14188 17187 14240 17196
rect 14188 17153 14197 17187
rect 14197 17153 14231 17187
rect 14231 17153 14240 17187
rect 20536 17280 20588 17332
rect 29184 17280 29236 17332
rect 29736 17280 29788 17332
rect 17960 17212 18012 17264
rect 14188 17144 14240 17153
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 14280 17119 14332 17128
rect 14280 17085 14289 17119
rect 14289 17085 14323 17119
rect 14323 17085 14332 17119
rect 14280 17076 14332 17085
rect 15016 17076 15068 17128
rect 16212 17119 16264 17128
rect 16212 17085 16221 17119
rect 16221 17085 16255 17119
rect 16255 17085 16264 17119
rect 16212 17076 16264 17085
rect 16488 17076 16540 17128
rect 17316 17119 17368 17128
rect 17316 17085 17325 17119
rect 17325 17085 17359 17119
rect 17359 17085 17368 17119
rect 17316 17076 17368 17085
rect 18328 17076 18380 17128
rect 23112 17187 23164 17196
rect 23112 17153 23121 17187
rect 23121 17153 23155 17187
rect 23155 17153 23164 17187
rect 23112 17144 23164 17153
rect 23296 17187 23348 17196
rect 23296 17153 23305 17187
rect 23305 17153 23339 17187
rect 23339 17153 23348 17187
rect 23296 17144 23348 17153
rect 24032 17144 24084 17196
rect 27804 17187 27856 17196
rect 27804 17153 27813 17187
rect 27813 17153 27847 17187
rect 27847 17153 27856 17187
rect 27804 17144 27856 17153
rect 28356 17212 28408 17264
rect 28816 17212 28868 17264
rect 28264 17187 28316 17196
rect 28264 17153 28273 17187
rect 28273 17153 28307 17187
rect 28307 17153 28316 17187
rect 28264 17144 28316 17153
rect 18972 17076 19024 17128
rect 12164 16940 12216 16992
rect 14004 16940 14056 16992
rect 14464 16983 14516 16992
rect 14464 16949 14473 16983
rect 14473 16949 14507 16983
rect 14507 16949 14516 16983
rect 14464 16940 14516 16949
rect 17040 16940 17092 16992
rect 19984 17008 20036 17060
rect 20076 16940 20128 16992
rect 20444 17076 20496 17128
rect 27436 17076 27488 17128
rect 28540 17187 28592 17196
rect 28540 17153 28549 17187
rect 28549 17153 28583 17187
rect 28583 17153 28592 17187
rect 28540 17144 28592 17153
rect 28908 17144 28960 17196
rect 29368 17144 29420 17196
rect 29828 17144 29880 17196
rect 30012 17187 30064 17196
rect 30012 17153 30021 17187
rect 30021 17153 30055 17187
rect 30055 17153 30064 17187
rect 30012 17144 30064 17153
rect 30196 17255 30248 17264
rect 30196 17221 30205 17255
rect 30205 17221 30239 17255
rect 30239 17221 30248 17255
rect 30196 17212 30248 17221
rect 30748 17280 30800 17332
rect 31024 17323 31076 17332
rect 31024 17289 31033 17323
rect 31033 17289 31067 17323
rect 31067 17289 31076 17323
rect 31024 17280 31076 17289
rect 32036 17280 32088 17332
rect 30656 17144 30708 17196
rect 33140 17280 33192 17332
rect 36452 17212 36504 17264
rect 29184 17076 29236 17128
rect 29736 17119 29788 17128
rect 29736 17085 29745 17119
rect 29745 17085 29779 17119
rect 29779 17085 29788 17119
rect 29736 17076 29788 17085
rect 31024 17119 31076 17128
rect 31024 17085 31033 17119
rect 31033 17085 31067 17119
rect 31067 17085 31076 17119
rect 31024 17076 31076 17085
rect 20536 17051 20588 17060
rect 20536 17017 20545 17051
rect 20545 17017 20579 17051
rect 20579 17017 20588 17051
rect 20536 17008 20588 17017
rect 20444 16940 20496 16992
rect 20628 16983 20680 16992
rect 20628 16949 20637 16983
rect 20637 16949 20671 16983
rect 20671 16949 20680 16983
rect 20628 16940 20680 16949
rect 20812 16983 20864 16992
rect 20812 16949 20821 16983
rect 20821 16949 20855 16983
rect 20855 16949 20864 16983
rect 20812 16940 20864 16949
rect 28172 17008 28224 17060
rect 28816 17008 28868 17060
rect 29092 17051 29144 17060
rect 27712 16940 27764 16992
rect 28632 16940 28684 16992
rect 29092 17017 29101 17051
rect 29101 17017 29135 17051
rect 29135 17017 29144 17051
rect 29092 17008 29144 17017
rect 29184 16940 29236 16992
rect 32588 17187 32640 17196
rect 32588 17153 32597 17187
rect 32597 17153 32631 17187
rect 32631 17153 32640 17187
rect 32588 17144 32640 17153
rect 32864 17144 32916 17196
rect 32956 17187 33008 17196
rect 32956 17153 32965 17187
rect 32965 17153 32999 17187
rect 32999 17153 33008 17187
rect 32956 17144 33008 17153
rect 33232 17144 33284 17196
rect 33600 17187 33652 17196
rect 33600 17153 33609 17187
rect 33609 17153 33643 17187
rect 33643 17153 33652 17187
rect 33600 17144 33652 17153
rect 34060 17144 34112 17196
rect 34520 17187 34572 17196
rect 34520 17153 34529 17187
rect 34529 17153 34563 17187
rect 34563 17153 34572 17187
rect 34520 17144 34572 17153
rect 34796 17187 34848 17196
rect 34796 17153 34805 17187
rect 34805 17153 34839 17187
rect 34839 17153 34848 17187
rect 34796 17144 34848 17153
rect 33416 17119 33468 17128
rect 33416 17085 33425 17119
rect 33425 17085 33459 17119
rect 33459 17085 33468 17119
rect 33416 17076 33468 17085
rect 34336 17076 34388 17128
rect 31760 16983 31812 16992
rect 31760 16949 31769 16983
rect 31769 16949 31803 16983
rect 31803 16949 31812 16983
rect 31760 16940 31812 16949
rect 32404 16983 32456 16992
rect 32404 16949 32413 16983
rect 32413 16949 32447 16983
rect 32447 16949 32456 16983
rect 32404 16940 32456 16949
rect 34060 17008 34112 17060
rect 37004 17187 37056 17196
rect 37004 17153 37013 17187
rect 37013 17153 37047 17187
rect 37047 17153 37056 17187
rect 37004 17144 37056 17153
rect 38752 17212 38804 17264
rect 41236 17212 41288 17264
rect 43076 17280 43128 17332
rect 42708 17212 42760 17264
rect 45652 17280 45704 17332
rect 46112 17280 46164 17332
rect 50528 17280 50580 17332
rect 50712 17280 50764 17332
rect 52368 17323 52420 17332
rect 52368 17289 52377 17323
rect 52377 17289 52411 17323
rect 52411 17289 52420 17323
rect 52368 17280 52420 17289
rect 53012 17280 53064 17332
rect 38384 17144 38436 17196
rect 38568 17187 38620 17196
rect 38568 17153 38577 17187
rect 38577 17153 38611 17187
rect 38611 17153 38620 17187
rect 38568 17144 38620 17153
rect 41052 17187 41104 17196
rect 38936 17076 38988 17128
rect 41052 17153 41061 17187
rect 41061 17153 41095 17187
rect 41095 17153 41104 17187
rect 41052 17144 41104 17153
rect 41328 17187 41380 17196
rect 41328 17153 41337 17187
rect 41337 17153 41371 17187
rect 41371 17153 41380 17187
rect 41328 17144 41380 17153
rect 41420 17144 41472 17196
rect 41696 17144 41748 17196
rect 42984 17144 43036 17196
rect 43444 17187 43496 17196
rect 43444 17153 43453 17187
rect 43453 17153 43487 17187
rect 43487 17153 43496 17187
rect 43444 17144 43496 17153
rect 43720 17187 43772 17196
rect 43720 17153 43729 17187
rect 43729 17153 43763 17187
rect 43763 17153 43772 17187
rect 43720 17144 43772 17153
rect 45468 17144 45520 17196
rect 45560 17187 45612 17196
rect 45560 17153 45569 17187
rect 45569 17153 45603 17187
rect 45603 17153 45612 17187
rect 45560 17144 45612 17153
rect 45744 17187 45796 17196
rect 45744 17153 45753 17187
rect 45753 17153 45787 17187
rect 45787 17153 45796 17187
rect 45744 17144 45796 17153
rect 45928 17255 45980 17264
rect 45928 17221 45937 17255
rect 45937 17221 45971 17255
rect 45971 17221 45980 17255
rect 45928 17212 45980 17221
rect 50620 17212 50672 17264
rect 54116 17255 54168 17264
rect 54116 17221 54125 17255
rect 54125 17221 54159 17255
rect 54159 17221 54168 17255
rect 54116 17212 54168 17221
rect 54484 17212 54536 17264
rect 46204 17144 46256 17196
rect 48044 17144 48096 17196
rect 49056 17144 49108 17196
rect 50344 17144 50396 17196
rect 40224 17076 40276 17128
rect 34152 16940 34204 16992
rect 34244 16983 34296 16992
rect 34244 16949 34253 16983
rect 34253 16949 34287 16983
rect 34287 16949 34296 16983
rect 34244 16940 34296 16949
rect 36452 16983 36504 16992
rect 36452 16949 36461 16983
rect 36461 16949 36495 16983
rect 36495 16949 36504 16983
rect 36452 16940 36504 16949
rect 37280 16940 37332 16992
rect 39948 16940 40000 16992
rect 42432 17076 42484 17128
rect 45008 17119 45060 17128
rect 45008 17085 45017 17119
rect 45017 17085 45051 17119
rect 45051 17085 45060 17119
rect 45008 17076 45060 17085
rect 46020 17076 46072 17128
rect 49700 17076 49752 17128
rect 41420 17008 41472 17060
rect 41328 16940 41380 16992
rect 41696 17051 41748 17060
rect 41696 17017 41705 17051
rect 41705 17017 41739 17051
rect 41739 17017 41748 17051
rect 41696 17008 41748 17017
rect 45836 17008 45888 17060
rect 50068 17008 50120 17060
rect 42340 16940 42392 16992
rect 43628 16983 43680 16992
rect 43628 16949 43637 16983
rect 43637 16949 43671 16983
rect 43671 16949 43680 16983
rect 43628 16940 43680 16949
rect 46296 16940 46348 16992
rect 48872 16940 48924 16992
rect 51264 16940 51316 16992
rect 53932 17187 53984 17196
rect 53932 17153 53942 17187
rect 53942 17153 53976 17187
rect 53976 17153 53984 17187
rect 53932 17144 53984 17153
rect 54208 17187 54260 17196
rect 54208 17153 54217 17187
rect 54217 17153 54251 17187
rect 54251 17153 54260 17187
rect 54208 17144 54260 17153
rect 54576 17144 54628 17196
rect 77852 17144 77904 17196
rect 78220 17051 78272 17060
rect 78220 17017 78229 17051
rect 78229 17017 78263 17051
rect 78263 17017 78272 17051
rect 78220 17008 78272 17017
rect 54116 16940 54168 16992
rect 54760 16940 54812 16992
rect 77852 16983 77904 16992
rect 77852 16949 77861 16983
rect 77861 16949 77895 16983
rect 77895 16949 77904 16983
rect 77852 16940 77904 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 14096 16736 14148 16788
rect 20444 16779 20496 16788
rect 20444 16745 20453 16779
rect 20453 16745 20487 16779
rect 20487 16745 20496 16779
rect 20444 16736 20496 16745
rect 17500 16668 17552 16720
rect 20628 16736 20680 16788
rect 20996 16736 21048 16788
rect 12624 16643 12676 16652
rect 12624 16609 12633 16643
rect 12633 16609 12667 16643
rect 12667 16609 12676 16643
rect 12624 16600 12676 16609
rect 12164 16532 12216 16584
rect 23480 16668 23532 16720
rect 18420 16600 18472 16652
rect 18972 16643 19024 16652
rect 18972 16609 18981 16643
rect 18981 16609 19015 16643
rect 19015 16609 19024 16643
rect 18972 16600 19024 16609
rect 22100 16600 22152 16652
rect 18052 16575 18104 16584
rect 18052 16541 18061 16575
rect 18061 16541 18095 16575
rect 18095 16541 18104 16575
rect 18052 16532 18104 16541
rect 19984 16532 20036 16584
rect 20076 16575 20128 16584
rect 20076 16541 20085 16575
rect 20085 16541 20119 16575
rect 20119 16541 20128 16575
rect 20076 16532 20128 16541
rect 21456 16532 21508 16584
rect 23112 16600 23164 16652
rect 23204 16575 23256 16584
rect 11520 16464 11572 16516
rect 12716 16464 12768 16516
rect 13636 16464 13688 16516
rect 18328 16464 18380 16516
rect 20812 16464 20864 16516
rect 23204 16541 23213 16575
rect 23213 16541 23247 16575
rect 23247 16541 23256 16575
rect 23204 16532 23256 16541
rect 25504 16736 25556 16788
rect 28172 16736 28224 16788
rect 28264 16779 28316 16788
rect 28264 16745 28273 16779
rect 28273 16745 28307 16779
rect 28307 16745 28316 16779
rect 28264 16736 28316 16745
rect 28540 16736 28592 16788
rect 29736 16736 29788 16788
rect 24768 16600 24820 16652
rect 28356 16668 28408 16720
rect 28908 16668 28960 16720
rect 32588 16736 32640 16788
rect 36544 16736 36596 16788
rect 38200 16736 38252 16788
rect 38384 16779 38436 16788
rect 38384 16745 38393 16779
rect 38393 16745 38427 16779
rect 38427 16745 38436 16779
rect 38384 16736 38436 16745
rect 41052 16736 41104 16788
rect 43168 16736 43220 16788
rect 45560 16736 45612 16788
rect 46020 16779 46072 16788
rect 46020 16745 46029 16779
rect 46029 16745 46063 16779
rect 46063 16745 46072 16779
rect 46020 16736 46072 16745
rect 46296 16779 46348 16788
rect 46296 16745 46305 16779
rect 46305 16745 46339 16779
rect 46339 16745 46348 16779
rect 46296 16736 46348 16745
rect 47676 16736 47728 16788
rect 37556 16668 37608 16720
rect 38476 16668 38528 16720
rect 24032 16532 24084 16584
rect 26240 16532 26292 16584
rect 26792 16575 26844 16584
rect 26792 16541 26801 16575
rect 26801 16541 26835 16575
rect 26835 16541 26844 16575
rect 26792 16532 26844 16541
rect 26884 16532 26936 16584
rect 36452 16643 36504 16652
rect 36452 16609 36461 16643
rect 36461 16609 36495 16643
rect 36495 16609 36504 16643
rect 36452 16600 36504 16609
rect 28540 16532 28592 16584
rect 31208 16532 31260 16584
rect 31576 16575 31628 16584
rect 31576 16541 31585 16575
rect 31585 16541 31619 16575
rect 31619 16541 31628 16575
rect 31576 16532 31628 16541
rect 33508 16532 33560 16584
rect 33876 16532 33928 16584
rect 40868 16600 40920 16652
rect 41328 16643 41380 16652
rect 41328 16609 41337 16643
rect 41337 16609 41371 16643
rect 41371 16609 41380 16643
rect 41328 16600 41380 16609
rect 42800 16600 42852 16652
rect 45008 16600 45060 16652
rect 45468 16668 45520 16720
rect 45744 16600 45796 16652
rect 38936 16575 38988 16584
rect 38936 16541 38944 16575
rect 38944 16541 38978 16575
rect 38978 16541 38988 16575
rect 38936 16532 38988 16541
rect 39028 16575 39080 16584
rect 39028 16541 39037 16575
rect 39037 16541 39071 16575
rect 39071 16541 39080 16575
rect 39028 16532 39080 16541
rect 39488 16532 39540 16584
rect 44364 16532 44416 16584
rect 49976 16736 50028 16788
rect 55312 16736 55364 16788
rect 12532 16396 12584 16448
rect 14924 16396 14976 16448
rect 17684 16439 17736 16448
rect 17684 16405 17693 16439
rect 17693 16405 17727 16439
rect 17727 16405 17736 16439
rect 17684 16396 17736 16405
rect 18512 16439 18564 16448
rect 18512 16405 18521 16439
rect 18521 16405 18555 16439
rect 18555 16405 18564 16439
rect 18512 16396 18564 16405
rect 20720 16396 20772 16448
rect 22744 16396 22796 16448
rect 26516 16507 26568 16516
rect 26516 16473 26525 16507
rect 26525 16473 26559 16507
rect 26559 16473 26568 16507
rect 26516 16464 26568 16473
rect 26608 16507 26660 16516
rect 26608 16473 26617 16507
rect 26617 16473 26651 16507
rect 26651 16473 26660 16507
rect 26608 16464 26660 16473
rect 27344 16464 27396 16516
rect 27804 16464 27856 16516
rect 31852 16507 31904 16516
rect 31852 16473 31861 16507
rect 31861 16473 31895 16507
rect 31895 16473 31904 16507
rect 31852 16464 31904 16473
rect 23572 16396 23624 16448
rect 23756 16439 23808 16448
rect 23756 16405 23765 16439
rect 23765 16405 23799 16439
rect 23799 16405 23808 16439
rect 23756 16396 23808 16405
rect 23848 16396 23900 16448
rect 25596 16396 25648 16448
rect 27528 16396 27580 16448
rect 27896 16396 27948 16448
rect 32680 16396 32732 16448
rect 35440 16464 35492 16516
rect 36084 16464 36136 16516
rect 36544 16464 36596 16516
rect 33508 16439 33560 16448
rect 33508 16405 33517 16439
rect 33517 16405 33551 16439
rect 33551 16405 33560 16439
rect 33508 16396 33560 16405
rect 35256 16396 35308 16448
rect 37096 16396 37148 16448
rect 39212 16464 39264 16516
rect 42616 16396 42668 16448
rect 44272 16396 44324 16448
rect 46112 16532 46164 16584
rect 46480 16575 46532 16584
rect 46480 16541 46489 16575
rect 46489 16541 46523 16575
rect 46523 16541 46532 16575
rect 46480 16532 46532 16541
rect 46848 16643 46900 16652
rect 46848 16609 46857 16643
rect 46857 16609 46891 16643
rect 46891 16609 46900 16643
rect 46848 16600 46900 16609
rect 47860 16600 47912 16652
rect 48228 16532 48280 16584
rect 48872 16575 48924 16584
rect 48872 16541 48881 16575
rect 48881 16541 48915 16575
rect 48915 16541 48924 16575
rect 48872 16532 48924 16541
rect 49332 16532 49384 16584
rect 47400 16464 47452 16516
rect 47308 16396 47360 16448
rect 48412 16396 48464 16448
rect 48688 16439 48740 16448
rect 48688 16405 48697 16439
rect 48697 16405 48731 16439
rect 48731 16405 48740 16439
rect 48688 16396 48740 16405
rect 48964 16507 49016 16516
rect 48964 16473 48973 16507
rect 48973 16473 49007 16507
rect 49007 16473 49016 16507
rect 48964 16464 49016 16473
rect 49056 16507 49108 16516
rect 49056 16473 49065 16507
rect 49065 16473 49099 16507
rect 49099 16473 49108 16507
rect 49056 16464 49108 16473
rect 49700 16507 49752 16516
rect 49700 16473 49709 16507
rect 49709 16473 49743 16507
rect 49743 16473 49752 16507
rect 49700 16464 49752 16473
rect 50344 16575 50396 16584
rect 50344 16541 50351 16575
rect 50351 16541 50396 16575
rect 50344 16532 50396 16541
rect 50804 16600 50856 16652
rect 51172 16600 51224 16652
rect 51356 16600 51408 16652
rect 51724 16600 51776 16652
rect 52644 16600 52696 16652
rect 50712 16532 50764 16584
rect 50068 16464 50120 16516
rect 50988 16464 51040 16516
rect 50896 16439 50948 16448
rect 50896 16405 50905 16439
rect 50905 16405 50939 16439
rect 50939 16405 50948 16439
rect 50896 16396 50948 16405
rect 51080 16396 51132 16448
rect 51264 16507 51316 16516
rect 51264 16473 51273 16507
rect 51273 16473 51307 16507
rect 51307 16473 51316 16507
rect 51264 16464 51316 16473
rect 51448 16575 51500 16584
rect 51448 16541 51457 16575
rect 51457 16541 51491 16575
rect 51491 16541 51500 16575
rect 51448 16532 51500 16541
rect 52552 16464 52604 16516
rect 54208 16532 54260 16584
rect 54760 16575 54812 16584
rect 54760 16541 54769 16575
rect 54769 16541 54803 16575
rect 54803 16541 54812 16575
rect 54760 16532 54812 16541
rect 54944 16575 54996 16584
rect 54944 16541 54953 16575
rect 54953 16541 54987 16575
rect 54987 16541 54996 16575
rect 54944 16532 54996 16541
rect 55036 16575 55088 16584
rect 55036 16541 55045 16575
rect 55045 16541 55079 16575
rect 55079 16541 55088 16575
rect 55036 16532 55088 16541
rect 55772 16575 55824 16584
rect 55772 16541 55781 16575
rect 55781 16541 55815 16575
rect 55815 16541 55824 16575
rect 55772 16532 55824 16541
rect 56416 16600 56468 16652
rect 55680 16464 55732 16516
rect 56140 16575 56192 16584
rect 56140 16541 56149 16575
rect 56149 16541 56183 16575
rect 56183 16541 56192 16575
rect 56140 16532 56192 16541
rect 51448 16396 51500 16448
rect 53748 16439 53800 16448
rect 53748 16405 53757 16439
rect 53757 16405 53791 16439
rect 53791 16405 53800 16439
rect 53748 16396 53800 16405
rect 53840 16439 53892 16448
rect 53840 16405 53849 16439
rect 53849 16405 53883 16439
rect 53883 16405 53892 16439
rect 53840 16396 53892 16405
rect 54576 16439 54628 16448
rect 54576 16405 54585 16439
rect 54585 16405 54619 16439
rect 54619 16405 54628 16439
rect 54576 16396 54628 16405
rect 57980 16396 58032 16448
rect 77852 16532 77904 16584
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 66314 16294 66366 16346
rect 66378 16294 66430 16346
rect 66442 16294 66494 16346
rect 66506 16294 66558 16346
rect 66570 16294 66622 16346
rect 1308 16056 1360 16108
rect 9496 16192 9548 16244
rect 12624 16192 12676 16244
rect 13360 16192 13412 16244
rect 17040 16235 17092 16244
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 17316 16192 17368 16244
rect 20812 16235 20864 16244
rect 20812 16201 20821 16235
rect 20821 16201 20855 16235
rect 20855 16201 20864 16235
rect 20812 16192 20864 16201
rect 23204 16192 23256 16244
rect 12256 16124 12308 16176
rect 14924 16124 14976 16176
rect 18512 16124 18564 16176
rect 11520 16099 11572 16108
rect 11520 16065 11529 16099
rect 11529 16065 11563 16099
rect 11563 16065 11572 16099
rect 11520 16056 11572 16065
rect 17132 16099 17184 16108
rect 17132 16065 17141 16099
rect 17141 16065 17175 16099
rect 17175 16065 17184 16099
rect 17132 16056 17184 16065
rect 17684 16056 17736 16108
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 20628 16056 20680 16108
rect 20720 16099 20772 16108
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 20812 16056 20864 16108
rect 21456 16056 21508 16108
rect 23296 16124 23348 16176
rect 24584 16235 24636 16244
rect 24584 16201 24593 16235
rect 24593 16201 24627 16235
rect 24627 16201 24636 16235
rect 24584 16192 24636 16201
rect 24768 16235 24820 16244
rect 24768 16201 24777 16235
rect 24777 16201 24811 16235
rect 24811 16201 24820 16235
rect 24768 16192 24820 16201
rect 26332 16192 26384 16244
rect 27252 16192 27304 16244
rect 23848 16124 23900 16176
rect 8300 15988 8352 16040
rect 11796 16031 11848 16040
rect 11796 15997 11805 16031
rect 11805 15997 11839 16031
rect 11839 15997 11848 16031
rect 11796 15988 11848 15997
rect 12256 15988 12308 16040
rect 12532 15988 12584 16040
rect 13636 16031 13688 16040
rect 13636 15997 13645 16031
rect 13645 15997 13679 16031
rect 13679 15997 13688 16031
rect 13636 15988 13688 15997
rect 14280 15988 14332 16040
rect 15752 15988 15804 16040
rect 20996 15988 21048 16040
rect 22928 15988 22980 16040
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 24400 16056 24452 16108
rect 24768 16056 24820 16108
rect 25596 16099 25648 16108
rect 25596 16065 25605 16099
rect 25605 16065 25639 16099
rect 25639 16065 25648 16099
rect 25596 16056 25648 16065
rect 26792 16124 26844 16176
rect 25964 16056 26016 16108
rect 27344 16124 27396 16176
rect 27528 16192 27580 16244
rect 31852 16192 31904 16244
rect 34796 16192 34848 16244
rect 38200 16192 38252 16244
rect 41512 16192 41564 16244
rect 42524 16192 42576 16244
rect 44456 16192 44508 16244
rect 27160 16056 27212 16108
rect 27988 16099 28040 16108
rect 27988 16065 27997 16099
rect 27997 16065 28031 16099
rect 28031 16065 28040 16099
rect 27988 16056 28040 16065
rect 29184 16124 29236 16176
rect 34244 16124 34296 16176
rect 29000 16056 29052 16108
rect 29552 16056 29604 16108
rect 32036 16056 32088 16108
rect 32404 16099 32456 16108
rect 32404 16065 32413 16099
rect 32413 16065 32447 16099
rect 32447 16065 32456 16099
rect 32404 16056 32456 16065
rect 32680 16099 32732 16108
rect 32680 16065 32689 16099
rect 32689 16065 32723 16099
rect 32723 16065 32732 16099
rect 32680 16056 32732 16065
rect 33232 16056 33284 16108
rect 33876 16099 33928 16108
rect 33876 16065 33885 16099
rect 33885 16065 33919 16099
rect 33919 16065 33928 16099
rect 33876 16056 33928 16065
rect 35256 16056 35308 16108
rect 44916 16235 44968 16244
rect 44916 16201 44925 16235
rect 44925 16201 44959 16235
rect 44959 16201 44968 16235
rect 44916 16192 44968 16201
rect 45652 16192 45704 16244
rect 46020 16192 46072 16244
rect 46480 16192 46532 16244
rect 26516 15988 26568 16040
rect 8116 15920 8168 15972
rect 16120 15920 16172 15972
rect 27252 15920 27304 15972
rect 27712 15920 27764 15972
rect 30012 15920 30064 15972
rect 33416 15988 33468 16040
rect 37004 15988 37056 16040
rect 45468 16099 45520 16108
rect 45468 16065 45477 16099
rect 45477 16065 45511 16099
rect 45511 16065 45520 16099
rect 45468 16056 45520 16065
rect 45744 16056 45796 16108
rect 46204 16056 46256 16108
rect 47400 16192 47452 16244
rect 47860 16124 47912 16176
rect 48412 16124 48464 16176
rect 49700 16124 49752 16176
rect 50160 16192 50212 16244
rect 50620 16192 50672 16244
rect 50804 16192 50856 16244
rect 45928 15988 45980 16040
rect 48504 16056 48556 16108
rect 48596 16099 48648 16108
rect 48596 16065 48605 16099
rect 48605 16065 48639 16099
rect 48639 16065 48648 16099
rect 48596 16056 48648 16065
rect 49516 16099 49568 16108
rect 49516 16065 49525 16099
rect 49525 16065 49559 16099
rect 49559 16065 49568 16099
rect 49516 16056 49568 16065
rect 50252 16056 50304 16108
rect 35256 15920 35308 15972
rect 36084 15920 36136 15972
rect 49056 15988 49108 16040
rect 49424 15988 49476 16040
rect 50436 16099 50488 16108
rect 50436 16065 50465 16099
rect 50465 16065 50488 16099
rect 50436 16056 50488 16065
rect 50896 16056 50948 16108
rect 14648 15852 14700 15904
rect 15476 15895 15528 15904
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 17408 15895 17460 15904
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 20536 15895 20588 15904
rect 20536 15861 20545 15895
rect 20545 15861 20579 15895
rect 20579 15861 20588 15895
rect 20536 15852 20588 15861
rect 21088 15895 21140 15904
rect 21088 15861 21097 15895
rect 21097 15861 21131 15895
rect 21131 15861 21140 15895
rect 21088 15852 21140 15861
rect 23388 15895 23440 15904
rect 23388 15861 23397 15895
rect 23397 15861 23431 15895
rect 23431 15861 23440 15895
rect 23388 15852 23440 15861
rect 25872 15895 25924 15904
rect 25872 15861 25881 15895
rect 25881 15861 25915 15895
rect 25915 15861 25924 15895
rect 25872 15852 25924 15861
rect 26332 15852 26384 15904
rect 29552 15852 29604 15904
rect 35992 15895 36044 15904
rect 35992 15861 36001 15895
rect 36001 15861 36035 15895
rect 36035 15861 36044 15895
rect 35992 15852 36044 15861
rect 39672 15852 39724 15904
rect 43352 15852 43404 15904
rect 46112 15852 46164 15904
rect 46756 15852 46808 15904
rect 48688 15852 48740 15904
rect 49332 15852 49384 15904
rect 49976 15895 50028 15904
rect 49976 15861 49985 15895
rect 49985 15861 50019 15895
rect 50019 15861 50028 15895
rect 49976 15852 50028 15861
rect 50712 15988 50764 16040
rect 51172 16099 51224 16108
rect 51172 16065 51181 16099
rect 51181 16065 51215 16099
rect 51215 16065 51224 16099
rect 51172 16056 51224 16065
rect 51356 16099 51408 16108
rect 51356 16065 51365 16099
rect 51365 16065 51399 16099
rect 51399 16065 51408 16099
rect 51356 16056 51408 16065
rect 51540 16056 51592 16108
rect 51908 16099 51960 16108
rect 51908 16065 51917 16099
rect 51917 16065 51951 16099
rect 51951 16065 51960 16099
rect 51908 16056 51960 16065
rect 52368 16192 52420 16244
rect 50436 15920 50488 15972
rect 52276 16099 52328 16108
rect 52276 16065 52285 16099
rect 52285 16065 52319 16099
rect 52319 16065 52328 16099
rect 52276 16056 52328 16065
rect 52460 16056 52512 16108
rect 52644 16192 52696 16244
rect 54944 16192 54996 16244
rect 56140 16192 56192 16244
rect 57980 16235 58032 16244
rect 57980 16201 57989 16235
rect 57989 16201 58023 16235
rect 58023 16201 58032 16235
rect 57980 16192 58032 16201
rect 53380 16167 53432 16176
rect 53380 16133 53389 16167
rect 53389 16133 53423 16167
rect 53423 16133 53432 16167
rect 53380 16124 53432 16133
rect 54576 16124 54628 16176
rect 55680 16124 55732 16176
rect 53840 16056 53892 16108
rect 54024 15988 54076 16040
rect 55036 15988 55088 16040
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 8300 15691 8352 15700
rect 8300 15657 8309 15691
rect 8309 15657 8343 15691
rect 8343 15657 8352 15691
rect 8300 15648 8352 15657
rect 11796 15691 11848 15700
rect 11796 15657 11805 15691
rect 11805 15657 11839 15691
rect 11839 15657 11848 15691
rect 11796 15648 11848 15657
rect 14280 15691 14332 15700
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 19708 15691 19760 15700
rect 12440 15555 12492 15564
rect 12440 15521 12449 15555
rect 12449 15521 12483 15555
rect 12483 15521 12492 15555
rect 12440 15512 12492 15521
rect 13360 15555 13412 15564
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13360 15512 13412 15521
rect 15476 15580 15528 15632
rect 15016 15512 15068 15564
rect 15752 15555 15804 15564
rect 15752 15521 15761 15555
rect 15761 15521 15795 15555
rect 15795 15521 15804 15555
rect 15752 15512 15804 15521
rect 19708 15657 19717 15691
rect 19717 15657 19751 15691
rect 19751 15657 19760 15691
rect 19708 15648 19760 15657
rect 24124 15648 24176 15700
rect 25136 15648 25188 15700
rect 27804 15648 27856 15700
rect 29000 15648 29052 15700
rect 19524 15580 19576 15632
rect 22100 15580 22152 15632
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 8116 15487 8168 15496
rect 8116 15453 8125 15487
rect 8125 15453 8159 15487
rect 8159 15453 8168 15487
rect 8116 15444 8168 15453
rect 12164 15487 12216 15496
rect 12164 15453 12173 15487
rect 12173 15453 12207 15487
rect 12207 15453 12216 15487
rect 12164 15444 12216 15453
rect 14648 15487 14700 15496
rect 14648 15453 14657 15487
rect 14657 15453 14691 15487
rect 14691 15453 14700 15487
rect 14648 15444 14700 15453
rect 18604 15444 18656 15496
rect 18972 15444 19024 15496
rect 19616 15444 19668 15496
rect 7932 15376 7984 15428
rect 20628 15512 20680 15564
rect 20352 15487 20404 15496
rect 20352 15453 20361 15487
rect 20361 15453 20395 15487
rect 20395 15453 20404 15487
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 21456 15512 21508 15564
rect 20352 15444 20404 15453
rect 20720 15419 20772 15428
rect 20720 15385 20729 15419
rect 20729 15385 20763 15419
rect 20763 15385 20772 15419
rect 20720 15376 20772 15385
rect 21088 15487 21140 15496
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 22744 15487 22796 15496
rect 22744 15453 22753 15487
rect 22753 15453 22787 15487
rect 22787 15453 22796 15487
rect 22744 15444 22796 15453
rect 24032 15580 24084 15632
rect 24768 15580 24820 15632
rect 27988 15580 28040 15632
rect 25320 15555 25372 15564
rect 25320 15521 25329 15555
rect 25329 15521 25363 15555
rect 25363 15521 25372 15555
rect 25320 15512 25372 15521
rect 25872 15512 25924 15564
rect 26148 15512 26200 15564
rect 23020 15487 23072 15496
rect 23020 15453 23029 15487
rect 23029 15453 23063 15487
rect 23063 15453 23072 15487
rect 23020 15444 23072 15453
rect 23204 15487 23256 15496
rect 23204 15453 23213 15487
rect 23213 15453 23247 15487
rect 23247 15453 23256 15487
rect 23204 15444 23256 15453
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 25504 15487 25556 15496
rect 25504 15453 25513 15487
rect 25513 15453 25547 15487
rect 25547 15453 25556 15487
rect 25504 15444 25556 15453
rect 25964 15444 26016 15496
rect 26424 15487 26476 15496
rect 26424 15453 26433 15487
rect 26433 15453 26467 15487
rect 26467 15453 26476 15487
rect 26424 15444 26476 15453
rect 27436 15512 27488 15564
rect 27252 15487 27304 15496
rect 27252 15453 27261 15487
rect 27261 15453 27295 15487
rect 27295 15453 27304 15487
rect 27252 15444 27304 15453
rect 27712 15487 27764 15496
rect 27712 15453 27721 15487
rect 27721 15453 27755 15487
rect 27755 15453 27764 15487
rect 27712 15444 27764 15453
rect 28816 15487 28868 15496
rect 28816 15453 28825 15487
rect 28825 15453 28859 15487
rect 28859 15453 28868 15487
rect 28816 15444 28868 15453
rect 21088 15308 21140 15360
rect 22928 15376 22980 15428
rect 27068 15376 27120 15428
rect 27528 15376 27580 15428
rect 29552 15444 29604 15496
rect 29736 15487 29788 15496
rect 29736 15453 29745 15487
rect 29745 15453 29779 15487
rect 29779 15453 29788 15487
rect 29736 15444 29788 15453
rect 31116 15444 31168 15496
rect 22468 15308 22520 15360
rect 23940 15308 23992 15360
rect 25504 15308 25556 15360
rect 26976 15308 27028 15360
rect 31576 15376 31628 15428
rect 33232 15376 33284 15428
rect 38752 15648 38804 15700
rect 40592 15648 40644 15700
rect 41420 15648 41472 15700
rect 42616 15648 42668 15700
rect 45928 15648 45980 15700
rect 46756 15648 46808 15700
rect 49884 15691 49936 15700
rect 49884 15657 49893 15691
rect 49893 15657 49927 15691
rect 49927 15657 49936 15691
rect 49884 15648 49936 15657
rect 51172 15648 51224 15700
rect 53380 15648 53432 15700
rect 34428 15580 34480 15632
rect 35992 15580 36044 15632
rect 35440 15555 35492 15564
rect 35440 15521 35449 15555
rect 35449 15521 35483 15555
rect 35483 15521 35492 15555
rect 35440 15512 35492 15521
rect 33692 15444 33744 15496
rect 34796 15444 34848 15496
rect 35348 15444 35400 15496
rect 33508 15308 33560 15360
rect 34244 15376 34296 15428
rect 34336 15376 34388 15428
rect 37372 15580 37424 15632
rect 37004 15444 37056 15496
rect 37280 15376 37332 15428
rect 37648 15376 37700 15428
rect 37740 15351 37792 15360
rect 37740 15317 37749 15351
rect 37749 15317 37783 15351
rect 37783 15317 37792 15351
rect 37740 15308 37792 15317
rect 37924 15487 37976 15496
rect 37924 15453 37933 15487
rect 37933 15453 37967 15487
rect 37967 15453 37976 15487
rect 37924 15444 37976 15453
rect 49608 15580 49660 15632
rect 50896 15580 50948 15632
rect 38568 15555 38620 15564
rect 38568 15521 38577 15555
rect 38577 15521 38611 15555
rect 38611 15521 38620 15555
rect 38568 15512 38620 15521
rect 40868 15512 40920 15564
rect 39304 15444 39356 15496
rect 45744 15512 45796 15564
rect 46848 15512 46900 15564
rect 49884 15512 49936 15564
rect 43536 15444 43588 15496
rect 48136 15444 48188 15496
rect 52276 15512 52328 15564
rect 54944 15512 54996 15564
rect 50896 15444 50948 15496
rect 54208 15444 54260 15496
rect 40040 15376 40092 15428
rect 40132 15419 40184 15428
rect 40132 15385 40141 15419
rect 40141 15385 40175 15419
rect 40175 15385 40184 15419
rect 40132 15376 40184 15385
rect 41420 15376 41472 15428
rect 41604 15351 41656 15360
rect 41604 15317 41613 15351
rect 41613 15317 41647 15351
rect 41647 15317 41656 15351
rect 41604 15308 41656 15317
rect 42156 15419 42208 15428
rect 42156 15385 42165 15419
rect 42165 15385 42199 15419
rect 42199 15385 42208 15419
rect 42156 15376 42208 15385
rect 42616 15376 42668 15428
rect 45836 15376 45888 15428
rect 48964 15376 49016 15428
rect 50988 15376 51040 15428
rect 53840 15376 53892 15428
rect 54668 15487 54720 15496
rect 54668 15453 54677 15487
rect 54677 15453 54711 15487
rect 54711 15453 54720 15487
rect 54668 15444 54720 15453
rect 55496 15487 55548 15496
rect 55496 15453 55505 15487
rect 55505 15453 55539 15487
rect 55539 15453 55548 15487
rect 55496 15444 55548 15453
rect 55772 15555 55824 15564
rect 55772 15521 55781 15555
rect 55781 15521 55815 15555
rect 55815 15521 55824 15555
rect 55772 15512 55824 15521
rect 54484 15419 54536 15428
rect 54484 15385 54493 15419
rect 54493 15385 54527 15419
rect 54527 15385 54536 15419
rect 54484 15376 54536 15385
rect 55956 15487 56008 15496
rect 55956 15453 55965 15487
rect 55965 15453 55999 15487
rect 55999 15453 56008 15487
rect 55956 15444 56008 15453
rect 43444 15308 43496 15360
rect 43536 15308 43588 15360
rect 43720 15351 43772 15360
rect 43720 15317 43729 15351
rect 43729 15317 43763 15351
rect 43763 15317 43772 15351
rect 43720 15308 43772 15317
rect 45468 15308 45520 15360
rect 47492 15308 47544 15360
rect 48596 15308 48648 15360
rect 49976 15308 50028 15360
rect 50896 15351 50948 15360
rect 50896 15317 50905 15351
rect 50905 15317 50939 15351
rect 50939 15317 50948 15351
rect 50896 15308 50948 15317
rect 56508 15376 56560 15428
rect 55220 15308 55272 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 66314 15206 66366 15258
rect 66378 15206 66430 15258
rect 66442 15206 66494 15258
rect 66506 15206 66558 15258
rect 66570 15206 66622 15258
rect 7656 14968 7708 15020
rect 8116 15104 8168 15156
rect 17132 15104 17184 15156
rect 7932 15011 7984 15020
rect 7932 14977 7941 15011
rect 7941 14977 7975 15011
rect 7975 14977 7984 15011
rect 7932 14968 7984 14977
rect 8576 14968 8628 15020
rect 9772 15036 9824 15088
rect 20352 15036 20404 15088
rect 20628 15036 20680 15088
rect 9496 15011 9548 15020
rect 9496 14977 9505 15011
rect 9505 14977 9539 15011
rect 9539 14977 9548 15011
rect 9496 14968 9548 14977
rect 10876 14968 10928 15020
rect 12256 14968 12308 15020
rect 12348 14968 12400 15020
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 13452 14900 13504 14952
rect 16948 14943 17000 14952
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 18604 15011 18656 15020
rect 18604 14977 18613 15011
rect 18613 14977 18647 15011
rect 18647 14977 18656 15011
rect 18604 14968 18656 14977
rect 23020 15036 23072 15088
rect 22744 14968 22796 15020
rect 22928 15011 22980 15020
rect 22928 14977 22937 15011
rect 22937 14977 22971 15011
rect 22971 14977 22980 15011
rect 22928 14968 22980 14977
rect 24032 15036 24084 15088
rect 26424 15104 26476 15156
rect 28908 15104 28960 15156
rect 33232 15104 33284 15156
rect 19616 14943 19668 14952
rect 19616 14909 19625 14943
rect 19625 14909 19659 14943
rect 19659 14909 19668 14943
rect 19616 14900 19668 14909
rect 19708 14900 19760 14952
rect 25320 15011 25372 15020
rect 25320 14977 25329 15011
rect 25329 14977 25363 15011
rect 25363 14977 25372 15011
rect 25320 14968 25372 14977
rect 25504 15011 25556 15020
rect 25504 14977 25513 15011
rect 25513 14977 25547 15011
rect 25547 14977 25556 15011
rect 25504 14968 25556 14977
rect 31484 15036 31536 15088
rect 26976 14968 27028 15020
rect 27068 15011 27120 15020
rect 27068 14977 27077 15011
rect 27077 14977 27111 15011
rect 27111 14977 27120 15011
rect 27068 14968 27120 14977
rect 27160 15011 27212 15020
rect 27160 14977 27170 15011
rect 27170 14977 27204 15011
rect 27204 14977 27212 15011
rect 27160 14968 27212 14977
rect 27712 14968 27764 15020
rect 28356 14968 28408 15020
rect 28632 15011 28684 15020
rect 28632 14977 28641 15011
rect 28641 14977 28675 15011
rect 28675 14977 28684 15011
rect 28632 14968 28684 14977
rect 28724 14968 28776 15020
rect 29184 14968 29236 15020
rect 32220 14968 32272 15020
rect 33140 14968 33192 15020
rect 33232 15011 33284 15020
rect 33232 14977 33241 15011
rect 33241 14977 33275 15011
rect 33275 14977 33284 15011
rect 33232 14968 33284 14977
rect 35440 15036 35492 15088
rect 37648 15104 37700 15156
rect 37740 15036 37792 15088
rect 39120 15036 39172 15088
rect 39396 15036 39448 15088
rect 14280 14764 14332 14816
rect 18972 14807 19024 14816
rect 18972 14773 18981 14807
rect 18981 14773 19015 14807
rect 19015 14773 19024 14807
rect 18972 14764 19024 14773
rect 19064 14807 19116 14816
rect 19064 14773 19073 14807
rect 19073 14773 19107 14807
rect 19107 14773 19116 14807
rect 19064 14764 19116 14773
rect 19248 14832 19300 14884
rect 19524 14832 19576 14884
rect 21088 14832 21140 14884
rect 22468 14832 22520 14884
rect 25596 14832 25648 14884
rect 25964 14832 26016 14884
rect 30012 14832 30064 14884
rect 33232 14832 33284 14884
rect 22652 14807 22704 14816
rect 22652 14773 22661 14807
rect 22661 14773 22695 14807
rect 22695 14773 22704 14807
rect 22652 14764 22704 14773
rect 22744 14764 22796 14816
rect 23296 14764 23348 14816
rect 25136 14764 25188 14816
rect 27804 14764 27856 14816
rect 28724 14807 28776 14816
rect 28724 14773 28733 14807
rect 28733 14773 28767 14807
rect 28767 14773 28776 14807
rect 28724 14764 28776 14773
rect 33508 14943 33560 14952
rect 33508 14909 33517 14943
rect 33517 14909 33551 14943
rect 33551 14909 33560 14943
rect 33508 14900 33560 14909
rect 34704 14832 34756 14884
rect 36084 14900 36136 14952
rect 39488 15011 39540 15020
rect 39488 14977 39497 15011
rect 39497 14977 39531 15011
rect 39531 14977 39540 15011
rect 39488 14968 39540 14977
rect 39672 15011 39724 15020
rect 39672 14977 39679 15011
rect 39679 14977 39724 15011
rect 39672 14968 39724 14977
rect 39764 15011 39816 15020
rect 39764 14977 39773 15011
rect 39773 14977 39807 15011
rect 39807 14977 39816 15011
rect 39764 14968 39816 14977
rect 40132 15104 40184 15156
rect 42156 15104 42208 15156
rect 43352 15147 43404 15156
rect 43352 15113 43361 15147
rect 43361 15113 43395 15147
rect 43395 15113 43404 15147
rect 43352 15104 43404 15113
rect 43444 15104 43496 15156
rect 48136 15104 48188 15156
rect 48228 15104 48280 15156
rect 55956 15104 56008 15156
rect 56508 15104 56560 15156
rect 41052 15011 41104 15020
rect 41052 14977 41061 15011
rect 41061 14977 41095 15011
rect 41095 14977 41104 15011
rect 41052 14968 41104 14977
rect 41604 14968 41656 15020
rect 41788 15011 41840 15020
rect 41788 14977 41797 15011
rect 41797 14977 41831 15011
rect 41831 14977 41840 15011
rect 41788 14968 41840 14977
rect 42064 14968 42116 15020
rect 42984 14968 43036 15020
rect 43996 14968 44048 15020
rect 45560 14968 45612 15020
rect 46664 14968 46716 15020
rect 48044 15011 48096 15020
rect 48044 14977 48053 15011
rect 48053 14977 48087 15011
rect 48087 14977 48096 15011
rect 48044 14968 48096 14977
rect 48136 15011 48188 15020
rect 48136 14977 48145 15011
rect 48145 14977 48179 15011
rect 48179 14977 48188 15011
rect 48136 14968 48188 14977
rect 55220 15036 55272 15088
rect 55588 15036 55640 15088
rect 43720 14900 43772 14952
rect 45376 14900 45428 14952
rect 47952 14900 48004 14952
rect 49700 14900 49752 14952
rect 41420 14832 41472 14884
rect 44364 14832 44416 14884
rect 34244 14764 34296 14816
rect 34796 14764 34848 14816
rect 36544 14764 36596 14816
rect 37004 14807 37056 14816
rect 37004 14773 37013 14807
rect 37013 14773 37047 14807
rect 37047 14773 37056 14807
rect 37004 14764 37056 14773
rect 39304 14807 39356 14816
rect 39304 14773 39313 14807
rect 39313 14773 39347 14807
rect 39347 14773 39356 14807
rect 39304 14764 39356 14773
rect 42156 14807 42208 14816
rect 42156 14773 42165 14807
rect 42165 14773 42199 14807
rect 42199 14773 42208 14807
rect 42156 14764 42208 14773
rect 43628 14764 43680 14816
rect 44088 14807 44140 14816
rect 44088 14773 44097 14807
rect 44097 14773 44131 14807
rect 44131 14773 44140 14807
rect 44088 14764 44140 14773
rect 45008 14764 45060 14816
rect 47124 14764 47176 14816
rect 47860 14807 47912 14816
rect 47860 14773 47869 14807
rect 47869 14773 47903 14807
rect 47903 14773 47912 14807
rect 47860 14764 47912 14773
rect 48780 14764 48832 14816
rect 49516 14764 49568 14816
rect 54024 14968 54076 15020
rect 51540 14832 51592 14884
rect 50620 14807 50672 14816
rect 50620 14773 50629 14807
rect 50629 14773 50663 14807
rect 50663 14773 50672 14807
rect 50620 14764 50672 14773
rect 51816 14764 51868 14816
rect 54208 14807 54260 14816
rect 54208 14773 54217 14807
rect 54217 14773 54251 14807
rect 54251 14773 54260 14807
rect 54208 14764 54260 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 8576 14560 8628 14612
rect 17960 14560 18012 14612
rect 18972 14560 19024 14612
rect 19708 14603 19760 14612
rect 19708 14569 19717 14603
rect 19717 14569 19751 14603
rect 19751 14569 19760 14603
rect 19708 14560 19760 14569
rect 20812 14560 20864 14612
rect 22652 14560 22704 14612
rect 23204 14603 23256 14612
rect 23204 14569 23213 14603
rect 23213 14569 23247 14603
rect 23247 14569 23256 14603
rect 23204 14560 23256 14569
rect 28172 14603 28224 14612
rect 28172 14569 28181 14603
rect 28181 14569 28215 14603
rect 28215 14569 28224 14603
rect 28172 14560 28224 14569
rect 30656 14560 30708 14612
rect 32036 14560 32088 14612
rect 33048 14560 33100 14612
rect 33232 14560 33284 14612
rect 34428 14560 34480 14612
rect 35348 14560 35400 14612
rect 37924 14560 37976 14612
rect 42064 14603 42116 14612
rect 42064 14569 42073 14603
rect 42073 14569 42107 14603
rect 42107 14569 42116 14603
rect 42064 14560 42116 14569
rect 42340 14560 42392 14612
rect 43076 14560 43128 14612
rect 43904 14560 43956 14612
rect 43996 14603 44048 14612
rect 43996 14569 44005 14603
rect 44005 14569 44039 14603
rect 44039 14569 44048 14603
rect 43996 14560 44048 14569
rect 14096 14535 14148 14544
rect 14096 14501 14105 14535
rect 14105 14501 14139 14535
rect 14139 14501 14148 14535
rect 14096 14492 14148 14501
rect 12440 14424 12492 14476
rect 1216 14356 1268 14408
rect 7656 14399 7708 14408
rect 7656 14365 7665 14399
rect 7665 14365 7699 14399
rect 7699 14365 7708 14399
rect 7656 14356 7708 14365
rect 12348 14399 12400 14408
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 16488 14424 16540 14476
rect 16948 14424 17000 14476
rect 19616 14424 19668 14476
rect 20536 14467 20588 14476
rect 20536 14433 20545 14467
rect 20545 14433 20579 14467
rect 20579 14433 20588 14467
rect 20536 14424 20588 14433
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 14464 14356 14516 14408
rect 18512 14356 18564 14408
rect 19064 14356 19116 14408
rect 21456 14356 21508 14408
rect 22376 14356 22428 14408
rect 24768 14492 24820 14544
rect 23296 14467 23348 14476
rect 23296 14433 23305 14467
rect 23305 14433 23339 14467
rect 23339 14433 23348 14467
rect 23296 14424 23348 14433
rect 23572 14424 23624 14476
rect 24860 14424 24912 14476
rect 23112 14356 23164 14408
rect 23388 14356 23440 14408
rect 27712 14492 27764 14544
rect 27160 14424 27212 14476
rect 26884 14356 26936 14408
rect 27344 14399 27396 14408
rect 27344 14365 27353 14399
rect 27353 14365 27387 14399
rect 27387 14365 27396 14399
rect 27344 14356 27396 14365
rect 27528 14356 27580 14408
rect 15108 14288 15160 14340
rect 15200 14331 15252 14340
rect 15200 14297 15209 14331
rect 15209 14297 15243 14331
rect 15243 14297 15252 14331
rect 15200 14288 15252 14297
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 11796 14220 11848 14272
rect 14464 14263 14516 14272
rect 14464 14229 14473 14263
rect 14473 14229 14507 14263
rect 14507 14229 14516 14263
rect 14464 14220 14516 14229
rect 14924 14220 14976 14272
rect 16764 14263 16816 14272
rect 16764 14229 16773 14263
rect 16773 14229 16807 14263
rect 16807 14229 16816 14263
rect 16764 14220 16816 14229
rect 23296 14288 23348 14340
rect 18328 14220 18380 14272
rect 20904 14220 20956 14272
rect 22560 14263 22612 14272
rect 22560 14229 22569 14263
rect 22569 14229 22603 14263
rect 22603 14229 22612 14263
rect 22560 14220 22612 14229
rect 22652 14220 22704 14272
rect 23388 14220 23440 14272
rect 23664 14220 23716 14272
rect 24768 14288 24820 14340
rect 26976 14288 27028 14340
rect 28080 14424 28132 14476
rect 33876 14492 33928 14544
rect 24308 14220 24360 14272
rect 26240 14220 26292 14272
rect 28080 14220 28132 14272
rect 29460 14424 29512 14476
rect 29736 14424 29788 14476
rect 31576 14424 31628 14476
rect 29552 14356 29604 14408
rect 30932 14356 30984 14408
rect 33140 14399 33192 14408
rect 33140 14365 33149 14399
rect 33149 14365 33183 14399
rect 33183 14365 33192 14399
rect 33140 14356 33192 14365
rect 33416 14399 33468 14408
rect 33416 14365 33425 14399
rect 33425 14365 33459 14399
rect 33459 14365 33468 14399
rect 33416 14356 33468 14365
rect 39672 14492 39724 14544
rect 35808 14424 35860 14476
rect 31576 14331 31628 14340
rect 31576 14297 31585 14331
rect 31585 14297 31619 14331
rect 31619 14297 31628 14331
rect 31576 14288 31628 14297
rect 32864 14288 32916 14340
rect 33508 14288 33560 14340
rect 34796 14288 34848 14340
rect 35808 14331 35860 14340
rect 35808 14297 35817 14331
rect 35817 14297 35851 14331
rect 35851 14297 35860 14331
rect 35808 14288 35860 14297
rect 30380 14220 30432 14272
rect 31944 14220 31996 14272
rect 33968 14220 34020 14272
rect 34152 14220 34204 14272
rect 35348 14220 35400 14272
rect 36176 14399 36228 14408
rect 36176 14365 36185 14399
rect 36185 14365 36219 14399
rect 36219 14365 36228 14399
rect 36176 14356 36228 14365
rect 36820 14424 36872 14476
rect 37188 14424 37240 14476
rect 37280 14424 37332 14476
rect 37556 14424 37608 14476
rect 36636 14399 36688 14408
rect 36636 14365 36645 14399
rect 36645 14365 36679 14399
rect 36679 14365 36688 14399
rect 36636 14356 36688 14365
rect 36360 14288 36412 14340
rect 36544 14331 36596 14340
rect 36544 14297 36553 14331
rect 36553 14297 36587 14331
rect 36587 14297 36596 14331
rect 36544 14288 36596 14297
rect 39764 14424 39816 14476
rect 39856 14424 39908 14476
rect 37004 14288 37056 14340
rect 36820 14263 36872 14272
rect 36820 14229 36829 14263
rect 36829 14229 36863 14263
rect 36863 14229 36872 14263
rect 36820 14220 36872 14229
rect 36912 14263 36964 14272
rect 36912 14229 36921 14263
rect 36921 14229 36955 14263
rect 36955 14229 36964 14263
rect 36912 14220 36964 14229
rect 37740 14220 37792 14272
rect 39488 14356 39540 14408
rect 42340 14424 42392 14476
rect 41512 14399 41564 14408
rect 41512 14365 41522 14399
rect 41522 14365 41556 14399
rect 41556 14365 41564 14399
rect 41512 14356 41564 14365
rect 41788 14399 41840 14408
rect 41788 14365 41797 14399
rect 41797 14365 41831 14399
rect 41831 14365 41840 14399
rect 41788 14356 41840 14365
rect 42156 14356 42208 14408
rect 43352 14492 43404 14544
rect 44916 14492 44968 14544
rect 47492 14603 47544 14612
rect 47492 14569 47501 14603
rect 47501 14569 47535 14603
rect 47535 14569 47544 14603
rect 47492 14560 47544 14569
rect 47768 14492 47820 14544
rect 42800 14399 42852 14408
rect 42800 14365 42809 14399
rect 42809 14365 42843 14399
rect 42843 14365 42852 14399
rect 42800 14356 42852 14365
rect 43628 14424 43680 14476
rect 41696 14331 41748 14340
rect 41696 14297 41705 14331
rect 41705 14297 41739 14331
rect 41739 14297 41748 14331
rect 41696 14288 41748 14297
rect 43536 14356 43588 14408
rect 44640 14424 44692 14476
rect 45100 14424 45152 14476
rect 45744 14467 45796 14476
rect 45744 14433 45753 14467
rect 45753 14433 45787 14467
rect 45787 14433 45796 14467
rect 45744 14424 45796 14433
rect 46756 14424 46808 14476
rect 41880 14220 41932 14272
rect 42248 14263 42300 14272
rect 42248 14229 42257 14263
rect 42257 14229 42291 14263
rect 42291 14229 42300 14263
rect 42248 14220 42300 14229
rect 44364 14288 44416 14340
rect 45008 14331 45060 14340
rect 45008 14297 45017 14331
rect 45017 14297 45051 14331
rect 45051 14297 45060 14331
rect 45008 14288 45060 14297
rect 45192 14331 45244 14340
rect 45192 14297 45201 14331
rect 45201 14297 45235 14331
rect 45235 14297 45244 14331
rect 45192 14288 45244 14297
rect 47308 14356 47360 14408
rect 47584 14356 47636 14408
rect 50804 14560 50856 14612
rect 48136 14399 48188 14408
rect 48136 14365 48150 14399
rect 48150 14365 48184 14399
rect 48184 14365 48188 14399
rect 50436 14492 50488 14544
rect 49700 14424 49752 14476
rect 49884 14424 49936 14476
rect 48136 14356 48188 14365
rect 48780 14399 48832 14408
rect 48780 14365 48789 14399
rect 48789 14365 48823 14399
rect 48823 14365 48832 14399
rect 48780 14356 48832 14365
rect 46020 14331 46072 14340
rect 46020 14297 46029 14331
rect 46029 14297 46063 14331
rect 46063 14297 46072 14331
rect 46020 14288 46072 14297
rect 47952 14331 48004 14340
rect 45284 14220 45336 14272
rect 47952 14297 47961 14331
rect 47961 14297 47995 14331
rect 47995 14297 48004 14331
rect 47952 14288 48004 14297
rect 50436 14399 50488 14408
rect 50436 14365 50445 14399
rect 50445 14365 50479 14399
rect 50479 14365 50488 14399
rect 50436 14356 50488 14365
rect 51080 14560 51132 14612
rect 53564 14603 53616 14612
rect 53564 14569 53573 14603
rect 53573 14569 53607 14603
rect 53607 14569 53616 14603
rect 53564 14560 53616 14569
rect 51356 14492 51408 14544
rect 50988 14424 51040 14476
rect 54208 14492 54260 14544
rect 51540 14399 51592 14408
rect 51540 14365 51573 14399
rect 51573 14365 51592 14399
rect 51540 14356 51592 14365
rect 51724 14356 51776 14408
rect 53564 14356 53616 14408
rect 54576 14399 54628 14408
rect 54576 14365 54580 14399
rect 54580 14365 54614 14399
rect 54614 14365 54628 14399
rect 47492 14220 47544 14272
rect 50988 14288 51040 14340
rect 52092 14331 52144 14340
rect 52092 14297 52101 14331
rect 52101 14297 52135 14331
rect 52135 14297 52144 14331
rect 52092 14288 52144 14297
rect 52552 14288 52604 14340
rect 53472 14288 53524 14340
rect 54576 14356 54628 14365
rect 54760 14399 54812 14408
rect 54760 14365 54769 14399
rect 54769 14365 54803 14399
rect 54803 14365 54812 14399
rect 54760 14356 54812 14365
rect 54944 14399 54996 14408
rect 54944 14365 54952 14399
rect 54952 14365 54986 14399
rect 54986 14365 54996 14399
rect 54944 14356 54996 14365
rect 48412 14263 48464 14272
rect 48412 14229 48421 14263
rect 48421 14229 48455 14263
rect 48455 14229 48464 14263
rect 48412 14220 48464 14229
rect 50252 14220 50304 14272
rect 50436 14220 50488 14272
rect 50620 14220 50672 14272
rect 51264 14220 51316 14272
rect 52184 14220 52236 14272
rect 54116 14220 54168 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 66314 14118 66366 14170
rect 66378 14118 66430 14170
rect 66442 14118 66494 14170
rect 66506 14118 66558 14170
rect 66570 14118 66622 14170
rect 7656 14016 7708 14068
rect 7840 13948 7892 14000
rect 10876 13948 10928 14000
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 12716 14016 12768 14068
rect 13452 14016 13504 14068
rect 15200 14016 15252 14068
rect 16764 14016 16816 14068
rect 21456 14059 21508 14068
rect 21456 14025 21465 14059
rect 21465 14025 21499 14059
rect 21499 14025 21508 14059
rect 21456 14016 21508 14025
rect 23112 14016 23164 14068
rect 11796 13991 11848 14000
rect 11796 13957 11805 13991
rect 11805 13957 11839 13991
rect 11839 13957 11848 13991
rect 11796 13948 11848 13957
rect 12256 13948 12308 14000
rect 1400 13880 1452 13889
rect 9404 13812 9456 13864
rect 16856 13880 16908 13932
rect 17408 13880 17460 13932
rect 17960 13923 18012 13932
rect 17960 13889 17969 13923
rect 17969 13889 18003 13923
rect 18003 13889 18012 13923
rect 17960 13880 18012 13889
rect 19248 13880 19300 13932
rect 22376 13923 22428 13932
rect 22376 13889 22385 13923
rect 22385 13889 22419 13923
rect 22419 13889 22428 13923
rect 22376 13880 22428 13889
rect 22468 13880 22520 13932
rect 22744 13923 22796 13932
rect 22744 13889 22753 13923
rect 22753 13889 22787 13923
rect 22787 13889 22796 13923
rect 22744 13880 22796 13889
rect 16396 13855 16448 13864
rect 16396 13821 16405 13855
rect 16405 13821 16439 13855
rect 16439 13821 16448 13855
rect 16396 13812 16448 13821
rect 23020 13880 23072 13932
rect 23388 13948 23440 14000
rect 25504 14016 25556 14068
rect 23480 13880 23532 13932
rect 23664 13923 23716 13932
rect 23664 13889 23673 13923
rect 23673 13889 23707 13923
rect 23707 13889 23716 13923
rect 23664 13880 23716 13889
rect 23848 13923 23900 13932
rect 23848 13889 23855 13923
rect 23855 13889 23900 13923
rect 23848 13880 23900 13889
rect 23940 13923 23992 13932
rect 23940 13889 23949 13923
rect 23949 13889 23983 13923
rect 23983 13889 23992 13923
rect 23940 13880 23992 13889
rect 24124 13923 24176 13932
rect 27528 13991 27580 14000
rect 27528 13957 27537 13991
rect 27537 13957 27571 13991
rect 27571 13957 27580 13991
rect 27528 13948 27580 13957
rect 28816 14016 28868 14068
rect 31576 14016 31628 14068
rect 31208 13948 31260 14000
rect 32128 13948 32180 14000
rect 24124 13889 24138 13923
rect 24138 13889 24172 13923
rect 24172 13889 24176 13923
rect 24124 13880 24176 13889
rect 24860 13923 24912 13932
rect 24860 13889 24874 13923
rect 24874 13889 24908 13923
rect 24908 13889 24912 13923
rect 24860 13880 24912 13889
rect 25320 13880 25372 13932
rect 25504 13923 25556 13932
rect 25504 13889 25513 13923
rect 25513 13889 25547 13923
rect 25547 13889 25556 13923
rect 25504 13880 25556 13889
rect 25596 13923 25648 13932
rect 25596 13889 25605 13923
rect 25605 13889 25639 13923
rect 25639 13889 25648 13923
rect 25596 13880 25648 13889
rect 24308 13787 24360 13796
rect 24308 13753 24317 13787
rect 24317 13753 24351 13787
rect 24351 13753 24360 13787
rect 24308 13744 24360 13753
rect 18052 13676 18104 13728
rect 18880 13676 18932 13728
rect 25964 13855 26016 13864
rect 25964 13821 25973 13855
rect 25973 13821 26007 13855
rect 26007 13821 26016 13855
rect 25964 13812 26016 13821
rect 26148 13923 26200 13932
rect 26148 13889 26157 13923
rect 26157 13889 26191 13923
rect 26191 13889 26200 13923
rect 26148 13880 26200 13889
rect 27344 13923 27396 13932
rect 27344 13889 27353 13923
rect 27353 13889 27387 13923
rect 27387 13889 27396 13923
rect 27344 13880 27396 13889
rect 27436 13923 27488 13932
rect 27436 13889 27445 13923
rect 27445 13889 27479 13923
rect 27479 13889 27488 13923
rect 27436 13880 27488 13889
rect 27712 13923 27764 13932
rect 27712 13889 27721 13923
rect 27721 13889 27755 13923
rect 27755 13889 27764 13923
rect 27712 13880 27764 13889
rect 27804 13923 27856 13932
rect 27804 13889 27813 13923
rect 27813 13889 27847 13923
rect 27847 13889 27856 13923
rect 27804 13880 27856 13889
rect 28080 13923 28132 13932
rect 28080 13889 28089 13923
rect 28089 13889 28123 13923
rect 28123 13889 28132 13923
rect 28080 13880 28132 13889
rect 32588 14016 32640 14068
rect 32864 14016 32916 14068
rect 36176 14016 36228 14068
rect 39856 14016 39908 14068
rect 32404 13923 32456 13932
rect 32404 13889 32408 13923
rect 32408 13889 32442 13923
rect 32442 13889 32456 13923
rect 26424 13812 26476 13864
rect 27068 13812 27120 13864
rect 32404 13880 32456 13889
rect 29460 13812 29512 13864
rect 29828 13855 29880 13864
rect 29828 13821 29837 13855
rect 29837 13821 29871 13855
rect 29871 13821 29880 13855
rect 29828 13812 29880 13821
rect 31944 13855 31996 13864
rect 31944 13821 31953 13855
rect 31953 13821 31987 13855
rect 31987 13821 31996 13855
rect 31944 13812 31996 13821
rect 33508 13948 33560 14000
rect 33048 13880 33100 13932
rect 33784 13880 33836 13932
rect 34060 13923 34112 13932
rect 34060 13889 34069 13923
rect 34069 13889 34103 13923
rect 34103 13889 34112 13923
rect 34060 13880 34112 13889
rect 34152 13923 34204 13932
rect 34152 13889 34161 13923
rect 34161 13889 34195 13923
rect 34195 13889 34204 13923
rect 34152 13880 34204 13889
rect 36268 13991 36320 14000
rect 36268 13957 36277 13991
rect 36277 13957 36311 13991
rect 36311 13957 36320 13991
rect 36268 13948 36320 13957
rect 36360 13991 36412 14000
rect 36360 13957 36369 13991
rect 36369 13957 36403 13991
rect 36403 13957 36412 13991
rect 36360 13948 36412 13957
rect 39304 13948 39356 14000
rect 39580 13948 39632 14000
rect 25044 13787 25096 13796
rect 25044 13753 25053 13787
rect 25053 13753 25087 13787
rect 25087 13753 25096 13787
rect 25044 13744 25096 13753
rect 25688 13744 25740 13796
rect 30932 13744 30984 13796
rect 33600 13812 33652 13864
rect 35992 13880 36044 13932
rect 36452 13923 36504 13932
rect 36452 13889 36461 13923
rect 36461 13889 36495 13923
rect 36495 13889 36504 13923
rect 36452 13880 36504 13889
rect 38844 13880 38896 13932
rect 40592 13923 40644 13932
rect 40592 13889 40601 13923
rect 40601 13889 40635 13923
rect 40635 13889 40644 13923
rect 40592 13880 40644 13889
rect 45744 14016 45796 14068
rect 46020 14016 46072 14068
rect 44088 13991 44140 14000
rect 44088 13957 44097 13991
rect 44097 13957 44131 13991
rect 44131 13957 44140 13991
rect 44088 13948 44140 13957
rect 46756 14016 46808 14068
rect 46940 14016 46992 14068
rect 47492 14016 47544 14068
rect 47676 14016 47728 14068
rect 47860 13948 47912 14000
rect 48412 13948 48464 14000
rect 36544 13812 36596 13864
rect 26608 13676 26660 13728
rect 26792 13676 26844 13728
rect 27160 13719 27212 13728
rect 27160 13685 27169 13719
rect 27169 13685 27203 13719
rect 27203 13685 27212 13719
rect 27160 13676 27212 13685
rect 27620 13676 27672 13728
rect 34244 13744 34296 13796
rect 36268 13744 36320 13796
rect 46940 13923 46992 13932
rect 46940 13889 46949 13923
rect 46949 13889 46983 13923
rect 46983 13889 46992 13923
rect 46940 13880 46992 13889
rect 49240 13880 49292 13932
rect 51724 14016 51776 14068
rect 52276 14016 52328 14068
rect 54208 14016 54260 14068
rect 51540 13948 51592 14000
rect 52092 13880 52144 13932
rect 52184 13923 52236 13932
rect 52184 13889 52193 13923
rect 52193 13889 52227 13923
rect 52227 13889 52236 13923
rect 52184 13880 52236 13889
rect 53472 13880 53524 13932
rect 54024 13948 54076 14000
rect 33140 13676 33192 13728
rect 33692 13676 33744 13728
rect 36636 13719 36688 13728
rect 36636 13685 36645 13719
rect 36645 13685 36679 13719
rect 36679 13685 36688 13719
rect 36636 13676 36688 13685
rect 39396 13676 39448 13728
rect 40408 13719 40460 13728
rect 40408 13685 40417 13719
rect 40417 13685 40451 13719
rect 40451 13685 40460 13719
rect 40408 13676 40460 13685
rect 42248 13744 42300 13796
rect 41972 13676 42024 13728
rect 46848 13812 46900 13864
rect 50160 13855 50212 13864
rect 50160 13821 50169 13855
rect 50169 13821 50203 13855
rect 50203 13821 50212 13855
rect 50160 13812 50212 13821
rect 50620 13812 50672 13864
rect 50804 13812 50856 13864
rect 51356 13812 51408 13864
rect 54944 13812 54996 13864
rect 55588 13880 55640 13932
rect 47124 13744 47176 13796
rect 47768 13744 47820 13796
rect 49884 13744 49936 13796
rect 51540 13744 51592 13796
rect 52552 13744 52604 13796
rect 45100 13676 45152 13728
rect 45376 13676 45428 13728
rect 46940 13676 46992 13728
rect 51172 13676 51224 13728
rect 51816 13676 51868 13728
rect 52368 13719 52420 13728
rect 52368 13685 52377 13719
rect 52377 13685 52411 13719
rect 52411 13685 52420 13719
rect 52368 13676 52420 13685
rect 53932 13719 53984 13728
rect 53932 13685 53962 13719
rect 53962 13685 53984 13719
rect 53932 13676 53984 13685
rect 55404 13719 55456 13728
rect 55404 13685 55413 13719
rect 55413 13685 55447 13719
rect 55447 13685 55456 13719
rect 55404 13676 55456 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 9404 13336 9456 13388
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 16396 13268 16448 13320
rect 10876 13200 10928 13252
rect 16948 13243 17000 13252
rect 16948 13209 16957 13243
rect 16957 13209 16991 13243
rect 16991 13209 17000 13243
rect 16948 13200 17000 13209
rect 17316 13311 17368 13320
rect 17316 13277 17325 13311
rect 17325 13277 17359 13311
rect 17359 13277 17368 13311
rect 17316 13268 17368 13277
rect 17408 13268 17460 13320
rect 21548 13515 21600 13524
rect 21548 13481 21557 13515
rect 21557 13481 21591 13515
rect 21591 13481 21600 13515
rect 21548 13472 21600 13481
rect 23020 13472 23072 13524
rect 23204 13515 23256 13524
rect 23204 13481 23213 13515
rect 23213 13481 23247 13515
rect 23247 13481 23256 13515
rect 23204 13472 23256 13481
rect 27436 13515 27488 13524
rect 27436 13481 27445 13515
rect 27445 13481 27479 13515
rect 27479 13481 27488 13515
rect 27436 13472 27488 13481
rect 29184 13515 29236 13524
rect 29184 13481 29193 13515
rect 29193 13481 29227 13515
rect 29227 13481 29236 13515
rect 29184 13472 29236 13481
rect 29828 13472 29880 13524
rect 32128 13472 32180 13524
rect 36636 13472 36688 13524
rect 37832 13472 37884 13524
rect 38384 13472 38436 13524
rect 39396 13515 39448 13524
rect 39396 13481 39405 13515
rect 39405 13481 39439 13515
rect 39439 13481 39448 13515
rect 39396 13472 39448 13481
rect 40408 13515 40460 13524
rect 40408 13481 40417 13515
rect 40417 13481 40451 13515
rect 40451 13481 40460 13515
rect 40408 13472 40460 13481
rect 40500 13515 40552 13524
rect 40500 13481 40509 13515
rect 40509 13481 40543 13515
rect 40543 13481 40552 13515
rect 40500 13472 40552 13481
rect 41696 13472 41748 13524
rect 42340 13472 42392 13524
rect 42708 13472 42760 13524
rect 44180 13472 44232 13524
rect 45008 13472 45060 13524
rect 50160 13515 50212 13524
rect 50160 13481 50169 13515
rect 50169 13481 50203 13515
rect 50203 13481 50212 13515
rect 50160 13472 50212 13481
rect 53932 13472 53984 13524
rect 18420 13404 18472 13456
rect 19432 13404 19484 13456
rect 21456 13404 21508 13456
rect 19248 13336 19300 13388
rect 23480 13336 23532 13388
rect 17960 13268 18012 13320
rect 18420 13243 18472 13252
rect 18420 13209 18429 13243
rect 18429 13209 18463 13243
rect 18463 13209 18472 13243
rect 18420 13200 18472 13209
rect 18788 13268 18840 13320
rect 19708 13311 19760 13320
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 23296 13268 23348 13320
rect 25964 13404 26016 13456
rect 26148 13404 26200 13456
rect 24124 13336 24176 13388
rect 24308 13336 24360 13388
rect 26700 13379 26752 13388
rect 26700 13345 26709 13379
rect 26709 13345 26743 13379
rect 26743 13345 26752 13379
rect 26700 13336 26752 13345
rect 26792 13379 26844 13388
rect 26792 13345 26801 13379
rect 26801 13345 26835 13379
rect 26835 13345 26844 13379
rect 26792 13336 26844 13345
rect 27160 13336 27212 13388
rect 32588 13404 32640 13456
rect 27528 13336 27580 13388
rect 27712 13268 27764 13320
rect 28356 13336 28408 13388
rect 13820 13132 13872 13184
rect 18144 13132 18196 13184
rect 19800 13200 19852 13252
rect 22376 13200 22428 13252
rect 19064 13132 19116 13184
rect 20720 13132 20772 13184
rect 21456 13132 21508 13184
rect 25044 13200 25096 13252
rect 27804 13200 27856 13252
rect 27896 13200 27948 13252
rect 24400 13132 24452 13184
rect 26792 13132 26844 13184
rect 28356 13200 28408 13252
rect 28724 13311 28776 13320
rect 28724 13277 28733 13311
rect 28733 13277 28767 13311
rect 28767 13277 28776 13311
rect 28724 13268 28776 13277
rect 30380 13311 30432 13320
rect 30380 13277 30389 13311
rect 30389 13277 30423 13311
rect 30423 13277 30432 13311
rect 30380 13268 30432 13277
rect 34152 13336 34204 13388
rect 31944 13268 31996 13320
rect 30288 13200 30340 13252
rect 31944 13132 31996 13184
rect 35440 13200 35492 13252
rect 36820 13404 36872 13456
rect 39764 13404 39816 13456
rect 40040 13404 40092 13456
rect 40776 13447 40828 13456
rect 40776 13413 40785 13447
rect 40785 13413 40819 13447
rect 40819 13413 40828 13447
rect 40776 13404 40828 13413
rect 42524 13404 42576 13456
rect 44548 13404 44600 13456
rect 44640 13404 44692 13456
rect 36360 13311 36412 13320
rect 36360 13277 36369 13311
rect 36369 13277 36403 13311
rect 36403 13277 36412 13311
rect 36360 13268 36412 13277
rect 36728 13311 36780 13320
rect 36728 13277 36737 13311
rect 36737 13277 36771 13311
rect 36771 13277 36780 13311
rect 36728 13268 36780 13277
rect 37004 13311 37056 13320
rect 37004 13277 37013 13311
rect 37013 13277 37047 13311
rect 37047 13277 37056 13311
rect 37004 13268 37056 13277
rect 37832 13268 37884 13320
rect 38200 13311 38252 13320
rect 38200 13277 38210 13311
rect 38210 13277 38244 13311
rect 38244 13277 38252 13311
rect 38200 13268 38252 13277
rect 38384 13311 38436 13320
rect 38384 13277 38393 13311
rect 38393 13277 38427 13311
rect 38427 13277 38436 13311
rect 38384 13268 38436 13277
rect 34704 13132 34756 13184
rect 36544 13132 36596 13184
rect 37096 13200 37148 13252
rect 38016 13200 38068 13252
rect 38292 13132 38344 13184
rect 39120 13311 39172 13320
rect 39120 13277 39129 13311
rect 39129 13277 39163 13311
rect 39163 13277 39172 13311
rect 39120 13268 39172 13277
rect 41512 13336 41564 13388
rect 51172 13404 51224 13456
rect 52368 13404 52420 13456
rect 39856 13311 39908 13320
rect 39856 13277 39865 13311
rect 39865 13277 39899 13311
rect 39899 13277 39908 13311
rect 39856 13268 39908 13277
rect 40040 13311 40092 13320
rect 40040 13277 40049 13311
rect 40049 13277 40083 13311
rect 40083 13277 40092 13311
rect 40040 13268 40092 13277
rect 40500 13268 40552 13320
rect 40776 13268 40828 13320
rect 41696 13268 41748 13320
rect 42892 13268 42944 13320
rect 44456 13311 44508 13320
rect 44456 13277 44465 13311
rect 44465 13277 44499 13311
rect 44499 13277 44508 13311
rect 44456 13268 44508 13277
rect 44916 13268 44968 13320
rect 40132 13243 40184 13252
rect 40132 13209 40141 13243
rect 40141 13209 40175 13243
rect 40175 13209 40184 13243
rect 40132 13200 40184 13209
rect 45284 13311 45336 13320
rect 45284 13277 45293 13311
rect 45293 13277 45327 13311
rect 45327 13277 45336 13311
rect 45284 13268 45336 13277
rect 48044 13336 48096 13388
rect 50252 13336 50304 13388
rect 47768 13268 47820 13320
rect 53840 13336 53892 13388
rect 55404 13336 55456 13388
rect 50620 13268 50672 13320
rect 54116 13268 54168 13320
rect 45376 13243 45428 13252
rect 40408 13132 40460 13184
rect 42984 13132 43036 13184
rect 45376 13209 45385 13243
rect 45385 13209 45419 13243
rect 45419 13209 45428 13243
rect 45376 13200 45428 13209
rect 44640 13175 44692 13184
rect 44640 13141 44649 13175
rect 44649 13141 44683 13175
rect 44683 13141 44692 13175
rect 44640 13132 44692 13141
rect 45560 13132 45612 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 66314 13030 66366 13082
rect 66378 13030 66430 13082
rect 66442 13030 66494 13082
rect 66506 13030 66558 13082
rect 66570 13030 66622 13082
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 14464 12928 14516 12980
rect 18420 12928 18472 12980
rect 19156 12928 19208 12980
rect 18512 12860 18564 12912
rect 17316 12792 17368 12844
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 18420 12792 18472 12844
rect 22192 12971 22244 12980
rect 22192 12937 22201 12971
rect 22201 12937 22235 12971
rect 22235 12937 22244 12971
rect 22192 12928 22244 12937
rect 22376 12928 22428 12980
rect 23940 12928 23992 12980
rect 25044 12928 25096 12980
rect 25504 12928 25556 12980
rect 27896 12928 27948 12980
rect 28540 12928 28592 12980
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 18880 12792 18932 12801
rect 19064 12835 19116 12844
rect 19064 12801 19073 12835
rect 19073 12801 19107 12835
rect 19107 12801 19116 12835
rect 19064 12792 19116 12801
rect 14832 12724 14884 12776
rect 16948 12724 17000 12776
rect 15016 12656 15068 12708
rect 16396 12656 16448 12708
rect 19800 12835 19852 12844
rect 19800 12801 19809 12835
rect 19809 12801 19843 12835
rect 19843 12801 19852 12835
rect 19800 12792 19852 12801
rect 21456 12860 21508 12912
rect 20076 12835 20128 12844
rect 20076 12801 20085 12835
rect 20085 12801 20119 12835
rect 20119 12801 20128 12835
rect 20076 12792 20128 12801
rect 21548 12792 21600 12844
rect 25228 12792 25280 12844
rect 26700 12860 26752 12912
rect 31668 12928 31720 12980
rect 32312 12928 32364 12980
rect 33324 12928 33376 12980
rect 19340 12656 19392 12708
rect 20720 12656 20772 12708
rect 23940 12724 23992 12776
rect 25688 12835 25740 12844
rect 25688 12801 25697 12835
rect 25697 12801 25731 12835
rect 25731 12801 25740 12835
rect 25688 12792 25740 12801
rect 25780 12835 25832 12844
rect 25780 12801 25789 12835
rect 25789 12801 25823 12835
rect 25823 12801 25832 12835
rect 25780 12792 25832 12801
rect 26976 12656 27028 12708
rect 27896 12656 27948 12708
rect 32036 12792 32088 12844
rect 32772 12792 32824 12844
rect 33876 12860 33928 12912
rect 34704 12903 34756 12912
rect 34704 12869 34713 12903
rect 34713 12869 34747 12903
rect 34747 12869 34756 12903
rect 34704 12860 34756 12869
rect 34796 12860 34848 12912
rect 36912 12928 36964 12980
rect 37004 12928 37056 12980
rect 37832 12971 37884 12980
rect 37832 12937 37841 12971
rect 37841 12937 37875 12971
rect 37875 12937 37884 12971
rect 37832 12928 37884 12937
rect 37924 12928 37976 12980
rect 38292 12928 38344 12980
rect 36360 12860 36412 12912
rect 33600 12835 33652 12844
rect 33600 12801 33609 12835
rect 33609 12801 33643 12835
rect 33643 12801 33652 12835
rect 33600 12792 33652 12801
rect 36820 12792 36872 12844
rect 37096 12792 37148 12844
rect 37464 12903 37516 12912
rect 37464 12869 37473 12903
rect 37473 12869 37507 12903
rect 37507 12869 37516 12903
rect 37464 12860 37516 12869
rect 37740 12860 37792 12912
rect 37648 12835 37700 12844
rect 37648 12801 37657 12835
rect 37657 12801 37691 12835
rect 37691 12801 37700 12835
rect 38108 12860 38160 12912
rect 40132 12860 40184 12912
rect 37648 12792 37700 12801
rect 38292 12792 38344 12844
rect 38568 12792 38620 12844
rect 32864 12656 32916 12708
rect 34428 12767 34480 12776
rect 34428 12733 34437 12767
rect 34437 12733 34471 12767
rect 34471 12733 34480 12767
rect 34428 12724 34480 12733
rect 35716 12656 35768 12708
rect 39856 12724 39908 12776
rect 40592 12835 40644 12844
rect 40592 12801 40601 12835
rect 40601 12801 40635 12835
rect 40635 12801 40644 12835
rect 40592 12792 40644 12801
rect 41420 12792 41472 12844
rect 42248 12792 42300 12844
rect 38200 12656 38252 12708
rect 42156 12724 42208 12776
rect 45100 12928 45152 12980
rect 42984 12903 43036 12912
rect 42984 12869 42993 12903
rect 42993 12869 43027 12903
rect 43027 12869 43036 12903
rect 42984 12860 43036 12869
rect 44272 12860 44324 12912
rect 46756 12860 46808 12912
rect 44548 12792 44600 12844
rect 45100 12835 45152 12844
rect 45100 12801 45109 12835
rect 45109 12801 45143 12835
rect 45143 12801 45152 12835
rect 45100 12792 45152 12801
rect 50344 12792 50396 12844
rect 54484 12792 54536 12844
rect 44456 12767 44508 12776
rect 44456 12733 44465 12767
rect 44465 12733 44499 12767
rect 44499 12733 44508 12767
rect 44456 12724 44508 12733
rect 45376 12767 45428 12776
rect 45376 12733 45385 12767
rect 45385 12733 45419 12767
rect 45419 12733 45428 12767
rect 45376 12724 45428 12733
rect 44272 12656 44324 12708
rect 44916 12656 44968 12708
rect 12992 12588 13044 12640
rect 17684 12631 17736 12640
rect 17684 12597 17693 12631
rect 17693 12597 17727 12631
rect 17727 12597 17736 12631
rect 17684 12588 17736 12597
rect 18420 12588 18472 12640
rect 19248 12588 19300 12640
rect 21180 12588 21232 12640
rect 27344 12588 27396 12640
rect 31024 12588 31076 12640
rect 31484 12631 31536 12640
rect 31484 12597 31493 12631
rect 31493 12597 31527 12631
rect 31527 12597 31536 12631
rect 31484 12588 31536 12597
rect 33416 12588 33468 12640
rect 36360 12588 36412 12640
rect 40684 12588 40736 12640
rect 46848 12631 46900 12640
rect 46848 12597 46857 12631
rect 46857 12597 46891 12631
rect 46891 12597 46900 12631
rect 46848 12588 46900 12597
rect 50988 12631 51040 12640
rect 50988 12597 50997 12631
rect 50997 12597 51031 12631
rect 51031 12597 51040 12631
rect 50988 12588 51040 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 14004 12384 14056 12436
rect 17316 12384 17368 12436
rect 20076 12384 20128 12436
rect 24216 12384 24268 12436
rect 24308 12384 24360 12436
rect 25780 12384 25832 12436
rect 12716 12248 12768 12300
rect 17132 12248 17184 12300
rect 18328 12316 18380 12368
rect 19340 12248 19392 12300
rect 14924 12180 14976 12232
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 17960 12180 18012 12232
rect 18052 12180 18104 12232
rect 19156 12180 19208 12232
rect 19432 12180 19484 12232
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 21456 12248 21508 12300
rect 24584 12316 24636 12368
rect 17500 12112 17552 12164
rect 17408 12044 17460 12096
rect 20536 12044 20588 12096
rect 23296 12087 23348 12096
rect 23296 12053 23305 12087
rect 23305 12053 23339 12087
rect 23339 12053 23348 12087
rect 23296 12044 23348 12053
rect 23388 12044 23440 12096
rect 24032 12180 24084 12232
rect 24124 12223 24176 12232
rect 24124 12189 24133 12223
rect 24133 12189 24167 12223
rect 24167 12189 24176 12223
rect 24124 12180 24176 12189
rect 24308 12180 24360 12232
rect 25044 12291 25096 12300
rect 25044 12257 25053 12291
rect 25053 12257 25087 12291
rect 25087 12257 25096 12291
rect 25044 12248 25096 12257
rect 25228 12248 25280 12300
rect 25780 12180 25832 12232
rect 28540 12384 28592 12436
rect 32864 12427 32916 12436
rect 32864 12393 32873 12427
rect 32873 12393 32907 12427
rect 32907 12393 32916 12427
rect 32864 12384 32916 12393
rect 26148 12316 26200 12368
rect 26700 12248 26752 12300
rect 27712 12316 27764 12368
rect 32772 12316 32824 12368
rect 34520 12384 34572 12436
rect 35440 12384 35492 12436
rect 35992 12384 36044 12436
rect 26148 12223 26200 12232
rect 26148 12189 26157 12223
rect 26157 12189 26191 12223
rect 26191 12189 26200 12223
rect 26148 12180 26200 12189
rect 26240 12223 26292 12232
rect 26240 12189 26249 12223
rect 26249 12189 26283 12223
rect 26283 12189 26292 12223
rect 26240 12180 26292 12189
rect 27712 12223 27764 12232
rect 27712 12189 27721 12223
rect 27721 12189 27755 12223
rect 27755 12189 27764 12223
rect 27712 12180 27764 12189
rect 27896 12223 27948 12232
rect 27896 12189 27905 12223
rect 27905 12189 27939 12223
rect 27939 12189 27948 12223
rect 27896 12180 27948 12189
rect 27988 12223 28040 12232
rect 27988 12189 27997 12223
rect 27997 12189 28031 12223
rect 28031 12189 28040 12223
rect 27988 12180 28040 12189
rect 28264 12180 28316 12232
rect 28632 12248 28684 12300
rect 31484 12248 31536 12300
rect 24216 12112 24268 12164
rect 28172 12112 28224 12164
rect 29460 12180 29512 12232
rect 33232 12316 33284 12368
rect 34244 12316 34296 12368
rect 33600 12248 33652 12300
rect 24032 12044 24084 12096
rect 25872 12044 25924 12096
rect 26608 12044 26660 12096
rect 27068 12087 27120 12096
rect 27068 12053 27077 12087
rect 27077 12053 27111 12087
rect 27111 12053 27120 12087
rect 27068 12044 27120 12053
rect 27896 12044 27948 12096
rect 31852 12112 31904 12164
rect 32864 12112 32916 12164
rect 33416 12223 33468 12232
rect 33416 12189 33425 12223
rect 33425 12189 33459 12223
rect 33459 12189 33468 12223
rect 33416 12180 33468 12189
rect 33508 12223 33560 12232
rect 33508 12189 33522 12223
rect 33522 12189 33556 12223
rect 33556 12189 33560 12223
rect 33508 12180 33560 12189
rect 29828 12044 29880 12096
rect 34152 12223 34204 12232
rect 34152 12189 34161 12223
rect 34161 12189 34195 12223
rect 34195 12189 34204 12223
rect 34152 12180 34204 12189
rect 34244 12223 34296 12232
rect 34244 12189 34253 12223
rect 34253 12189 34287 12223
rect 34287 12189 34296 12223
rect 34244 12180 34296 12189
rect 35716 12316 35768 12368
rect 36636 12316 36688 12368
rect 37372 12316 37424 12368
rect 35348 12248 35400 12300
rect 37556 12248 37608 12300
rect 42156 12427 42208 12436
rect 42156 12393 42165 12427
rect 42165 12393 42199 12427
rect 42199 12393 42208 12427
rect 42156 12384 42208 12393
rect 42892 12427 42944 12436
rect 42892 12393 42901 12427
rect 42901 12393 42935 12427
rect 42935 12393 42944 12427
rect 42892 12384 42944 12393
rect 44548 12384 44600 12436
rect 45376 12384 45428 12436
rect 40684 12291 40736 12300
rect 40684 12257 40693 12291
rect 40693 12257 40727 12291
rect 40727 12257 40736 12291
rect 40684 12248 40736 12257
rect 42156 12248 42208 12300
rect 42800 12316 42852 12368
rect 34520 12112 34572 12164
rect 37280 12223 37332 12232
rect 37280 12189 37289 12223
rect 37289 12189 37323 12223
rect 37323 12189 37332 12223
rect 37280 12180 37332 12189
rect 33968 12044 34020 12096
rect 35992 12112 36044 12164
rect 37832 12223 37884 12232
rect 37832 12189 37842 12223
rect 37842 12189 37876 12223
rect 37876 12189 37884 12223
rect 37832 12180 37884 12189
rect 38108 12223 38160 12232
rect 38108 12189 38117 12223
rect 38117 12189 38151 12223
rect 38151 12189 38160 12223
rect 38108 12180 38160 12189
rect 38476 12180 38528 12232
rect 40224 12180 40276 12232
rect 44180 12316 44232 12368
rect 46940 12384 46992 12436
rect 50344 12384 50396 12436
rect 46848 12248 46900 12300
rect 51816 12248 51868 12300
rect 54024 12248 54076 12300
rect 54208 12248 54260 12300
rect 39120 12112 39172 12164
rect 38108 12044 38160 12096
rect 38384 12087 38436 12096
rect 38384 12053 38393 12087
rect 38393 12053 38427 12087
rect 38427 12053 38436 12087
rect 38384 12044 38436 12053
rect 42524 12155 42576 12164
rect 42524 12121 42533 12155
rect 42533 12121 42567 12155
rect 42567 12121 42576 12155
rect 42524 12112 42576 12121
rect 43628 12180 43680 12232
rect 45560 12180 45612 12232
rect 47124 12223 47176 12232
rect 47124 12189 47133 12223
rect 47133 12189 47167 12223
rect 47167 12189 47176 12223
rect 47124 12180 47176 12189
rect 55404 12223 55456 12232
rect 55404 12189 55413 12223
rect 55413 12189 55447 12223
rect 55447 12189 55456 12223
rect 55404 12180 55456 12189
rect 47676 12112 47728 12164
rect 49240 12112 49292 12164
rect 50344 12112 50396 12164
rect 50712 12112 50764 12164
rect 44272 12044 44324 12096
rect 48320 12044 48372 12096
rect 51540 12044 51592 12096
rect 52276 12044 52328 12096
rect 52644 12112 52696 12164
rect 55864 12112 55916 12164
rect 54116 12044 54168 12096
rect 54944 12044 54996 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 66314 11942 66366 11994
rect 66378 11942 66430 11994
rect 66442 11942 66494 11994
rect 66506 11942 66558 11994
rect 66570 11942 66622 11994
rect 14832 11840 14884 11892
rect 15568 11840 15620 11892
rect 12992 11815 13044 11824
rect 12992 11781 13001 11815
rect 13001 11781 13035 11815
rect 13035 11781 13044 11815
rect 12992 11772 13044 11781
rect 14004 11772 14056 11824
rect 18880 11840 18932 11892
rect 17408 11815 17460 11824
rect 17408 11781 17417 11815
rect 17417 11781 17451 11815
rect 17451 11781 17460 11815
rect 17408 11772 17460 11781
rect 18144 11772 18196 11824
rect 22192 11772 22244 11824
rect 12716 11747 12768 11756
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 12716 11704 12768 11713
rect 16948 11704 17000 11756
rect 17684 11747 17736 11756
rect 17684 11713 17693 11747
rect 17693 11713 17727 11747
rect 17727 11713 17736 11747
rect 17684 11704 17736 11713
rect 21180 11704 21232 11756
rect 22652 11747 22704 11756
rect 22652 11713 22661 11747
rect 22661 11713 22695 11747
rect 22695 11713 22704 11747
rect 22652 11704 22704 11713
rect 22928 11704 22980 11756
rect 23388 11772 23440 11824
rect 24124 11840 24176 11892
rect 23296 11747 23348 11756
rect 23296 11713 23305 11747
rect 23305 11713 23339 11747
rect 23339 11713 23348 11747
rect 23296 11704 23348 11713
rect 20536 11636 20588 11688
rect 23664 11747 23716 11756
rect 23664 11713 23673 11747
rect 23673 11713 23707 11747
rect 23707 11713 23716 11747
rect 23664 11704 23716 11713
rect 22928 11568 22980 11620
rect 23296 11568 23348 11620
rect 24952 11772 25004 11824
rect 25872 11772 25924 11824
rect 26240 11772 26292 11824
rect 27988 11772 28040 11824
rect 23940 11747 23992 11756
rect 23940 11713 23949 11747
rect 23949 11713 23983 11747
rect 23983 11713 23992 11747
rect 23940 11704 23992 11713
rect 24308 11747 24360 11756
rect 24308 11713 24317 11747
rect 24317 11713 24351 11747
rect 24351 11713 24360 11747
rect 24308 11704 24360 11713
rect 24492 11747 24544 11756
rect 24492 11713 24501 11747
rect 24501 11713 24535 11747
rect 24535 11713 24544 11747
rect 24492 11704 24544 11713
rect 25228 11747 25280 11756
rect 25228 11713 25237 11747
rect 25237 11713 25271 11747
rect 25271 11713 25280 11747
rect 25228 11704 25280 11713
rect 25320 11704 25372 11756
rect 24216 11679 24268 11688
rect 24216 11645 24225 11679
rect 24225 11645 24259 11679
rect 24259 11645 24268 11679
rect 24216 11636 24268 11645
rect 24584 11636 24636 11688
rect 25872 11679 25924 11688
rect 25872 11645 25881 11679
rect 25881 11645 25915 11679
rect 25915 11645 25924 11679
rect 25872 11636 25924 11645
rect 26056 11636 26108 11688
rect 26516 11636 26568 11688
rect 27528 11747 27580 11756
rect 27528 11713 27537 11747
rect 27537 11713 27571 11747
rect 27571 11713 27580 11747
rect 27528 11704 27580 11713
rect 27620 11747 27672 11756
rect 27620 11713 27629 11747
rect 27629 11713 27663 11747
rect 27663 11713 27672 11747
rect 27620 11704 27672 11713
rect 27712 11747 27764 11756
rect 27712 11713 27721 11747
rect 27721 11713 27755 11747
rect 27755 11713 27764 11747
rect 27712 11704 27764 11713
rect 31852 11772 31904 11824
rect 32128 11772 32180 11824
rect 34796 11840 34848 11892
rect 36544 11840 36596 11892
rect 37096 11840 37148 11892
rect 37464 11840 37516 11892
rect 33968 11815 34020 11824
rect 33968 11781 33977 11815
rect 33977 11781 34011 11815
rect 34011 11781 34020 11815
rect 33968 11772 34020 11781
rect 29460 11747 29512 11756
rect 29460 11713 29469 11747
rect 29469 11713 29503 11747
rect 29503 11713 29512 11747
rect 29460 11704 29512 11713
rect 34520 11704 34572 11756
rect 29736 11679 29788 11688
rect 29736 11645 29745 11679
rect 29745 11645 29779 11679
rect 29779 11645 29788 11679
rect 29736 11636 29788 11645
rect 31392 11636 31444 11688
rect 36636 11747 36688 11756
rect 36636 11713 36640 11747
rect 36640 11713 36674 11747
rect 36674 11713 36688 11747
rect 36636 11704 36688 11713
rect 36544 11636 36596 11688
rect 36912 11747 36964 11756
rect 37556 11772 37608 11824
rect 38476 11772 38528 11824
rect 36912 11713 36957 11747
rect 36957 11713 36964 11747
rect 36912 11704 36964 11713
rect 37832 11747 37884 11756
rect 37832 11713 37841 11747
rect 37841 11713 37875 11747
rect 37875 11713 37884 11747
rect 37832 11704 37884 11713
rect 38384 11747 38436 11756
rect 38384 11713 38393 11747
rect 38393 11713 38427 11747
rect 38427 11713 38436 11747
rect 38384 11704 38436 11713
rect 39488 11704 39540 11756
rect 17960 11500 18012 11552
rect 18696 11500 18748 11552
rect 23388 11543 23440 11552
rect 23388 11509 23397 11543
rect 23397 11509 23431 11543
rect 23431 11509 23440 11543
rect 23388 11500 23440 11509
rect 24124 11543 24176 11552
rect 24124 11509 24133 11543
rect 24133 11509 24167 11543
rect 24167 11509 24176 11543
rect 24124 11500 24176 11509
rect 25872 11500 25924 11552
rect 28264 11568 28316 11620
rect 26424 11543 26476 11552
rect 26424 11509 26433 11543
rect 26433 11509 26467 11543
rect 26467 11509 26476 11543
rect 26424 11500 26476 11509
rect 27252 11543 27304 11552
rect 27252 11509 27261 11543
rect 27261 11509 27295 11543
rect 27295 11509 27304 11543
rect 27252 11500 27304 11509
rect 31208 11543 31260 11552
rect 31208 11509 31217 11543
rect 31217 11509 31251 11543
rect 31251 11509 31260 11543
rect 31208 11500 31260 11509
rect 31668 11500 31720 11552
rect 33232 11500 33284 11552
rect 33600 11500 33652 11552
rect 34428 11500 34480 11552
rect 36544 11500 36596 11552
rect 37280 11679 37332 11688
rect 37280 11645 37289 11679
rect 37289 11645 37323 11679
rect 37323 11645 37332 11679
rect 37280 11636 37332 11645
rect 37096 11568 37148 11620
rect 39672 11568 39724 11620
rect 38108 11500 38160 11552
rect 38200 11543 38252 11552
rect 38200 11509 38209 11543
rect 38209 11509 38243 11543
rect 38243 11509 38252 11543
rect 38200 11500 38252 11509
rect 38568 11543 38620 11552
rect 38568 11509 38577 11543
rect 38577 11509 38611 11543
rect 38611 11509 38620 11543
rect 38568 11500 38620 11509
rect 40592 11840 40644 11892
rect 47676 11883 47728 11892
rect 47676 11849 47685 11883
rect 47685 11849 47719 11883
rect 47719 11849 47728 11883
rect 47676 11840 47728 11849
rect 47952 11840 48004 11892
rect 42524 11772 42576 11824
rect 45836 11772 45888 11824
rect 50712 11883 50764 11892
rect 50712 11849 50721 11883
rect 50721 11849 50755 11883
rect 50755 11849 50764 11883
rect 50712 11840 50764 11849
rect 50988 11840 51040 11892
rect 47860 11747 47912 11756
rect 47860 11713 47869 11747
rect 47869 11713 47903 11747
rect 47903 11713 47912 11747
rect 47860 11704 47912 11713
rect 47952 11747 48004 11756
rect 47952 11713 47961 11747
rect 47961 11713 47995 11747
rect 47995 11713 48004 11747
rect 47952 11704 48004 11713
rect 48504 11747 48556 11756
rect 48504 11713 48513 11747
rect 48513 11713 48547 11747
rect 48547 11713 48556 11747
rect 48504 11704 48556 11713
rect 48596 11747 48648 11756
rect 48596 11713 48605 11747
rect 48605 11713 48639 11747
rect 48639 11713 48648 11747
rect 48596 11704 48648 11713
rect 48872 11747 48924 11756
rect 48872 11713 48881 11747
rect 48881 11713 48915 11747
rect 48915 11713 48924 11747
rect 48872 11704 48924 11713
rect 48320 11636 48372 11688
rect 40132 11568 40184 11620
rect 46572 11568 46624 11620
rect 49332 11747 49384 11756
rect 49332 11713 49341 11747
rect 49341 11713 49375 11747
rect 49375 11713 49384 11747
rect 49332 11704 49384 11713
rect 49700 11704 49752 11756
rect 49976 11704 50028 11756
rect 52828 11772 52880 11824
rect 54392 11772 54444 11824
rect 54944 11772 54996 11824
rect 50988 11747 51040 11756
rect 50988 11713 50997 11747
rect 50997 11713 51031 11747
rect 51031 11713 51040 11747
rect 50988 11704 51040 11713
rect 52000 11704 52052 11756
rect 52276 11747 52328 11756
rect 52276 11713 52285 11747
rect 52285 11713 52319 11747
rect 52319 11713 52328 11747
rect 52276 11704 52328 11713
rect 53012 11747 53064 11756
rect 53012 11713 53021 11747
rect 53021 11713 53055 11747
rect 53055 11713 53064 11747
rect 53012 11704 53064 11713
rect 54208 11747 54260 11756
rect 54208 11713 54217 11747
rect 54217 11713 54251 11747
rect 54251 11713 54260 11747
rect 54208 11704 54260 11713
rect 49884 11679 49936 11688
rect 49884 11645 49893 11679
rect 49893 11645 49927 11679
rect 49927 11645 49936 11679
rect 49884 11636 49936 11645
rect 41696 11500 41748 11552
rect 46940 11500 46992 11552
rect 48136 11543 48188 11552
rect 48136 11509 48145 11543
rect 48145 11509 48179 11543
rect 48179 11509 48188 11543
rect 48136 11500 48188 11509
rect 52000 11568 52052 11620
rect 54484 11679 54536 11688
rect 54484 11645 54493 11679
rect 54493 11645 54527 11679
rect 54527 11645 54536 11679
rect 54484 11636 54536 11645
rect 51080 11500 51132 11552
rect 51172 11543 51224 11552
rect 51172 11509 51181 11543
rect 51181 11509 51215 11543
rect 51215 11509 51224 11543
rect 51172 11500 51224 11509
rect 51908 11500 51960 11552
rect 52460 11543 52512 11552
rect 52460 11509 52469 11543
rect 52469 11509 52503 11543
rect 52503 11509 52512 11543
rect 52460 11500 52512 11509
rect 55036 11500 55088 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 19156 11296 19208 11348
rect 22468 11296 22520 11348
rect 23388 11296 23440 11348
rect 24400 11296 24452 11348
rect 24032 11228 24084 11280
rect 26148 11296 26200 11348
rect 27804 11339 27856 11348
rect 27804 11305 27813 11339
rect 27813 11305 27847 11339
rect 27847 11305 27856 11339
rect 27804 11296 27856 11305
rect 29736 11339 29788 11348
rect 29736 11305 29745 11339
rect 29745 11305 29779 11339
rect 29779 11305 29788 11339
rect 29736 11296 29788 11305
rect 29828 11296 29880 11348
rect 41788 11296 41840 11348
rect 42248 11339 42300 11348
rect 42248 11305 42257 11339
rect 42257 11305 42291 11339
rect 42291 11305 42300 11339
rect 42248 11296 42300 11305
rect 44180 11296 44232 11348
rect 45652 11339 45704 11348
rect 45652 11305 45661 11339
rect 45661 11305 45695 11339
rect 45695 11305 45704 11339
rect 45652 11296 45704 11305
rect 46296 11296 46348 11348
rect 48320 11339 48372 11348
rect 48320 11305 48329 11339
rect 48329 11305 48363 11339
rect 48363 11305 48372 11339
rect 48320 11296 48372 11305
rect 49700 11296 49752 11348
rect 50988 11296 51040 11348
rect 17132 11203 17184 11212
rect 17132 11169 17141 11203
rect 17141 11169 17175 11203
rect 17175 11169 17184 11203
rect 17132 11160 17184 11169
rect 20536 11160 20588 11212
rect 21456 11160 21508 11212
rect 22928 11160 22980 11212
rect 24124 11160 24176 11212
rect 27620 11160 27672 11212
rect 27896 11203 27948 11212
rect 27896 11169 27905 11203
rect 27905 11169 27939 11203
rect 27939 11169 27948 11203
rect 27896 11160 27948 11169
rect 29460 11160 29512 11212
rect 30288 11203 30340 11212
rect 30288 11169 30297 11203
rect 30297 11169 30331 11203
rect 30331 11169 30340 11203
rect 30288 11160 30340 11169
rect 22008 11092 22060 11144
rect 18696 11024 18748 11076
rect 19248 11024 19300 11076
rect 20904 11067 20956 11076
rect 20904 11033 20913 11067
rect 20913 11033 20947 11067
rect 20947 11033 20956 11067
rect 20904 11024 20956 11033
rect 24492 11092 24544 11144
rect 26240 11092 26292 11144
rect 20720 10956 20772 11008
rect 23296 11067 23348 11076
rect 23296 11033 23321 11067
rect 23321 11033 23348 11067
rect 23296 11024 23348 11033
rect 22652 10956 22704 11008
rect 24216 11024 24268 11076
rect 26424 11135 26476 11144
rect 26424 11101 26433 11135
rect 26433 11101 26467 11135
rect 26467 11101 26476 11135
rect 26424 11092 26476 11101
rect 26608 11135 26660 11144
rect 26608 11101 26617 11135
rect 26617 11101 26651 11135
rect 26651 11101 26660 11135
rect 26608 11092 26660 11101
rect 27344 11092 27396 11144
rect 28172 11092 28224 11144
rect 26516 11024 26568 11076
rect 27252 11024 27304 11076
rect 28448 11067 28500 11076
rect 28448 11033 28457 11067
rect 28457 11033 28491 11067
rect 28491 11033 28500 11067
rect 28448 11024 28500 11033
rect 31208 11092 31260 11144
rect 26056 10956 26108 11008
rect 28172 10999 28224 11008
rect 28172 10965 28181 10999
rect 28181 10965 28215 10999
rect 28215 10965 28224 10999
rect 28172 10956 28224 10965
rect 28632 10999 28684 11008
rect 28632 10965 28641 10999
rect 28641 10965 28675 10999
rect 28675 10965 28684 10999
rect 28632 10956 28684 10965
rect 37832 11228 37884 11280
rect 39672 11271 39724 11280
rect 39672 11237 39681 11271
rect 39681 11237 39715 11271
rect 39715 11237 39724 11271
rect 39672 11228 39724 11237
rect 34428 11160 34480 11212
rect 37648 11160 37700 11212
rect 38200 11203 38252 11212
rect 38200 11169 38209 11203
rect 38209 11169 38243 11203
rect 38243 11169 38252 11203
rect 38200 11160 38252 11169
rect 41788 11160 41840 11212
rect 42064 11135 42116 11144
rect 42064 11101 42073 11135
rect 42073 11101 42107 11135
rect 42107 11101 42116 11135
rect 42064 11092 42116 11101
rect 43352 11092 43404 11144
rect 35992 11067 36044 11076
rect 35992 11033 36001 11067
rect 36001 11033 36035 11067
rect 36035 11033 36044 11067
rect 35992 11024 36044 11033
rect 37464 10956 37516 11008
rect 38660 11024 38712 11076
rect 44180 11135 44232 11144
rect 44180 11101 44189 11135
rect 44189 11101 44223 11135
rect 44223 11101 44232 11135
rect 44180 11092 44232 11101
rect 47860 11160 47912 11212
rect 48504 11160 48556 11212
rect 50436 11160 50488 11212
rect 44824 11092 44876 11144
rect 46572 11092 46624 11144
rect 48596 11135 48648 11144
rect 48596 11101 48605 11135
rect 48605 11101 48639 11135
rect 48639 11101 48648 11135
rect 48596 11092 48648 11101
rect 50620 11160 50672 11212
rect 50896 11160 50948 11212
rect 54484 11339 54536 11348
rect 54484 11305 54493 11339
rect 54493 11305 54527 11339
rect 54527 11305 54536 11339
rect 54484 11296 54536 11305
rect 54576 11228 54628 11280
rect 45652 11024 45704 11076
rect 48780 11067 48832 11076
rect 48780 11033 48789 11067
rect 48789 11033 48823 11067
rect 48823 11033 48832 11067
rect 48780 11024 48832 11033
rect 49332 11024 49384 11076
rect 50896 11024 50948 11076
rect 52000 11135 52052 11144
rect 52000 11101 52009 11135
rect 52009 11101 52043 11135
rect 52043 11101 52052 11135
rect 52000 11092 52052 11101
rect 51724 11024 51776 11076
rect 39028 10956 39080 11008
rect 41972 10956 42024 11008
rect 42248 10956 42300 11008
rect 44272 10956 44324 11008
rect 45744 10956 45796 11008
rect 46112 10956 46164 11008
rect 50712 10956 50764 11008
rect 52644 11135 52696 11144
rect 52644 11101 52653 11135
rect 52653 11101 52687 11135
rect 52687 11101 52696 11135
rect 52644 11092 52696 11101
rect 52828 11135 52880 11144
rect 52828 11101 52837 11135
rect 52837 11101 52871 11135
rect 52871 11101 52880 11135
rect 52828 11092 52880 11101
rect 53564 11160 53616 11212
rect 54208 11203 54260 11212
rect 54208 11169 54217 11203
rect 54217 11169 54251 11203
rect 54251 11169 54260 11203
rect 54208 11160 54260 11169
rect 55772 11296 55824 11348
rect 54392 11092 54444 11144
rect 53012 11024 53064 11076
rect 54300 11024 54352 11076
rect 54760 11135 54812 11144
rect 54760 11101 54769 11135
rect 54769 11101 54803 11135
rect 54803 11101 54812 11135
rect 54760 11092 54812 11101
rect 55036 11135 55088 11144
rect 55036 11101 55045 11135
rect 55045 11101 55079 11135
rect 55079 11101 55088 11135
rect 55036 11092 55088 11101
rect 54944 11024 54996 11076
rect 55036 10956 55088 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 66314 10854 66366 10906
rect 66378 10854 66430 10906
rect 66442 10854 66494 10906
rect 66506 10854 66558 10906
rect 66570 10854 66622 10906
rect 19156 10752 19208 10804
rect 19892 10752 19944 10804
rect 22008 10684 22060 10736
rect 17132 10616 17184 10668
rect 19248 10616 19300 10668
rect 19708 10616 19760 10668
rect 25780 10616 25832 10668
rect 26332 10659 26384 10668
rect 26332 10625 26341 10659
rect 26341 10625 26375 10659
rect 26375 10625 26384 10659
rect 26332 10616 26384 10625
rect 26976 10684 27028 10736
rect 32956 10752 33008 10804
rect 35992 10752 36044 10804
rect 38844 10752 38896 10804
rect 39580 10752 39632 10804
rect 42064 10795 42116 10804
rect 42064 10761 42073 10795
rect 42073 10761 42107 10795
rect 42107 10761 42116 10795
rect 42064 10752 42116 10761
rect 44180 10752 44232 10804
rect 45652 10752 45704 10804
rect 33784 10684 33836 10736
rect 34428 10684 34480 10736
rect 28632 10659 28684 10668
rect 28632 10625 28641 10659
rect 28641 10625 28675 10659
rect 28675 10625 28684 10659
rect 28632 10616 28684 10625
rect 29460 10616 29512 10668
rect 29552 10659 29604 10668
rect 29552 10625 29561 10659
rect 29561 10625 29595 10659
rect 29595 10625 29604 10659
rect 29552 10616 29604 10625
rect 32956 10659 33008 10668
rect 32956 10625 32965 10659
rect 32965 10625 32999 10659
rect 32999 10625 33008 10659
rect 32956 10616 33008 10625
rect 20720 10548 20772 10600
rect 21180 10591 21232 10600
rect 21180 10557 21189 10591
rect 21189 10557 21223 10591
rect 21223 10557 21232 10591
rect 21180 10548 21232 10557
rect 21456 10591 21508 10600
rect 21456 10557 21465 10591
rect 21465 10557 21499 10591
rect 21499 10557 21508 10591
rect 21456 10548 21508 10557
rect 28172 10548 28224 10600
rect 29828 10548 29880 10600
rect 32128 10548 32180 10600
rect 33232 10659 33284 10668
rect 33232 10625 33241 10659
rect 33241 10625 33275 10659
rect 33275 10625 33284 10659
rect 33232 10616 33284 10625
rect 33324 10659 33376 10668
rect 33324 10625 33333 10659
rect 33333 10625 33367 10659
rect 33367 10625 33376 10659
rect 33324 10616 33376 10625
rect 36544 10616 36596 10668
rect 38568 10684 38620 10736
rect 38660 10684 38712 10736
rect 39028 10684 39080 10736
rect 41696 10727 41748 10736
rect 41696 10693 41705 10727
rect 41705 10693 41739 10727
rect 41739 10693 41748 10727
rect 41696 10684 41748 10693
rect 37280 10616 37332 10668
rect 37832 10659 37884 10668
rect 37832 10625 37841 10659
rect 37841 10625 37875 10659
rect 37875 10625 37884 10659
rect 37832 10616 37884 10625
rect 38752 10616 38804 10668
rect 41420 10659 41472 10668
rect 41420 10625 41429 10659
rect 41429 10625 41463 10659
rect 41463 10625 41472 10659
rect 41420 10616 41472 10625
rect 41788 10659 41840 10668
rect 41788 10625 41797 10659
rect 41797 10625 41831 10659
rect 41831 10625 41840 10659
rect 41788 10616 41840 10625
rect 42064 10616 42116 10668
rect 33600 10591 33652 10600
rect 33600 10557 33609 10591
rect 33609 10557 33643 10591
rect 33643 10557 33652 10591
rect 33600 10548 33652 10557
rect 33876 10591 33928 10600
rect 33876 10557 33885 10591
rect 33885 10557 33919 10591
rect 33919 10557 33928 10591
rect 33876 10548 33928 10557
rect 34888 10548 34940 10600
rect 37648 10548 37700 10600
rect 40224 10548 40276 10600
rect 41696 10548 41748 10600
rect 42248 10548 42300 10600
rect 44272 10727 44324 10736
rect 44272 10693 44281 10727
rect 44281 10693 44315 10727
rect 44315 10693 44324 10727
rect 44272 10684 44324 10693
rect 48872 10752 48924 10804
rect 49240 10752 49292 10804
rect 46296 10727 46348 10736
rect 46296 10693 46305 10727
rect 46305 10693 46339 10727
rect 46339 10693 46348 10727
rect 46296 10684 46348 10693
rect 46664 10684 46716 10736
rect 43352 10659 43404 10668
rect 43352 10625 43361 10659
rect 43361 10625 43395 10659
rect 43395 10625 43404 10659
rect 43352 10616 43404 10625
rect 43628 10659 43680 10668
rect 43628 10625 43637 10659
rect 43637 10625 43671 10659
rect 43671 10625 43680 10659
rect 43628 10616 43680 10625
rect 43720 10659 43772 10668
rect 43720 10625 43729 10659
rect 43729 10625 43763 10659
rect 43763 10625 43772 10659
rect 43720 10616 43772 10625
rect 46112 10659 46164 10668
rect 22008 10412 22060 10464
rect 26608 10412 26660 10464
rect 28448 10455 28500 10464
rect 28448 10421 28457 10455
rect 28457 10421 28491 10455
rect 28491 10421 28500 10455
rect 28448 10412 28500 10421
rect 32404 10455 32456 10464
rect 32404 10421 32413 10455
rect 32413 10421 32447 10455
rect 32447 10421 32456 10455
rect 32404 10412 32456 10421
rect 34612 10412 34664 10464
rect 43996 10591 44048 10600
rect 43996 10557 44005 10591
rect 44005 10557 44039 10591
rect 44039 10557 44048 10591
rect 43996 10548 44048 10557
rect 46112 10625 46116 10659
rect 46116 10625 46150 10659
rect 46150 10625 46164 10659
rect 46112 10616 46164 10625
rect 46572 10659 46624 10668
rect 46572 10625 46581 10659
rect 46581 10625 46615 10659
rect 46615 10625 46624 10659
rect 46572 10616 46624 10625
rect 47124 10616 47176 10668
rect 51356 10752 51408 10804
rect 51724 10752 51776 10804
rect 50804 10727 50856 10736
rect 50804 10693 50813 10727
rect 50813 10693 50847 10727
rect 50847 10693 50856 10727
rect 50804 10684 50856 10693
rect 51448 10684 51500 10736
rect 51816 10727 51868 10736
rect 51816 10693 51825 10727
rect 51825 10693 51859 10727
rect 51859 10693 51868 10727
rect 51816 10684 51868 10693
rect 45284 10480 45336 10532
rect 47032 10548 47084 10600
rect 47952 10548 48004 10600
rect 49424 10548 49476 10600
rect 44272 10412 44324 10464
rect 48228 10412 48280 10464
rect 49424 10455 49476 10464
rect 49424 10421 49433 10455
rect 49433 10421 49467 10455
rect 49467 10421 49476 10455
rect 49424 10412 49476 10421
rect 49608 10412 49660 10464
rect 50804 10412 50856 10464
rect 53104 10616 53156 10668
rect 53380 10616 53432 10668
rect 54760 10795 54812 10804
rect 54760 10761 54769 10795
rect 54769 10761 54803 10795
rect 54803 10761 54812 10795
rect 54760 10752 54812 10761
rect 54300 10684 54352 10736
rect 54208 10659 54260 10668
rect 54208 10625 54217 10659
rect 54217 10625 54251 10659
rect 54251 10625 54260 10659
rect 54208 10616 54260 10625
rect 52092 10548 52144 10600
rect 54576 10659 54628 10668
rect 54576 10625 54585 10659
rect 54585 10625 54619 10659
rect 54619 10625 54628 10659
rect 54576 10616 54628 10625
rect 56600 10548 56652 10600
rect 54852 10455 54904 10464
rect 54852 10421 54861 10455
rect 54861 10421 54895 10455
rect 54895 10421 54904 10455
rect 54852 10412 54904 10421
rect 55772 10412 55824 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 25412 10251 25464 10260
rect 25412 10217 25421 10251
rect 25421 10217 25455 10251
rect 25455 10217 25464 10251
rect 25412 10208 25464 10217
rect 30104 10208 30156 10260
rect 32680 10208 32732 10260
rect 32956 10251 33008 10260
rect 32956 10217 32965 10251
rect 32965 10217 32999 10251
rect 32999 10217 33008 10251
rect 32956 10208 33008 10217
rect 33876 10251 33928 10260
rect 33876 10217 33885 10251
rect 33885 10217 33919 10251
rect 33919 10217 33928 10251
rect 33876 10208 33928 10217
rect 39672 10251 39724 10260
rect 39672 10217 39681 10251
rect 39681 10217 39715 10251
rect 39715 10217 39724 10251
rect 39672 10208 39724 10217
rect 43352 10208 43404 10260
rect 43536 10251 43588 10260
rect 43536 10217 43545 10251
rect 43545 10217 43579 10251
rect 43579 10217 43588 10251
rect 43536 10208 43588 10217
rect 47952 10251 48004 10260
rect 47952 10217 47961 10251
rect 47961 10217 47995 10251
rect 47995 10217 48004 10251
rect 47952 10208 48004 10217
rect 48136 10208 48188 10260
rect 21456 10072 21508 10124
rect 26516 10072 26568 10124
rect 25412 10004 25464 10056
rect 26608 10047 26660 10056
rect 26608 10013 26617 10047
rect 26617 10013 26651 10047
rect 26651 10013 26660 10047
rect 26608 10004 26660 10013
rect 26792 10047 26844 10056
rect 26792 10013 26801 10047
rect 26801 10013 26835 10047
rect 26835 10013 26844 10047
rect 26792 10004 26844 10013
rect 26976 10047 27028 10056
rect 26976 10013 26985 10047
rect 26985 10013 27019 10047
rect 27019 10013 27028 10047
rect 26976 10004 27028 10013
rect 30932 10047 30984 10056
rect 30932 10013 30941 10047
rect 30941 10013 30975 10047
rect 30975 10013 30984 10047
rect 30932 10004 30984 10013
rect 32496 10004 32548 10056
rect 34612 10072 34664 10124
rect 39764 10140 39816 10192
rect 48688 10208 48740 10260
rect 49332 10208 49384 10260
rect 50068 10208 50120 10260
rect 51816 10208 51868 10260
rect 33048 10004 33100 10056
rect 34520 10047 34572 10056
rect 34520 10013 34529 10047
rect 34529 10013 34563 10047
rect 34563 10013 34572 10047
rect 34520 10004 34572 10013
rect 38844 10047 38896 10056
rect 38844 10013 38848 10047
rect 38848 10013 38882 10047
rect 38882 10013 38896 10047
rect 38844 10004 38896 10013
rect 39856 10072 39908 10124
rect 40224 10072 40276 10124
rect 43996 10072 44048 10124
rect 46940 10072 46992 10124
rect 47032 10115 47084 10124
rect 47032 10081 47041 10115
rect 47041 10081 47075 10115
rect 47075 10081 47084 10115
rect 47032 10072 47084 10081
rect 47216 10072 47268 10124
rect 47860 10072 47912 10124
rect 39212 10047 39264 10056
rect 39212 10013 39220 10047
rect 39220 10013 39254 10047
rect 39254 10013 39264 10047
rect 39212 10004 39264 10013
rect 39672 10004 39724 10056
rect 43352 10004 43404 10056
rect 43904 10004 43956 10056
rect 47676 10047 47728 10056
rect 47676 10013 47685 10047
rect 47685 10013 47719 10047
rect 47719 10013 47728 10047
rect 47676 10004 47728 10013
rect 48872 10140 48924 10192
rect 49424 10072 49476 10124
rect 48596 10004 48648 10056
rect 48872 10047 48924 10056
rect 48872 10013 48881 10047
rect 48881 10013 48915 10047
rect 48915 10013 48924 10047
rect 48872 10004 48924 10013
rect 26884 9979 26936 9988
rect 26884 9945 26893 9979
rect 26893 9945 26927 9979
rect 26927 9945 26936 9979
rect 26884 9936 26936 9945
rect 31208 9979 31260 9988
rect 31208 9945 31217 9979
rect 31217 9945 31251 9979
rect 31251 9945 31260 9979
rect 31208 9936 31260 9945
rect 32680 9936 32732 9988
rect 34796 9936 34848 9988
rect 40224 9979 40276 9988
rect 40224 9945 40233 9979
rect 40233 9945 40267 9979
rect 40267 9945 40276 9979
rect 40224 9936 40276 9945
rect 19708 9911 19760 9920
rect 19708 9877 19717 9911
rect 19717 9877 19751 9911
rect 19751 9877 19760 9911
rect 19708 9868 19760 9877
rect 27160 9911 27212 9920
rect 27160 9877 27169 9911
rect 27169 9877 27203 9911
rect 27203 9877 27212 9911
rect 27160 9868 27212 9877
rect 33876 9868 33928 9920
rect 34336 9868 34388 9920
rect 34704 9911 34756 9920
rect 34704 9877 34713 9911
rect 34713 9877 34747 9911
rect 34747 9877 34756 9911
rect 34704 9868 34756 9877
rect 37280 9868 37332 9920
rect 41236 9868 41288 9920
rect 41696 9911 41748 9920
rect 41696 9877 41705 9911
rect 41705 9877 41739 9911
rect 41739 9877 41748 9911
rect 41696 9868 41748 9877
rect 41972 9936 42024 9988
rect 44272 9936 44324 9988
rect 45192 9936 45244 9988
rect 45560 9979 45612 9988
rect 45560 9945 45569 9979
rect 45569 9945 45603 9979
rect 45603 9945 45612 9979
rect 45560 9936 45612 9945
rect 46572 9936 46624 9988
rect 47124 9911 47176 9920
rect 47124 9877 47133 9911
rect 47133 9877 47167 9911
rect 47167 9877 47176 9911
rect 47124 9868 47176 9877
rect 48320 9936 48372 9988
rect 49240 10047 49292 10056
rect 49240 10013 49249 10047
rect 49249 10013 49283 10047
rect 49283 10013 49292 10047
rect 49240 10004 49292 10013
rect 50160 10072 50212 10124
rect 51356 10140 51408 10192
rect 51632 10140 51684 10192
rect 49976 10004 50028 10056
rect 50344 10047 50396 10056
rect 50344 10013 50353 10047
rect 50353 10013 50387 10047
rect 50387 10013 50396 10047
rect 50344 10004 50396 10013
rect 50436 10047 50488 10056
rect 50436 10013 50446 10047
rect 50446 10013 50480 10047
rect 50480 10013 50488 10047
rect 50436 10004 50488 10013
rect 50712 10047 50764 10056
rect 50712 10013 50721 10047
rect 50721 10013 50755 10047
rect 50755 10013 50764 10047
rect 50712 10004 50764 10013
rect 50804 10047 50856 10056
rect 50804 10013 50818 10047
rect 50818 10013 50852 10047
rect 50852 10013 50856 10047
rect 50804 10004 50856 10013
rect 51264 10047 51316 10056
rect 51264 10013 51268 10047
rect 51268 10013 51302 10047
rect 51302 10013 51316 10047
rect 51264 10004 51316 10013
rect 51448 10047 51500 10056
rect 51448 10013 51457 10047
rect 51457 10013 51491 10047
rect 51491 10013 51500 10047
rect 51448 10004 51500 10013
rect 51540 10047 51592 10056
rect 51540 10013 51585 10047
rect 51585 10013 51592 10047
rect 51540 10004 51592 10013
rect 51724 10047 51776 10056
rect 51724 10013 51733 10047
rect 51733 10013 51767 10047
rect 51767 10013 51776 10047
rect 51724 10004 51776 10013
rect 52000 10140 52052 10192
rect 52184 10140 52236 10192
rect 56600 10072 56652 10124
rect 49332 9936 49384 9988
rect 52092 10004 52144 10056
rect 52368 10047 52420 10056
rect 52368 10013 52382 10047
rect 52382 10013 52416 10047
rect 52416 10013 52420 10047
rect 52368 10004 52420 10013
rect 54852 10004 54904 10056
rect 52184 9979 52236 9988
rect 52184 9945 52193 9979
rect 52193 9945 52227 9979
rect 52227 9945 52236 9979
rect 52184 9936 52236 9945
rect 49700 9868 49752 9920
rect 49792 9911 49844 9920
rect 49792 9877 49801 9911
rect 49801 9877 49835 9911
rect 49835 9877 49844 9911
rect 49792 9868 49844 9877
rect 50988 9911 51040 9920
rect 50988 9877 50997 9911
rect 50997 9877 51031 9911
rect 51031 9877 51040 9911
rect 50988 9868 51040 9877
rect 51264 9868 51316 9920
rect 51448 9868 51500 9920
rect 52920 9979 52972 9988
rect 52920 9945 52929 9979
rect 52929 9945 52963 9979
rect 52963 9945 52972 9979
rect 52920 9936 52972 9945
rect 54208 9936 54260 9988
rect 53012 9868 53064 9920
rect 54392 9911 54444 9920
rect 54392 9877 54401 9911
rect 54401 9877 54435 9911
rect 54435 9877 54444 9911
rect 55588 9979 55640 9988
rect 55588 9945 55597 9979
rect 55597 9945 55631 9979
rect 55631 9945 55640 9979
rect 55588 9936 55640 9945
rect 54392 9868 54444 9877
rect 55772 9868 55824 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 66314 9766 66366 9818
rect 66378 9766 66430 9818
rect 66442 9766 66494 9818
rect 66506 9766 66558 9818
rect 66570 9766 66622 9818
rect 26884 9664 26936 9716
rect 31208 9664 31260 9716
rect 28448 9596 28500 9648
rect 28816 9596 28868 9648
rect 26516 9528 26568 9580
rect 27988 9503 28040 9512
rect 27988 9469 27997 9503
rect 27997 9469 28031 9503
rect 28031 9469 28040 9503
rect 27988 9460 28040 9469
rect 31024 9528 31076 9580
rect 32404 9596 32456 9648
rect 31852 9528 31904 9580
rect 34704 9596 34756 9648
rect 35716 9639 35768 9648
rect 35716 9605 35725 9639
rect 35725 9605 35759 9639
rect 35759 9605 35768 9639
rect 35716 9596 35768 9605
rect 40224 9664 40276 9716
rect 38200 9596 38252 9648
rect 38936 9596 38988 9648
rect 40040 9596 40092 9648
rect 34336 9571 34388 9580
rect 34336 9537 34345 9571
rect 34345 9537 34379 9571
rect 34379 9537 34388 9571
rect 34336 9528 34388 9537
rect 34796 9528 34848 9580
rect 28816 9460 28868 9512
rect 33048 9460 33100 9512
rect 33416 9460 33468 9512
rect 34244 9460 34296 9512
rect 34612 9460 34664 9512
rect 35256 9571 35308 9580
rect 35256 9537 35265 9571
rect 35265 9537 35299 9571
rect 35299 9537 35308 9571
rect 35256 9528 35308 9537
rect 37648 9571 37700 9580
rect 37648 9537 37657 9571
rect 37657 9537 37691 9571
rect 37691 9537 37700 9571
rect 37648 9528 37700 9537
rect 40684 9528 40736 9580
rect 35900 9460 35952 9512
rect 36636 9460 36688 9512
rect 37280 9460 37332 9512
rect 37924 9503 37976 9512
rect 37924 9469 37933 9503
rect 37933 9469 37967 9503
rect 37967 9469 37976 9503
rect 37924 9460 37976 9469
rect 30932 9392 30984 9444
rect 31760 9392 31812 9444
rect 32680 9392 32732 9444
rect 33784 9435 33836 9444
rect 33784 9401 33793 9435
rect 33793 9401 33827 9435
rect 33827 9401 33836 9435
rect 33784 9392 33836 9401
rect 29828 9367 29880 9376
rect 29828 9333 29837 9367
rect 29837 9333 29871 9367
rect 29871 9333 29880 9367
rect 29828 9324 29880 9333
rect 33232 9324 33284 9376
rect 36176 9392 36228 9444
rect 37464 9392 37516 9444
rect 35440 9324 35492 9376
rect 35900 9367 35952 9376
rect 35900 9333 35909 9367
rect 35909 9333 35943 9367
rect 35943 9333 35952 9367
rect 35900 9324 35952 9333
rect 36268 9324 36320 9376
rect 38384 9324 38436 9376
rect 39304 9324 39356 9376
rect 42340 9528 42392 9580
rect 42800 9571 42852 9580
rect 42800 9537 42809 9571
rect 42809 9537 42843 9571
rect 42843 9537 42852 9571
rect 42800 9528 42852 9537
rect 43260 9571 43312 9580
rect 43260 9537 43264 9571
rect 43264 9537 43298 9571
rect 43298 9537 43312 9571
rect 41696 9460 41748 9512
rect 42708 9460 42760 9512
rect 43260 9528 43312 9537
rect 43536 9571 43588 9580
rect 43536 9537 43581 9571
rect 43581 9537 43588 9571
rect 43536 9528 43588 9537
rect 45284 9664 45336 9716
rect 45560 9664 45612 9716
rect 46112 9664 46164 9716
rect 49976 9664 50028 9716
rect 50344 9664 50396 9716
rect 48688 9596 48740 9648
rect 49148 9596 49200 9648
rect 45928 9571 45980 9580
rect 45928 9537 45937 9571
rect 45937 9537 45971 9571
rect 45971 9537 45980 9571
rect 45928 9528 45980 9537
rect 47124 9528 47176 9580
rect 39488 9367 39540 9376
rect 39488 9333 39497 9367
rect 39497 9333 39531 9367
rect 39531 9333 39540 9367
rect 39488 9324 39540 9333
rect 40316 9367 40368 9376
rect 40316 9333 40325 9367
rect 40325 9333 40359 9367
rect 40359 9333 40368 9367
rect 40316 9324 40368 9333
rect 41972 9324 42024 9376
rect 47216 9460 47268 9512
rect 49516 9528 49568 9580
rect 49700 9596 49752 9648
rect 50252 9596 50304 9648
rect 50712 9664 50764 9716
rect 51172 9664 51224 9716
rect 51724 9664 51776 9716
rect 52000 9664 52052 9716
rect 52920 9664 52972 9716
rect 54944 9664 54996 9716
rect 50068 9460 50120 9512
rect 50344 9571 50396 9580
rect 50344 9537 50353 9571
rect 50353 9537 50387 9571
rect 50387 9537 50396 9571
rect 50344 9528 50396 9537
rect 50436 9460 50488 9512
rect 49976 9392 50028 9444
rect 43720 9324 43772 9376
rect 46848 9324 46900 9376
rect 48872 9324 48924 9376
rect 50160 9324 50212 9376
rect 50344 9392 50396 9444
rect 51632 9639 51684 9648
rect 50896 9528 50948 9580
rect 51632 9605 51641 9639
rect 51641 9605 51675 9639
rect 51675 9605 51684 9639
rect 51632 9596 51684 9605
rect 55496 9634 55548 9686
rect 55588 9664 55640 9716
rect 51356 9528 51408 9580
rect 53012 9571 53064 9580
rect 53012 9537 53021 9571
rect 53021 9537 53055 9571
rect 53055 9537 53064 9571
rect 53012 9528 53064 9537
rect 54208 9528 54260 9580
rect 54484 9571 54536 9580
rect 54484 9537 54493 9571
rect 54493 9537 54527 9571
rect 54527 9537 54536 9571
rect 54484 9528 54536 9537
rect 54668 9571 54720 9580
rect 54668 9537 54677 9571
rect 54677 9537 54711 9571
rect 54711 9537 54720 9571
rect 54668 9528 54720 9537
rect 54392 9460 54444 9512
rect 54944 9528 54996 9580
rect 55312 9528 55364 9580
rect 55496 9571 55548 9580
rect 55496 9537 55505 9571
rect 55505 9537 55539 9571
rect 55539 9537 55548 9571
rect 55496 9528 55548 9537
rect 56600 9571 56652 9580
rect 56600 9537 56609 9571
rect 56609 9537 56643 9571
rect 56643 9537 56652 9571
rect 56600 9528 56652 9537
rect 50804 9392 50856 9444
rect 51172 9392 51224 9444
rect 51448 9392 51500 9444
rect 52368 9392 52420 9444
rect 51908 9324 51960 9376
rect 53196 9367 53248 9376
rect 53196 9333 53205 9367
rect 53205 9333 53239 9367
rect 53239 9333 53248 9367
rect 53196 9324 53248 9333
rect 55036 9367 55088 9376
rect 55036 9333 55045 9367
rect 55045 9333 55079 9367
rect 55079 9333 55088 9367
rect 55036 9324 55088 9333
rect 55496 9324 55548 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 28264 9163 28316 9172
rect 28264 9129 28273 9163
rect 28273 9129 28307 9163
rect 28307 9129 28316 9163
rect 28264 9120 28316 9129
rect 31300 9120 31352 9172
rect 31484 9120 31536 9172
rect 31852 9163 31904 9172
rect 31852 9129 31861 9163
rect 31861 9129 31895 9163
rect 31895 9129 31904 9163
rect 31852 9120 31904 9129
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 27160 8984 27212 9036
rect 31208 8916 31260 8968
rect 33600 8984 33652 9036
rect 37924 9120 37976 9172
rect 38384 9120 38436 9172
rect 42616 9120 42668 9172
rect 42892 9163 42944 9172
rect 42892 9129 42901 9163
rect 42901 9129 42935 9163
rect 42935 9129 42944 9163
rect 42892 9120 42944 9129
rect 43260 9120 43312 9172
rect 49516 9120 49568 9172
rect 49700 9163 49752 9172
rect 49700 9129 49709 9163
rect 49709 9129 49743 9163
rect 49743 9129 49752 9163
rect 49700 9120 49752 9129
rect 49884 9120 49936 9172
rect 50896 9120 50948 9172
rect 55036 9120 55088 9172
rect 55312 9120 55364 9172
rect 35992 9052 36044 9104
rect 35164 8984 35216 9036
rect 31484 8959 31536 8968
rect 31484 8925 31493 8959
rect 31493 8925 31527 8959
rect 31527 8925 31536 8959
rect 31484 8916 31536 8925
rect 31668 8959 31720 8968
rect 31668 8925 31677 8959
rect 31677 8925 31711 8959
rect 31711 8925 31720 8959
rect 31668 8916 31720 8925
rect 32220 8959 32272 8968
rect 32220 8925 32227 8959
rect 32227 8925 32272 8959
rect 22008 8780 22060 8832
rect 31392 8848 31444 8900
rect 31576 8891 31628 8900
rect 31576 8857 31585 8891
rect 31585 8857 31619 8891
rect 31619 8857 31628 8891
rect 31576 8848 31628 8857
rect 28816 8780 28868 8832
rect 31484 8780 31536 8832
rect 32220 8916 32272 8925
rect 32404 8959 32456 8968
rect 32404 8925 32410 8959
rect 32410 8925 32444 8959
rect 32444 8925 32456 8959
rect 32404 8916 32456 8925
rect 35900 8959 35952 8968
rect 35900 8925 35909 8959
rect 35909 8925 35943 8959
rect 35943 8925 35952 8959
rect 35900 8916 35952 8925
rect 37004 9052 37056 9104
rect 37280 9095 37332 9104
rect 37280 9061 37289 9095
rect 37289 9061 37323 9095
rect 37323 9061 37332 9095
rect 37280 9052 37332 9061
rect 38568 9052 38620 9104
rect 40316 9052 40368 9104
rect 36820 8984 36872 9036
rect 36360 8959 36412 8968
rect 36360 8925 36374 8959
rect 36374 8925 36408 8959
rect 36408 8925 36412 8959
rect 36360 8916 36412 8925
rect 36636 8959 36688 8968
rect 36636 8925 36645 8959
rect 36645 8925 36679 8959
rect 36679 8925 36688 8959
rect 36636 8916 36688 8925
rect 37464 8984 37516 9036
rect 38016 8984 38068 9036
rect 42616 8984 42668 9036
rect 32220 8780 32272 8832
rect 32772 8848 32824 8900
rect 33048 8891 33100 8900
rect 33048 8857 33057 8891
rect 33057 8857 33091 8891
rect 33091 8857 33100 8891
rect 33048 8848 33100 8857
rect 32588 8780 32640 8832
rect 32680 8823 32732 8832
rect 32680 8789 32689 8823
rect 32689 8789 32723 8823
rect 32723 8789 32732 8823
rect 32680 8780 32732 8789
rect 33968 8780 34020 8832
rect 34428 8848 34480 8900
rect 36176 8891 36228 8900
rect 36176 8857 36185 8891
rect 36185 8857 36219 8891
rect 36219 8857 36228 8891
rect 36176 8848 36228 8857
rect 34704 8823 34756 8832
rect 34704 8789 34713 8823
rect 34713 8789 34747 8823
rect 34747 8789 34756 8823
rect 34704 8780 34756 8789
rect 36544 8823 36596 8832
rect 36544 8789 36553 8823
rect 36553 8789 36587 8823
rect 36587 8789 36596 8823
rect 36544 8780 36596 8789
rect 36636 8780 36688 8832
rect 37648 8848 37700 8900
rect 38292 8916 38344 8968
rect 38384 8959 38436 8968
rect 38384 8925 38393 8959
rect 38393 8925 38427 8959
rect 38427 8925 38436 8959
rect 38384 8916 38436 8925
rect 38476 8959 38528 8968
rect 38476 8925 38485 8959
rect 38485 8925 38519 8959
rect 38519 8925 38528 8959
rect 38476 8916 38528 8925
rect 39488 8916 39540 8968
rect 41972 8959 42024 8968
rect 41972 8925 41981 8959
rect 41981 8925 42015 8959
rect 42015 8925 42024 8959
rect 41972 8916 42024 8925
rect 42064 8959 42116 8968
rect 42064 8925 42073 8959
rect 42073 8925 42107 8959
rect 42107 8925 42116 8959
rect 42064 8916 42116 8925
rect 41696 8848 41748 8900
rect 46296 9052 46348 9104
rect 50344 9052 50396 9104
rect 50712 9052 50764 9104
rect 51080 9052 51132 9104
rect 44180 8984 44232 9036
rect 49608 8984 49660 9036
rect 49700 8984 49752 9036
rect 50988 8984 51040 9036
rect 44088 8959 44140 8968
rect 44088 8925 44097 8959
rect 44097 8925 44131 8959
rect 44131 8925 44140 8959
rect 44088 8916 44140 8925
rect 44364 8959 44416 8968
rect 44364 8925 44372 8959
rect 44372 8925 44406 8959
rect 44406 8925 44416 8959
rect 44364 8916 44416 8925
rect 44456 8959 44508 8968
rect 44456 8925 44465 8959
rect 44465 8925 44499 8959
rect 44499 8925 44508 8959
rect 44456 8916 44508 8925
rect 45468 8916 45520 8968
rect 49056 8916 49108 8968
rect 51080 8916 51132 8968
rect 44916 8848 44968 8900
rect 49700 8848 49752 8900
rect 50344 8848 50396 8900
rect 50988 8891 51040 8900
rect 50988 8857 50997 8891
rect 50997 8857 51031 8891
rect 51031 8857 51040 8891
rect 50988 8848 51040 8857
rect 51264 8959 51316 8968
rect 51264 8925 51273 8959
rect 51273 8925 51307 8959
rect 51307 8925 51316 8959
rect 51264 8916 51316 8925
rect 51632 8848 51684 8900
rect 38384 8780 38436 8832
rect 38844 8780 38896 8832
rect 40684 8780 40736 8832
rect 40868 8780 40920 8832
rect 41788 8780 41840 8832
rect 42340 8780 42392 8832
rect 43812 8823 43864 8832
rect 43812 8789 43821 8823
rect 43821 8789 43855 8823
rect 43855 8789 43864 8823
rect 43812 8780 43864 8789
rect 46848 8780 46900 8832
rect 48964 8780 49016 8832
rect 50160 8823 50212 8832
rect 50160 8789 50169 8823
rect 50169 8789 50203 8823
rect 50203 8789 50212 8823
rect 50160 8780 50212 8789
rect 51356 8780 51408 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 66314 8678 66366 8730
rect 66378 8678 66430 8730
rect 66442 8678 66494 8730
rect 66506 8678 66558 8730
rect 66570 8678 66622 8730
rect 29460 8508 29512 8560
rect 31760 8576 31812 8628
rect 33048 8576 33100 8628
rect 35348 8576 35400 8628
rect 35440 8576 35492 8628
rect 35532 8576 35584 8628
rect 31300 8508 31352 8560
rect 32128 8508 32180 8560
rect 32588 8508 32640 8560
rect 32772 8508 32824 8560
rect 31024 8483 31076 8492
rect 31024 8449 31028 8483
rect 31028 8449 31062 8483
rect 31062 8449 31076 8483
rect 31024 8440 31076 8449
rect 31116 8483 31168 8492
rect 31116 8449 31125 8483
rect 31125 8449 31159 8483
rect 31159 8449 31168 8483
rect 31116 8440 31168 8449
rect 31392 8483 31444 8492
rect 31392 8449 31400 8483
rect 31400 8449 31434 8483
rect 31434 8449 31444 8483
rect 31392 8440 31444 8449
rect 31484 8483 31536 8492
rect 31484 8449 31493 8483
rect 31493 8449 31527 8483
rect 31527 8449 31536 8483
rect 31484 8440 31536 8449
rect 32680 8440 32732 8492
rect 34704 8440 34756 8492
rect 29184 8415 29236 8424
rect 29184 8381 29193 8415
rect 29193 8381 29227 8415
rect 29227 8381 29236 8415
rect 29184 8372 29236 8381
rect 32220 8372 32272 8424
rect 32956 8372 33008 8424
rect 33232 8415 33284 8424
rect 33232 8381 33241 8415
rect 33241 8381 33275 8415
rect 33275 8381 33284 8415
rect 33232 8372 33284 8381
rect 33692 8372 33744 8424
rect 33876 8372 33928 8424
rect 31116 8304 31168 8356
rect 31392 8304 31444 8356
rect 32772 8304 32824 8356
rect 35164 8483 35216 8492
rect 35164 8449 35174 8483
rect 35174 8449 35208 8483
rect 35208 8449 35216 8483
rect 35164 8440 35216 8449
rect 35440 8483 35492 8492
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 35716 8440 35768 8492
rect 36176 8483 36228 8492
rect 36176 8449 36185 8483
rect 36185 8449 36219 8483
rect 36219 8449 36228 8483
rect 36176 8440 36228 8449
rect 36268 8483 36320 8492
rect 36268 8449 36282 8483
rect 36282 8449 36316 8483
rect 36316 8449 36320 8483
rect 36544 8576 36596 8628
rect 37556 8576 37608 8628
rect 38476 8576 38528 8628
rect 36728 8551 36780 8560
rect 36728 8517 36737 8551
rect 36737 8517 36771 8551
rect 36771 8517 36780 8551
rect 36728 8508 36780 8517
rect 37188 8508 37240 8560
rect 37280 8551 37332 8560
rect 37280 8517 37289 8551
rect 37289 8517 37323 8551
rect 37323 8517 37332 8551
rect 37280 8508 37332 8517
rect 38108 8508 38160 8560
rect 42800 8576 42852 8628
rect 43168 8576 43220 8628
rect 43536 8576 43588 8628
rect 45468 8619 45520 8628
rect 36268 8440 36320 8449
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 37648 8440 37700 8492
rect 35440 8304 35492 8356
rect 30380 8236 30432 8288
rect 37188 8372 37240 8424
rect 37280 8372 37332 8424
rect 36084 8236 36136 8288
rect 37464 8304 37516 8356
rect 38016 8304 38068 8356
rect 40316 8372 40368 8424
rect 40868 8415 40920 8424
rect 40868 8381 40877 8415
rect 40877 8381 40911 8415
rect 40911 8381 40920 8415
rect 40868 8372 40920 8381
rect 37372 8236 37424 8288
rect 38292 8236 38344 8288
rect 39212 8304 39264 8356
rect 41420 8508 41472 8560
rect 41512 8483 41564 8492
rect 40132 8236 40184 8288
rect 41512 8449 41520 8483
rect 41520 8449 41554 8483
rect 41554 8449 41564 8483
rect 41512 8440 41564 8449
rect 41696 8508 41748 8560
rect 42340 8440 42392 8492
rect 42616 8483 42668 8492
rect 42616 8449 42625 8483
rect 42625 8449 42659 8483
rect 42659 8449 42668 8483
rect 42616 8440 42668 8449
rect 42708 8483 42760 8492
rect 42708 8449 42718 8483
rect 42718 8449 42752 8483
rect 42752 8449 42760 8483
rect 42708 8440 42760 8449
rect 42892 8483 42944 8492
rect 42892 8449 42901 8483
rect 42901 8449 42935 8483
rect 42935 8449 42944 8483
rect 42892 8440 42944 8449
rect 42984 8483 43036 8492
rect 42984 8449 42993 8483
rect 42993 8449 43027 8483
rect 43027 8449 43036 8483
rect 42984 8440 43036 8449
rect 43720 8508 43772 8560
rect 43352 8440 43404 8492
rect 43812 8440 43864 8492
rect 43720 8415 43772 8424
rect 43720 8381 43729 8415
rect 43729 8381 43763 8415
rect 43763 8381 43772 8415
rect 43720 8372 43772 8381
rect 44180 8483 44232 8492
rect 44180 8449 44189 8483
rect 44189 8449 44223 8483
rect 44223 8449 44232 8483
rect 44180 8440 44232 8449
rect 45468 8585 45477 8619
rect 45477 8585 45511 8619
rect 45511 8585 45520 8619
rect 45468 8576 45520 8585
rect 42064 8236 42116 8288
rect 42708 8236 42760 8288
rect 44732 8483 44784 8492
rect 44732 8449 44742 8483
rect 44742 8449 44776 8483
rect 44776 8449 44784 8483
rect 44732 8440 44784 8449
rect 45376 8508 45428 8560
rect 44916 8483 44968 8492
rect 44916 8449 44925 8483
rect 44925 8449 44959 8483
rect 44959 8449 44968 8483
rect 44916 8440 44968 8449
rect 45100 8483 45152 8492
rect 45100 8449 45114 8483
rect 45114 8449 45148 8483
rect 45148 8449 45152 8483
rect 48780 8576 48832 8628
rect 50528 8576 50580 8628
rect 50804 8576 50856 8628
rect 50896 8576 50948 8628
rect 51172 8619 51224 8628
rect 51172 8585 51181 8619
rect 51181 8585 51215 8619
rect 51215 8585 51224 8619
rect 51172 8576 51224 8585
rect 46572 8508 46624 8560
rect 47216 8508 47268 8560
rect 50712 8551 50764 8560
rect 50712 8517 50721 8551
rect 50721 8517 50755 8551
rect 50755 8517 50764 8551
rect 50712 8508 50764 8517
rect 45100 8440 45152 8449
rect 48872 8483 48924 8492
rect 48872 8449 48881 8483
rect 48881 8449 48915 8483
rect 48915 8449 48924 8483
rect 48872 8440 48924 8449
rect 49792 8440 49844 8492
rect 50528 8483 50580 8492
rect 50528 8449 50535 8483
rect 50535 8449 50580 8483
rect 50528 8440 50580 8449
rect 51080 8508 51132 8560
rect 52184 8508 52236 8560
rect 45652 8372 45704 8424
rect 47124 8415 47176 8424
rect 47124 8381 47133 8415
rect 47133 8381 47167 8415
rect 47167 8381 47176 8415
rect 47124 8372 47176 8381
rect 45284 8279 45336 8288
rect 45284 8245 45293 8279
rect 45293 8245 45327 8279
rect 45327 8245 45336 8279
rect 45284 8236 45336 8245
rect 46940 8236 46992 8288
rect 48044 8372 48096 8424
rect 48964 8372 49016 8424
rect 50252 8415 50304 8424
rect 50252 8381 50261 8415
rect 50261 8381 50295 8415
rect 50295 8381 50304 8415
rect 50252 8372 50304 8381
rect 50620 8372 50672 8424
rect 51264 8483 51316 8492
rect 51264 8449 51273 8483
rect 51273 8449 51307 8483
rect 51307 8449 51316 8483
rect 51264 8440 51316 8449
rect 51632 8483 51684 8492
rect 51632 8449 51641 8483
rect 51641 8449 51675 8483
rect 51675 8449 51684 8483
rect 51632 8440 51684 8449
rect 51724 8483 51776 8492
rect 51724 8449 51738 8483
rect 51738 8449 51772 8483
rect 51772 8449 51776 8483
rect 51724 8440 51776 8449
rect 53472 8483 53524 8492
rect 53472 8449 53481 8483
rect 53481 8449 53515 8483
rect 53515 8449 53524 8483
rect 53472 8440 53524 8449
rect 54852 8440 54904 8492
rect 78036 8483 78088 8492
rect 78036 8449 78045 8483
rect 78045 8449 78079 8483
rect 78079 8449 78088 8483
rect 78036 8440 78088 8449
rect 51264 8304 51316 8356
rect 52000 8347 52052 8356
rect 52000 8313 52009 8347
rect 52009 8313 52043 8347
rect 52043 8313 52052 8347
rect 52000 8304 52052 8313
rect 52920 8304 52972 8356
rect 53564 8304 53616 8356
rect 78220 8347 78272 8356
rect 78220 8313 78229 8347
rect 78229 8313 78263 8347
rect 78263 8313 78272 8347
rect 78220 8304 78272 8313
rect 48504 8236 48556 8288
rect 50068 8236 50120 8288
rect 50896 8236 50948 8288
rect 51724 8236 51776 8288
rect 53288 8279 53340 8288
rect 53288 8245 53297 8279
rect 53297 8245 53331 8279
rect 53331 8245 53340 8279
rect 53288 8236 53340 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 29184 8032 29236 8084
rect 35440 8075 35492 8084
rect 35440 8041 35449 8075
rect 35449 8041 35483 8075
rect 35483 8041 35492 8075
rect 35440 8032 35492 8041
rect 31116 7896 31168 7948
rect 30380 7871 30432 7880
rect 30380 7837 30389 7871
rect 30389 7837 30423 7871
rect 30423 7837 30432 7871
rect 30380 7828 30432 7837
rect 30564 7871 30616 7880
rect 30564 7837 30573 7871
rect 30573 7837 30607 7871
rect 30607 7837 30616 7871
rect 30564 7828 30616 7837
rect 31024 7828 31076 7880
rect 31484 7828 31536 7880
rect 31668 7871 31720 7880
rect 31668 7837 31677 7871
rect 31677 7837 31711 7871
rect 31711 7837 31720 7871
rect 31668 7828 31720 7837
rect 32312 7896 32364 7948
rect 32036 7871 32088 7880
rect 32036 7837 32045 7871
rect 32045 7837 32079 7871
rect 32079 7837 32088 7871
rect 32036 7828 32088 7837
rect 34428 7828 34480 7880
rect 31024 7692 31076 7744
rect 31760 7692 31812 7744
rect 32588 7760 32640 7812
rect 34704 7760 34756 7812
rect 36084 8007 36136 8016
rect 36084 7973 36093 8007
rect 36093 7973 36127 8007
rect 36127 7973 36136 8007
rect 36084 7964 36136 7973
rect 36268 7964 36320 8016
rect 41972 8032 42024 8084
rect 42616 8075 42668 8084
rect 42616 8041 42625 8075
rect 42625 8041 42659 8075
rect 42659 8041 42668 8075
rect 42616 8032 42668 8041
rect 35900 7939 35952 7948
rect 35900 7905 35909 7939
rect 35909 7905 35943 7939
rect 35943 7905 35952 7939
rect 35900 7896 35952 7905
rect 37280 7896 37332 7948
rect 37648 7939 37700 7948
rect 37648 7905 37657 7939
rect 37657 7905 37691 7939
rect 37691 7905 37700 7939
rect 37648 7896 37700 7905
rect 38476 7939 38528 7948
rect 38476 7905 38485 7939
rect 38485 7905 38519 7939
rect 38519 7905 38528 7939
rect 38476 7896 38528 7905
rect 38844 7828 38896 7880
rect 38660 7692 38712 7744
rect 38752 7692 38804 7744
rect 41880 7964 41932 8016
rect 39856 7939 39908 7948
rect 39856 7905 39865 7939
rect 39865 7905 39899 7939
rect 39899 7905 39908 7939
rect 39856 7896 39908 7905
rect 40132 7939 40184 7948
rect 40132 7905 40141 7939
rect 40141 7905 40175 7939
rect 40175 7905 40184 7939
rect 40132 7896 40184 7905
rect 39212 7871 39264 7880
rect 39212 7837 39221 7871
rect 39221 7837 39255 7871
rect 39255 7837 39264 7871
rect 39212 7828 39264 7837
rect 39304 7871 39356 7880
rect 39304 7837 39313 7871
rect 39313 7837 39347 7871
rect 39347 7837 39356 7871
rect 39304 7828 39356 7837
rect 41236 7828 41288 7880
rect 41880 7828 41932 7880
rect 43076 8032 43128 8084
rect 43352 8075 43404 8084
rect 43352 8041 43361 8075
rect 43361 8041 43395 8075
rect 43395 8041 43404 8075
rect 43352 8032 43404 8041
rect 45100 8032 45152 8084
rect 45928 8075 45980 8084
rect 45928 8041 45937 8075
rect 45937 8041 45971 8075
rect 45971 8041 45980 8075
rect 45928 8032 45980 8041
rect 47124 8032 47176 8084
rect 49976 8075 50028 8084
rect 49976 8041 49985 8075
rect 49985 8041 50019 8075
rect 50019 8041 50028 8075
rect 49976 8032 50028 8041
rect 50252 8032 50304 8084
rect 50804 8032 50856 8084
rect 51264 8032 51316 8084
rect 51448 8032 51500 8084
rect 52184 8032 52236 8084
rect 54852 8075 54904 8084
rect 54852 8041 54861 8075
rect 54861 8041 54895 8075
rect 54895 8041 54904 8075
rect 54852 8032 54904 8041
rect 44180 7964 44232 8016
rect 55772 7964 55824 8016
rect 46848 7939 46900 7948
rect 46848 7905 46857 7939
rect 46857 7905 46891 7939
rect 46891 7905 46900 7939
rect 46848 7896 46900 7905
rect 48044 7896 48096 7948
rect 48504 7939 48556 7948
rect 48504 7905 48513 7939
rect 48513 7905 48547 7939
rect 48547 7905 48556 7939
rect 48504 7896 48556 7905
rect 50620 7896 50672 7948
rect 51816 7896 51868 7948
rect 53380 7896 53432 7948
rect 54024 7896 54076 7948
rect 54668 7896 54720 7948
rect 42340 7803 42392 7812
rect 42340 7769 42349 7803
rect 42349 7769 42383 7803
rect 42383 7769 42392 7803
rect 42340 7760 42392 7769
rect 45376 7871 45428 7880
rect 45376 7837 45385 7871
rect 45385 7837 45419 7871
rect 45419 7837 45428 7871
rect 45376 7828 45428 7837
rect 45652 7871 45704 7880
rect 45652 7837 45661 7871
rect 45661 7837 45695 7871
rect 45695 7837 45704 7871
rect 45652 7828 45704 7837
rect 45744 7871 45796 7880
rect 45744 7837 45753 7871
rect 45753 7837 45787 7871
rect 45787 7837 45796 7871
rect 45744 7828 45796 7837
rect 42616 7760 42668 7812
rect 45836 7760 45888 7812
rect 47124 7871 47176 7880
rect 47124 7837 47133 7871
rect 47133 7837 47167 7871
rect 47167 7837 47176 7871
rect 47124 7828 47176 7837
rect 42708 7692 42760 7744
rect 47676 7871 47728 7880
rect 47676 7837 47685 7871
rect 47685 7837 47719 7871
rect 47719 7837 47728 7871
rect 47676 7828 47728 7837
rect 48228 7760 48280 7812
rect 51540 7760 51592 7812
rect 53288 7760 53340 7812
rect 52920 7692 52972 7744
rect 53656 7692 53708 7744
rect 54944 7828 54996 7880
rect 78036 8075 78088 8084
rect 78036 8041 78045 8075
rect 78045 8041 78079 8075
rect 78079 8041 78088 8075
rect 78036 8032 78088 8041
rect 55588 7803 55640 7812
rect 55588 7769 55597 7803
rect 55597 7769 55631 7803
rect 55631 7769 55640 7803
rect 55588 7760 55640 7769
rect 55036 7692 55088 7744
rect 77668 7692 77720 7744
rect 78404 7735 78456 7744
rect 78404 7701 78413 7735
rect 78413 7701 78447 7735
rect 78447 7701 78456 7735
rect 78404 7692 78456 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 66314 7590 66366 7642
rect 66378 7590 66430 7642
rect 66442 7590 66494 7642
rect 66506 7590 66558 7642
rect 66570 7590 66622 7642
rect 31852 7488 31904 7540
rect 37280 7531 37332 7540
rect 37280 7497 37289 7531
rect 37289 7497 37323 7531
rect 37323 7497 37332 7531
rect 37280 7488 37332 7497
rect 38660 7488 38712 7540
rect 40776 7488 40828 7540
rect 42524 7488 42576 7540
rect 37372 7420 37424 7472
rect 41972 7420 42024 7472
rect 30932 7395 30984 7404
rect 30932 7361 30941 7395
rect 30941 7361 30975 7395
rect 30975 7361 30984 7395
rect 30932 7352 30984 7361
rect 31024 7395 31076 7404
rect 31024 7361 31033 7395
rect 31033 7361 31067 7395
rect 31067 7361 31076 7395
rect 31024 7352 31076 7361
rect 32772 7395 32824 7404
rect 32772 7361 32781 7395
rect 32781 7361 32815 7395
rect 32815 7361 32824 7395
rect 32772 7352 32824 7361
rect 33692 7395 33744 7404
rect 30564 7284 30616 7336
rect 33692 7361 33701 7395
rect 33701 7361 33735 7395
rect 33735 7361 33744 7395
rect 33692 7352 33744 7361
rect 33876 7395 33928 7404
rect 33876 7361 33885 7395
rect 33885 7361 33919 7395
rect 33919 7361 33928 7395
rect 33876 7352 33928 7361
rect 39856 7352 39908 7404
rect 40776 7352 40828 7404
rect 41512 7352 41564 7404
rect 41696 7352 41748 7404
rect 42340 7352 42392 7404
rect 42616 7395 42668 7404
rect 42616 7361 42625 7395
rect 42625 7361 42659 7395
rect 42659 7361 42668 7395
rect 42616 7352 42668 7361
rect 33048 7284 33100 7336
rect 38752 7327 38804 7336
rect 38752 7293 38761 7327
rect 38761 7293 38795 7327
rect 38795 7293 38804 7327
rect 38752 7284 38804 7293
rect 41788 7284 41840 7336
rect 43352 7216 43404 7268
rect 30748 7191 30800 7200
rect 30748 7157 30757 7191
rect 30757 7157 30791 7191
rect 30791 7157 30800 7191
rect 30748 7148 30800 7157
rect 34060 7191 34112 7200
rect 34060 7157 34069 7191
rect 34069 7157 34103 7191
rect 34103 7157 34112 7191
rect 34060 7148 34112 7157
rect 38752 7148 38804 7200
rect 41420 7148 41472 7200
rect 43076 7148 43128 7200
rect 43720 7395 43772 7404
rect 43720 7361 43729 7395
rect 43729 7361 43763 7395
rect 43763 7361 43772 7395
rect 43720 7352 43772 7361
rect 44456 7488 44508 7540
rect 46480 7488 46532 7540
rect 47676 7488 47728 7540
rect 51540 7531 51592 7540
rect 51540 7497 51549 7531
rect 51549 7497 51583 7531
rect 51583 7497 51592 7531
rect 51540 7488 51592 7497
rect 53472 7531 53524 7540
rect 53472 7497 53481 7531
rect 53481 7497 53515 7531
rect 53515 7497 53524 7531
rect 53472 7488 53524 7497
rect 53748 7488 53800 7540
rect 54208 7488 54260 7540
rect 49976 7463 50028 7472
rect 49976 7429 49985 7463
rect 49985 7429 50019 7463
rect 50019 7429 50028 7463
rect 49976 7420 50028 7429
rect 50068 7463 50120 7472
rect 50068 7429 50077 7463
rect 50077 7429 50111 7463
rect 50111 7429 50120 7463
rect 50068 7420 50120 7429
rect 44640 7352 44692 7404
rect 49884 7395 49936 7404
rect 49884 7361 49893 7395
rect 49893 7361 49927 7395
rect 49927 7361 49936 7395
rect 49884 7352 49936 7361
rect 50344 7352 50396 7404
rect 51172 7352 51224 7404
rect 51724 7395 51776 7404
rect 51724 7361 51733 7395
rect 51733 7361 51767 7395
rect 51767 7361 51776 7395
rect 51724 7352 51776 7361
rect 52184 7352 52236 7404
rect 53656 7395 53708 7404
rect 53656 7361 53660 7395
rect 53660 7361 53694 7395
rect 53694 7361 53708 7395
rect 53656 7352 53708 7361
rect 53748 7395 53800 7404
rect 53748 7361 53757 7395
rect 53757 7361 53791 7395
rect 53791 7361 53800 7395
rect 53748 7352 53800 7361
rect 53840 7395 53892 7404
rect 53840 7361 53849 7395
rect 53849 7361 53883 7395
rect 53883 7361 53892 7395
rect 53840 7352 53892 7361
rect 54116 7395 54168 7404
rect 54116 7361 54125 7395
rect 54125 7361 54159 7395
rect 54159 7361 54168 7395
rect 54116 7352 54168 7361
rect 55036 7488 55088 7540
rect 55772 7420 55824 7472
rect 54760 7395 54812 7404
rect 54760 7361 54769 7395
rect 54769 7361 54803 7395
rect 54803 7361 54812 7395
rect 54760 7352 54812 7361
rect 77668 7352 77720 7404
rect 45744 7216 45796 7268
rect 50528 7216 50580 7268
rect 53380 7216 53432 7268
rect 54208 7216 54260 7268
rect 44824 7148 44876 7200
rect 49700 7191 49752 7200
rect 49700 7157 49709 7191
rect 49709 7157 49743 7191
rect 49743 7157 49752 7191
rect 49700 7148 49752 7157
rect 52552 7148 52604 7200
rect 53564 7148 53616 7200
rect 55772 7148 55824 7200
rect 77668 7191 77720 7200
rect 77668 7157 77677 7191
rect 77677 7157 77711 7191
rect 77711 7157 77720 7191
rect 77668 7148 77720 7157
rect 78220 7191 78272 7200
rect 78220 7157 78229 7191
rect 78229 7157 78263 7191
rect 78263 7157 78272 7191
rect 78220 7148 78272 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 30748 6944 30800 6996
rect 31760 6944 31812 6996
rect 33416 6944 33468 6996
rect 34060 6987 34112 6996
rect 34060 6953 34081 6987
rect 34081 6953 34112 6987
rect 34060 6944 34112 6953
rect 44272 6944 44324 6996
rect 46204 6987 46256 6996
rect 46204 6953 46213 6987
rect 46213 6953 46247 6987
rect 46247 6953 46256 6987
rect 46204 6944 46256 6953
rect 46296 6944 46348 6996
rect 46848 6944 46900 6996
rect 50804 6944 50856 6996
rect 54116 6944 54168 6996
rect 29460 6808 29512 6860
rect 31392 6808 31444 6860
rect 31668 6783 31720 6792
rect 31668 6749 31677 6783
rect 31677 6749 31711 6783
rect 31711 6749 31720 6783
rect 31668 6740 31720 6749
rect 31852 6740 31904 6792
rect 33324 6808 33376 6860
rect 33692 6808 33744 6860
rect 37372 6876 37424 6928
rect 38292 6876 38344 6928
rect 34796 6740 34848 6792
rect 35348 6740 35400 6792
rect 33600 6672 33652 6724
rect 33968 6672 34020 6724
rect 35164 6672 35216 6724
rect 37188 6808 37240 6860
rect 36636 6783 36688 6792
rect 36636 6749 36645 6783
rect 36645 6749 36679 6783
rect 36679 6749 36688 6783
rect 36636 6740 36688 6749
rect 38108 6808 38160 6860
rect 37464 6740 37516 6792
rect 38292 6783 38344 6792
rect 38292 6749 38296 6783
rect 38296 6749 38330 6783
rect 38330 6749 38344 6783
rect 38292 6740 38344 6749
rect 39304 6808 39356 6860
rect 41144 6876 41196 6928
rect 44640 6876 44692 6928
rect 45652 6876 45704 6928
rect 33048 6604 33100 6656
rect 33324 6604 33376 6656
rect 34244 6604 34296 6656
rect 35072 6647 35124 6656
rect 35072 6613 35081 6647
rect 35081 6613 35115 6647
rect 35115 6613 35124 6647
rect 35072 6604 35124 6613
rect 35992 6604 36044 6656
rect 36912 6604 36964 6656
rect 38108 6647 38160 6656
rect 38108 6613 38117 6647
rect 38117 6613 38151 6647
rect 38151 6613 38160 6647
rect 38108 6604 38160 6613
rect 38384 6715 38436 6724
rect 38384 6681 38393 6715
rect 38393 6681 38427 6715
rect 38427 6681 38436 6715
rect 38384 6672 38436 6681
rect 38752 6783 38804 6792
rect 38752 6749 38761 6783
rect 38761 6749 38795 6783
rect 38795 6749 38804 6783
rect 38752 6740 38804 6749
rect 40500 6783 40552 6792
rect 40500 6749 40509 6783
rect 40509 6749 40543 6783
rect 40543 6749 40552 6783
rect 40500 6740 40552 6749
rect 41512 6808 41564 6860
rect 40960 6740 41012 6792
rect 42432 6808 42484 6860
rect 43352 6808 43404 6860
rect 45008 6851 45060 6860
rect 45008 6817 45017 6851
rect 45017 6817 45051 6851
rect 45051 6817 45060 6851
rect 45008 6808 45060 6817
rect 45836 6808 45888 6860
rect 46664 6808 46716 6860
rect 40684 6715 40736 6724
rect 40684 6681 40693 6715
rect 40693 6681 40727 6715
rect 40727 6681 40736 6715
rect 40684 6672 40736 6681
rect 40776 6715 40828 6724
rect 40776 6681 40785 6715
rect 40785 6681 40819 6715
rect 40819 6681 40828 6715
rect 40776 6672 40828 6681
rect 41144 6672 41196 6724
rect 42800 6740 42852 6792
rect 46204 6740 46256 6792
rect 46480 6783 46532 6792
rect 46480 6749 46490 6783
rect 46490 6749 46524 6783
rect 46524 6749 46532 6783
rect 46480 6740 46532 6749
rect 49884 6876 49936 6928
rect 49792 6851 49844 6860
rect 49792 6817 49801 6851
rect 49801 6817 49835 6851
rect 49835 6817 49844 6851
rect 49792 6808 49844 6817
rect 50988 6808 51040 6860
rect 51632 6808 51684 6860
rect 43260 6715 43312 6724
rect 43260 6681 43269 6715
rect 43269 6681 43303 6715
rect 43303 6681 43312 6715
rect 43260 6672 43312 6681
rect 44272 6672 44324 6724
rect 45560 6672 45612 6724
rect 45744 6672 45796 6724
rect 41512 6604 41564 6656
rect 41604 6604 41656 6656
rect 44916 6604 44968 6656
rect 45836 6604 45888 6656
rect 46664 6715 46716 6724
rect 46664 6681 46673 6715
rect 46673 6681 46707 6715
rect 46707 6681 46716 6715
rect 46664 6672 46716 6681
rect 46756 6715 46808 6724
rect 46756 6681 46765 6715
rect 46765 6681 46799 6715
rect 46799 6681 46808 6715
rect 46756 6672 46808 6681
rect 47308 6740 47360 6792
rect 49700 6740 49752 6792
rect 50436 6740 50488 6792
rect 77852 6783 77904 6792
rect 77852 6749 77861 6783
rect 77861 6749 77895 6783
rect 77895 6749 77904 6783
rect 77852 6740 77904 6749
rect 51908 6672 51960 6724
rect 49056 6604 49108 6656
rect 49700 6604 49752 6656
rect 78036 6647 78088 6656
rect 78036 6613 78045 6647
rect 78045 6613 78079 6647
rect 78079 6613 78088 6647
rect 78036 6604 78088 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 66314 6502 66366 6554
rect 66378 6502 66430 6554
rect 66442 6502 66494 6554
rect 66506 6502 66558 6554
rect 66570 6502 66622 6554
rect 30104 6443 30156 6452
rect 30104 6409 30113 6443
rect 30113 6409 30147 6443
rect 30147 6409 30156 6443
rect 30104 6400 30156 6409
rect 31484 6400 31536 6452
rect 33508 6400 33560 6452
rect 33876 6400 33928 6452
rect 31392 6332 31444 6384
rect 31760 6332 31812 6384
rect 31484 6307 31536 6316
rect 31484 6273 31493 6307
rect 31493 6273 31527 6307
rect 31527 6273 31536 6307
rect 31484 6264 31536 6273
rect 36636 6400 36688 6452
rect 40960 6400 41012 6452
rect 41696 6400 41748 6452
rect 42432 6400 42484 6452
rect 35072 6375 35124 6384
rect 35072 6341 35081 6375
rect 35081 6341 35115 6375
rect 35115 6341 35124 6375
rect 35072 6332 35124 6341
rect 35164 6332 35216 6384
rect 32956 6264 33008 6316
rect 29460 6196 29512 6248
rect 33324 6307 33376 6316
rect 33324 6273 33333 6307
rect 33333 6273 33367 6307
rect 33367 6273 33376 6307
rect 33324 6264 33376 6273
rect 33508 6307 33560 6316
rect 33508 6273 33522 6307
rect 33522 6273 33556 6307
rect 33556 6273 33560 6307
rect 33508 6264 33560 6273
rect 34796 6307 34848 6316
rect 34796 6273 34805 6307
rect 34805 6273 34839 6307
rect 34839 6273 34848 6307
rect 34796 6264 34848 6273
rect 36636 6264 36688 6316
rect 38752 6332 38804 6384
rect 41144 6332 41196 6384
rect 41604 6375 41656 6384
rect 41604 6341 41613 6375
rect 41613 6341 41647 6375
rect 41647 6341 41656 6375
rect 41604 6332 41656 6341
rect 38108 6264 38160 6316
rect 43260 6400 43312 6452
rect 44180 6400 44232 6452
rect 44456 6400 44508 6452
rect 43076 6332 43128 6384
rect 44916 6400 44968 6452
rect 45008 6400 45060 6452
rect 44824 6375 44876 6384
rect 44824 6341 44833 6375
rect 44833 6341 44867 6375
rect 44867 6341 44876 6375
rect 44824 6332 44876 6341
rect 43352 6264 43404 6316
rect 44456 6307 44508 6316
rect 44456 6273 44465 6307
rect 44465 6273 44499 6307
rect 44499 6273 44508 6307
rect 44456 6264 44508 6273
rect 44640 6307 44692 6316
rect 44640 6273 44647 6307
rect 44647 6273 44692 6307
rect 44640 6264 44692 6273
rect 45560 6264 45612 6316
rect 47308 6400 47360 6452
rect 46572 6332 46624 6384
rect 47768 6332 47820 6384
rect 49056 6375 49108 6384
rect 49056 6341 49065 6375
rect 49065 6341 49099 6375
rect 49099 6341 49108 6375
rect 49056 6332 49108 6341
rect 49700 6375 49752 6384
rect 49700 6341 49709 6375
rect 49709 6341 49743 6375
rect 49743 6341 49752 6375
rect 49700 6332 49752 6341
rect 50436 6400 50488 6452
rect 55128 6400 55180 6452
rect 49976 6332 50028 6384
rect 51632 6264 51684 6316
rect 53656 6264 53708 6316
rect 34428 6196 34480 6248
rect 31208 6060 31260 6112
rect 32956 6060 33008 6112
rect 34152 6060 34204 6112
rect 36912 6196 36964 6248
rect 38200 6196 38252 6248
rect 39764 6239 39816 6248
rect 39764 6205 39773 6239
rect 39773 6205 39807 6239
rect 39807 6205 39816 6239
rect 39764 6196 39816 6205
rect 37556 6128 37608 6180
rect 38476 6128 38528 6180
rect 41052 6196 41104 6248
rect 41144 6196 41196 6248
rect 42800 6196 42852 6248
rect 45100 6196 45152 6248
rect 42248 6128 42300 6180
rect 46112 6196 46164 6248
rect 46756 6196 46808 6248
rect 48044 6196 48096 6248
rect 50712 6196 50764 6248
rect 53288 6196 53340 6248
rect 54024 6264 54076 6316
rect 54208 6264 54260 6316
rect 36084 6060 36136 6112
rect 38108 6060 38160 6112
rect 41512 6060 41564 6112
rect 42524 6060 42576 6112
rect 43720 6060 43772 6112
rect 46296 6103 46348 6112
rect 46296 6069 46305 6103
rect 46305 6069 46339 6103
rect 46339 6069 46348 6103
rect 46296 6060 46348 6069
rect 46480 6060 46532 6112
rect 46756 6060 46808 6112
rect 49516 6060 49568 6112
rect 52460 6060 52512 6112
rect 52828 6103 52880 6112
rect 52828 6069 52837 6103
rect 52837 6069 52871 6103
rect 52871 6069 52880 6103
rect 52828 6060 52880 6069
rect 53656 6060 53708 6112
rect 53748 6060 53800 6112
rect 78036 6307 78088 6316
rect 78036 6273 78045 6307
rect 78045 6273 78079 6307
rect 78079 6273 78088 6307
rect 78036 6264 78088 6273
rect 78220 6171 78272 6180
rect 78220 6137 78229 6171
rect 78229 6137 78263 6171
rect 78263 6137 78272 6171
rect 78220 6128 78272 6137
rect 55312 6060 55364 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 31852 5856 31904 5908
rect 34244 5856 34296 5908
rect 32036 5788 32088 5840
rect 35348 5899 35400 5908
rect 35348 5865 35357 5899
rect 35357 5865 35391 5899
rect 35391 5865 35400 5899
rect 35348 5856 35400 5865
rect 36820 5856 36872 5908
rect 39764 5856 39816 5908
rect 44364 5856 44416 5908
rect 46112 5856 46164 5908
rect 50068 5856 50120 5908
rect 50344 5856 50396 5908
rect 50988 5856 51040 5908
rect 53288 5899 53340 5908
rect 53288 5865 53297 5899
rect 53297 5865 53331 5899
rect 53331 5865 53340 5899
rect 53288 5856 53340 5865
rect 29460 5720 29512 5772
rect 30288 5720 30340 5772
rect 33048 5720 33100 5772
rect 31760 5652 31812 5704
rect 33508 5652 33560 5704
rect 34060 5695 34112 5704
rect 34060 5661 34068 5695
rect 34068 5661 34102 5695
rect 34102 5661 34112 5695
rect 34060 5652 34112 5661
rect 34152 5695 34204 5704
rect 34152 5661 34161 5695
rect 34161 5661 34195 5695
rect 34195 5661 34204 5695
rect 34152 5652 34204 5661
rect 34612 5652 34664 5704
rect 34796 5695 34848 5704
rect 34796 5661 34806 5695
rect 34806 5661 34840 5695
rect 34840 5661 34848 5695
rect 34796 5652 34848 5661
rect 30656 5627 30708 5636
rect 30656 5593 30665 5627
rect 30665 5593 30699 5627
rect 30699 5593 30708 5627
rect 30656 5584 30708 5593
rect 33324 5584 33376 5636
rect 34520 5584 34572 5636
rect 34888 5584 34940 5636
rect 35992 5788 36044 5840
rect 36176 5788 36228 5840
rect 37464 5788 37516 5840
rect 41420 5788 41472 5840
rect 36084 5720 36136 5772
rect 38108 5763 38160 5772
rect 38108 5729 38117 5763
rect 38117 5729 38151 5763
rect 38151 5729 38160 5763
rect 38108 5720 38160 5729
rect 35164 5695 35216 5704
rect 35164 5661 35178 5695
rect 35178 5661 35212 5695
rect 35212 5661 35216 5695
rect 35164 5652 35216 5661
rect 36636 5695 36688 5704
rect 36636 5661 36645 5695
rect 36645 5661 36679 5695
rect 36679 5661 36688 5695
rect 36636 5652 36688 5661
rect 36820 5695 36872 5704
rect 36820 5661 36827 5695
rect 36827 5661 36872 5695
rect 36820 5652 36872 5661
rect 36912 5695 36964 5704
rect 36912 5661 36921 5695
rect 36921 5661 36955 5695
rect 36955 5661 36964 5695
rect 36912 5652 36964 5661
rect 37464 5652 37516 5704
rect 40684 5652 40736 5704
rect 35440 5584 35492 5636
rect 33140 5516 33192 5568
rect 34612 5516 34664 5568
rect 37372 5584 37424 5636
rect 37188 5516 37240 5568
rect 37464 5516 37516 5568
rect 41236 5584 41288 5636
rect 41696 5695 41748 5704
rect 41696 5661 41705 5695
rect 41705 5661 41739 5695
rect 41739 5661 41748 5695
rect 41696 5652 41748 5661
rect 41880 5695 41932 5704
rect 46480 5763 46532 5772
rect 46480 5729 46489 5763
rect 46489 5729 46523 5763
rect 46523 5729 46532 5763
rect 46480 5720 46532 5729
rect 46756 5763 46808 5772
rect 46756 5729 46765 5763
rect 46765 5729 46799 5763
rect 46799 5729 46808 5763
rect 46756 5720 46808 5729
rect 51448 5788 51500 5840
rect 41880 5661 41925 5695
rect 41925 5661 41932 5695
rect 41880 5652 41932 5661
rect 46572 5584 46624 5636
rect 41144 5516 41196 5568
rect 41420 5559 41472 5568
rect 41420 5525 41429 5559
rect 41429 5525 41463 5559
rect 41463 5525 41472 5559
rect 41420 5516 41472 5525
rect 41788 5516 41840 5568
rect 46204 5516 46256 5568
rect 50344 5695 50396 5704
rect 50344 5661 50348 5695
rect 50348 5661 50382 5695
rect 50382 5661 50396 5695
rect 50344 5652 50396 5661
rect 50436 5695 50488 5704
rect 50436 5661 50445 5695
rect 50445 5661 50479 5695
rect 50479 5661 50488 5695
rect 50436 5652 50488 5661
rect 50712 5695 50764 5704
rect 50712 5661 50720 5695
rect 50720 5661 50754 5695
rect 50754 5661 50764 5695
rect 50712 5652 50764 5661
rect 50804 5695 50856 5704
rect 50804 5661 50813 5695
rect 50813 5661 50847 5695
rect 50847 5661 50856 5695
rect 50804 5652 50856 5661
rect 51080 5720 51132 5772
rect 51172 5695 51224 5704
rect 51172 5661 51181 5695
rect 51181 5661 51215 5695
rect 51215 5661 51224 5695
rect 51172 5652 51224 5661
rect 50068 5584 50120 5636
rect 49516 5559 49568 5568
rect 49516 5525 49525 5559
rect 49525 5525 49559 5559
rect 49559 5525 49568 5559
rect 49516 5516 49568 5525
rect 49700 5516 49752 5568
rect 54024 5720 54076 5772
rect 55036 5720 55088 5772
rect 55588 5720 55640 5772
rect 51448 5559 51500 5568
rect 51448 5525 51457 5559
rect 51457 5525 51491 5559
rect 51491 5525 51500 5559
rect 51448 5516 51500 5525
rect 52920 5652 52972 5704
rect 53380 5695 53432 5704
rect 53380 5661 53389 5695
rect 53389 5661 53423 5695
rect 53423 5661 53432 5695
rect 53380 5652 53432 5661
rect 51724 5584 51776 5636
rect 52092 5516 52144 5568
rect 53564 5584 53616 5636
rect 53748 5516 53800 5568
rect 55404 5627 55456 5636
rect 55404 5593 55413 5627
rect 55413 5593 55447 5627
rect 55447 5593 55456 5627
rect 55404 5584 55456 5593
rect 55772 5516 55824 5568
rect 77668 5559 77720 5568
rect 77668 5525 77677 5559
rect 77677 5525 77711 5559
rect 77711 5525 77720 5559
rect 77668 5516 77720 5525
rect 78404 5559 78456 5568
rect 78404 5525 78413 5559
rect 78413 5525 78447 5559
rect 78447 5525 78456 5559
rect 78404 5516 78456 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 66314 5414 66366 5466
rect 66378 5414 66430 5466
rect 66442 5414 66494 5466
rect 66506 5414 66558 5466
rect 66570 5414 66622 5466
rect 30656 5312 30708 5364
rect 36268 5312 36320 5364
rect 36544 5312 36596 5364
rect 36912 5312 36964 5364
rect 42616 5312 42668 5364
rect 30932 5176 30984 5228
rect 31208 5219 31260 5228
rect 31208 5185 31217 5219
rect 31217 5185 31251 5219
rect 31251 5185 31260 5219
rect 31208 5176 31260 5185
rect 32036 5176 32088 5228
rect 33140 5219 33192 5228
rect 33140 5185 33149 5219
rect 33149 5185 33183 5219
rect 33183 5185 33192 5219
rect 33140 5176 33192 5185
rect 33692 5244 33744 5296
rect 34428 5244 34480 5296
rect 34888 5219 34940 5228
rect 34888 5185 34897 5219
rect 34897 5185 34931 5219
rect 34931 5185 34940 5219
rect 34888 5176 34940 5185
rect 35164 5176 35216 5228
rect 36176 5176 36228 5228
rect 36360 5219 36412 5228
rect 36360 5185 36369 5219
rect 36369 5185 36403 5219
rect 36403 5185 36412 5219
rect 36360 5176 36412 5185
rect 36544 5176 36596 5228
rect 38384 5244 38436 5296
rect 37096 5108 37148 5160
rect 35992 5083 36044 5092
rect 35992 5049 36001 5083
rect 36001 5049 36035 5083
rect 36035 5049 36044 5083
rect 37372 5176 37424 5228
rect 37464 5219 37516 5228
rect 37464 5185 37473 5219
rect 37473 5185 37507 5219
rect 37507 5185 37516 5219
rect 37464 5176 37516 5185
rect 41880 5244 41932 5296
rect 42892 5287 42944 5296
rect 42892 5253 42901 5287
rect 42901 5253 42935 5287
rect 42935 5253 42944 5287
rect 42892 5244 42944 5253
rect 44180 5312 44232 5364
rect 53104 5355 53156 5364
rect 53104 5321 53113 5355
rect 53113 5321 53147 5355
rect 53147 5321 53156 5355
rect 53104 5312 53156 5321
rect 41788 5176 41840 5228
rect 43076 5219 43128 5228
rect 44548 5244 44600 5296
rect 43076 5185 43121 5219
rect 43121 5185 43128 5219
rect 43076 5176 43128 5185
rect 43904 5176 43956 5228
rect 49516 5176 49568 5228
rect 49700 5219 49752 5228
rect 49700 5185 49709 5219
rect 49709 5185 49743 5219
rect 49743 5185 49752 5219
rect 49700 5176 49752 5185
rect 50988 5176 51040 5228
rect 45652 5108 45704 5160
rect 49792 5108 49844 5160
rect 35992 5040 36044 5049
rect 32312 4972 32364 5024
rect 35532 4972 35584 5024
rect 36452 4972 36504 5024
rect 37188 4972 37240 5024
rect 37556 4972 37608 5024
rect 43444 4972 43496 5024
rect 46296 4972 46348 5024
rect 47400 4972 47452 5024
rect 49516 5015 49568 5024
rect 49516 4981 49525 5015
rect 49525 4981 49559 5015
rect 49559 4981 49568 5015
rect 49516 4972 49568 4981
rect 51448 5244 51500 5296
rect 51908 5219 51960 5228
rect 51908 5185 51917 5219
rect 51917 5185 51951 5219
rect 51951 5185 51960 5219
rect 51908 5176 51960 5185
rect 52828 5176 52880 5228
rect 55128 5219 55180 5228
rect 55128 5185 55137 5219
rect 55137 5185 55171 5219
rect 55171 5185 55180 5219
rect 55128 5176 55180 5185
rect 78312 5219 78364 5228
rect 78312 5185 78321 5219
rect 78321 5185 78355 5219
rect 78355 5185 78364 5219
rect 78312 5176 78364 5185
rect 51724 5151 51776 5160
rect 51724 5117 51733 5151
rect 51733 5117 51767 5151
rect 51767 5117 51776 5151
rect 51724 5108 51776 5117
rect 52092 5108 52144 5160
rect 53380 5108 53432 5160
rect 56048 5108 56100 5160
rect 55404 5040 55456 5092
rect 52552 4972 52604 5024
rect 78128 5015 78180 5024
rect 78128 4981 78137 5015
rect 78137 4981 78171 5015
rect 78171 4981 78180 5015
rect 78128 4972 78180 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 30012 4768 30064 4820
rect 30288 4632 30340 4684
rect 32312 4675 32364 4684
rect 32312 4641 32321 4675
rect 32321 4641 32355 4675
rect 32355 4641 32364 4675
rect 32312 4632 32364 4641
rect 30012 4607 30064 4616
rect 30012 4573 30021 4607
rect 30021 4573 30055 4607
rect 30055 4573 30064 4607
rect 30012 4564 30064 4573
rect 31484 4564 31536 4616
rect 33600 4496 33652 4548
rect 31668 4428 31720 4480
rect 43628 4768 43680 4820
rect 44732 4768 44784 4820
rect 44824 4768 44876 4820
rect 34428 4700 34480 4752
rect 34060 4632 34112 4684
rect 33784 4564 33836 4616
rect 35256 4471 35308 4480
rect 35256 4437 35265 4471
rect 35265 4437 35299 4471
rect 35299 4437 35308 4471
rect 35256 4428 35308 4437
rect 35532 4607 35584 4616
rect 35532 4573 35541 4607
rect 35541 4573 35575 4607
rect 35575 4573 35584 4607
rect 35532 4564 35584 4573
rect 38384 4700 38436 4752
rect 41328 4700 41380 4752
rect 41972 4700 42024 4752
rect 37188 4675 37240 4684
rect 37188 4641 37197 4675
rect 37197 4641 37231 4675
rect 37231 4641 37240 4675
rect 37188 4632 37240 4641
rect 40776 4632 40828 4684
rect 44272 4632 44324 4684
rect 36360 4564 36412 4616
rect 35992 4496 36044 4548
rect 36084 4496 36136 4548
rect 39856 4607 39908 4616
rect 39856 4573 39865 4607
rect 39865 4573 39899 4607
rect 39899 4573 39908 4607
rect 39856 4564 39908 4573
rect 41236 4564 41288 4616
rect 42800 4607 42852 4616
rect 42800 4573 42809 4607
rect 42809 4573 42843 4607
rect 42843 4573 42852 4607
rect 42800 4564 42852 4573
rect 44824 4564 44876 4616
rect 45836 4632 45888 4684
rect 46848 4632 46900 4684
rect 37648 4496 37700 4548
rect 40132 4539 40184 4548
rect 40132 4505 40141 4539
rect 40141 4505 40175 4539
rect 40175 4505 40184 4539
rect 40132 4496 40184 4505
rect 36360 4428 36412 4480
rect 43076 4539 43128 4548
rect 43076 4505 43085 4539
rect 43085 4505 43119 4539
rect 43119 4505 43128 4539
rect 43076 4496 43128 4505
rect 45560 4564 45612 4616
rect 46112 4564 46164 4616
rect 47400 4811 47452 4820
rect 47400 4777 47409 4811
rect 47409 4777 47443 4811
rect 47443 4777 47452 4811
rect 47400 4768 47452 4777
rect 49516 4768 49568 4820
rect 53564 4768 53616 4820
rect 47308 4607 47360 4616
rect 47308 4573 47317 4607
rect 47317 4573 47351 4607
rect 47351 4573 47360 4607
rect 47308 4564 47360 4573
rect 52552 4700 52604 4752
rect 50988 4632 51040 4684
rect 52092 4632 52144 4684
rect 47676 4607 47728 4616
rect 47676 4573 47685 4607
rect 47685 4573 47719 4607
rect 47719 4573 47728 4607
rect 47676 4564 47728 4573
rect 52000 4564 52052 4616
rect 54760 4632 54812 4684
rect 53656 4607 53708 4616
rect 53656 4573 53665 4607
rect 53665 4573 53699 4607
rect 53699 4573 53708 4607
rect 53656 4564 53708 4573
rect 42984 4428 43036 4480
rect 44732 4428 44784 4480
rect 46848 4539 46900 4548
rect 46848 4505 46857 4539
rect 46857 4505 46891 4539
rect 46891 4505 46900 4539
rect 46848 4496 46900 4505
rect 45560 4471 45612 4480
rect 45560 4437 45569 4471
rect 45569 4437 45603 4471
rect 45603 4437 45612 4471
rect 45560 4428 45612 4437
rect 45652 4428 45704 4480
rect 46756 4428 46808 4480
rect 49976 4496 50028 4548
rect 50344 4496 50396 4548
rect 51540 4496 51592 4548
rect 55036 4564 55088 4616
rect 78496 4607 78548 4616
rect 78496 4573 78505 4607
rect 78505 4573 78539 4607
rect 78539 4573 78548 4607
rect 78496 4564 78548 4573
rect 49056 4428 49108 4480
rect 78312 4471 78364 4480
rect 78312 4437 78321 4471
rect 78321 4437 78355 4471
rect 78355 4437 78364 4471
rect 78312 4428 78364 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 66314 4326 66366 4378
rect 66378 4326 66430 4378
rect 66442 4326 66494 4378
rect 66506 4326 66558 4378
rect 66570 4326 66622 4378
rect 33600 4156 33652 4208
rect 35992 4224 36044 4276
rect 37832 4224 37884 4276
rect 40132 4224 40184 4276
rect 43076 4224 43128 4276
rect 47308 4224 47360 4276
rect 36268 4156 36320 4208
rect 37648 4156 37700 4208
rect 38200 4156 38252 4208
rect 39580 4156 39632 4208
rect 30840 4088 30892 4140
rect 36084 4131 36136 4140
rect 36084 4097 36093 4131
rect 36093 4097 36127 4131
rect 36127 4097 36136 4131
rect 36084 4088 36136 4097
rect 36360 4131 36412 4140
rect 36360 4097 36369 4131
rect 36369 4097 36403 4131
rect 36403 4097 36412 4131
rect 36360 4088 36412 4097
rect 36452 4131 36504 4140
rect 36452 4097 36461 4131
rect 36461 4097 36495 4131
rect 36495 4097 36504 4131
rect 36452 4088 36504 4097
rect 41144 4088 41196 4140
rect 41788 4156 41840 4208
rect 41972 4199 42024 4208
rect 41972 4165 41981 4199
rect 41981 4165 42015 4199
rect 42015 4165 42024 4199
rect 41972 4156 42024 4165
rect 42616 4156 42668 4208
rect 47768 4156 47820 4208
rect 34060 4020 34112 4072
rect 35256 4020 35308 4072
rect 19708 3884 19760 3936
rect 31852 3884 31904 3936
rect 31944 3927 31996 3936
rect 31944 3893 31953 3927
rect 31953 3893 31987 3927
rect 31987 3893 31996 3927
rect 31944 3884 31996 3893
rect 36176 3927 36228 3936
rect 36176 3893 36185 3927
rect 36185 3893 36219 3927
rect 36219 3893 36228 3927
rect 36176 3884 36228 3893
rect 37096 4020 37148 4072
rect 37556 3952 37608 4004
rect 40868 3995 40920 4004
rect 40868 3961 40877 3995
rect 40877 3961 40911 3995
rect 40911 3961 40920 3995
rect 40868 3952 40920 3961
rect 38844 3884 38896 3936
rect 39580 3884 39632 3936
rect 40776 3884 40828 3936
rect 42892 4088 42944 4140
rect 43444 4088 43496 4140
rect 44732 4131 44784 4140
rect 44732 4097 44741 4131
rect 44741 4097 44775 4131
rect 44775 4097 44784 4131
rect 44732 4088 44784 4097
rect 45560 4088 45612 4140
rect 45652 4131 45704 4140
rect 45652 4097 45661 4131
rect 45661 4097 45695 4131
rect 45695 4097 45704 4131
rect 45652 4088 45704 4097
rect 54024 4088 54076 4140
rect 68192 4088 68244 4140
rect 47124 4020 47176 4072
rect 47676 4020 47728 4072
rect 49056 4063 49108 4072
rect 49056 4029 49065 4063
rect 49065 4029 49099 4063
rect 49099 4029 49108 4063
rect 49056 4020 49108 4029
rect 51080 4020 51132 4072
rect 52092 4020 52144 4072
rect 59360 4020 59412 4072
rect 78312 4020 78364 4072
rect 43720 3995 43772 4004
rect 43720 3961 43729 3995
rect 43729 3961 43763 3995
rect 43763 3961 43772 3995
rect 43720 3952 43772 3961
rect 46296 3952 46348 4004
rect 51448 3952 51500 4004
rect 58992 3952 59044 4004
rect 41420 3884 41472 3936
rect 41512 3927 41564 3936
rect 41512 3893 41521 3927
rect 41521 3893 41555 3927
rect 41555 3893 41564 3927
rect 41512 3884 41564 3893
rect 45284 3884 45336 3936
rect 56416 3927 56468 3936
rect 56416 3893 56425 3927
rect 56425 3893 56459 3927
rect 56459 3893 56468 3927
rect 56416 3884 56468 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 30012 3723 30064 3732
rect 30012 3689 30021 3723
rect 30021 3689 30055 3723
rect 30055 3689 30064 3723
rect 30012 3680 30064 3689
rect 31944 3680 31996 3732
rect 30196 3587 30248 3596
rect 30196 3553 30205 3587
rect 30205 3553 30239 3587
rect 30239 3553 30248 3587
rect 30196 3544 30248 3553
rect 31760 3612 31812 3664
rect 38200 3612 38252 3664
rect 42892 3655 42944 3664
rect 42892 3621 42901 3655
rect 42901 3621 42935 3655
rect 42935 3621 42944 3655
rect 42892 3612 42944 3621
rect 42984 3612 43036 3664
rect 43260 3612 43312 3664
rect 44272 3612 44324 3664
rect 44548 3612 44600 3664
rect 46756 3723 46808 3732
rect 46756 3689 46765 3723
rect 46765 3689 46799 3723
rect 46799 3689 46808 3723
rect 46756 3680 46808 3689
rect 50344 3723 50396 3732
rect 50344 3689 50353 3723
rect 50353 3689 50387 3723
rect 50387 3689 50396 3723
rect 50344 3680 50396 3689
rect 51356 3680 51408 3732
rect 59360 3723 59412 3732
rect 55312 3612 55364 3664
rect 42800 3544 42852 3596
rect 44824 3544 44876 3596
rect 45008 3587 45060 3596
rect 45008 3553 45017 3587
rect 45017 3553 45051 3587
rect 45051 3553 45060 3587
rect 45008 3544 45060 3553
rect 45284 3587 45336 3596
rect 45284 3553 45293 3587
rect 45293 3553 45327 3587
rect 45327 3553 45336 3587
rect 45284 3544 45336 3553
rect 55404 3544 55456 3596
rect 56416 3544 56468 3596
rect 57796 3612 57848 3664
rect 59360 3689 59369 3723
rect 59369 3689 59403 3723
rect 59403 3689 59412 3723
rect 59360 3680 59412 3689
rect 72608 3723 72660 3732
rect 72608 3689 72617 3723
rect 72617 3689 72651 3723
rect 72651 3689 72660 3723
rect 72608 3680 72660 3689
rect 68928 3612 68980 3664
rect 77668 3612 77720 3664
rect 31852 3476 31904 3528
rect 38936 3451 38988 3460
rect 38936 3417 38945 3451
rect 38945 3417 38979 3451
rect 38979 3417 38988 3451
rect 38936 3408 38988 3417
rect 41420 3451 41472 3460
rect 41420 3417 41429 3451
rect 41429 3417 41463 3451
rect 41463 3417 41472 3451
rect 41420 3408 41472 3417
rect 42708 3408 42760 3460
rect 31944 3383 31996 3392
rect 31944 3349 31953 3383
rect 31953 3349 31987 3383
rect 31987 3349 31996 3383
rect 31944 3340 31996 3349
rect 44916 3476 44968 3528
rect 52920 3476 52972 3528
rect 54300 3476 54352 3528
rect 55496 3476 55548 3528
rect 57704 3544 57756 3596
rect 43628 3451 43680 3460
rect 43628 3417 43637 3451
rect 43637 3417 43671 3451
rect 43671 3417 43680 3451
rect 43628 3408 43680 3417
rect 43904 3408 43956 3460
rect 44548 3408 44600 3460
rect 47768 3408 47820 3460
rect 50344 3408 50396 3460
rect 58164 3519 58216 3528
rect 58164 3485 58173 3519
rect 58173 3485 58207 3519
rect 58207 3485 58216 3519
rect 58164 3476 58216 3485
rect 58256 3408 58308 3460
rect 74448 3544 74500 3596
rect 58992 3519 59044 3528
rect 58992 3485 59001 3519
rect 59001 3485 59035 3519
rect 59035 3485 59044 3519
rect 58992 3476 59044 3485
rect 68468 3476 68520 3528
rect 72424 3476 72476 3528
rect 73528 3476 73580 3528
rect 76196 3476 76248 3528
rect 50804 3383 50856 3392
rect 50804 3349 50813 3383
rect 50813 3349 50847 3383
rect 50847 3349 50856 3383
rect 50804 3340 50856 3349
rect 50988 3383 51040 3392
rect 50988 3349 51015 3383
rect 51015 3349 51040 3383
rect 50988 3340 51040 3349
rect 56784 3383 56836 3392
rect 56784 3349 56793 3383
rect 56793 3349 56827 3383
rect 56827 3349 56836 3383
rect 56784 3340 56836 3349
rect 56968 3383 57020 3392
rect 56968 3349 56977 3383
rect 56977 3349 57011 3383
rect 57011 3349 57020 3383
rect 56968 3340 57020 3349
rect 57796 3340 57848 3392
rect 58440 3340 58492 3392
rect 72148 3383 72200 3392
rect 72148 3349 72157 3383
rect 72157 3349 72191 3383
rect 72191 3349 72200 3383
rect 72148 3340 72200 3349
rect 72516 3408 72568 3460
rect 78128 3408 78180 3460
rect 72884 3383 72936 3392
rect 72884 3349 72893 3383
rect 72893 3349 72927 3383
rect 72927 3349 72936 3383
rect 72884 3340 72936 3349
rect 73068 3340 73120 3392
rect 77760 3340 77812 3392
rect 77944 3340 77996 3392
rect 78496 3383 78548 3392
rect 78496 3349 78505 3383
rect 78505 3349 78539 3383
rect 78539 3349 78548 3383
rect 78496 3340 78548 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 66314 3238 66366 3290
rect 66378 3238 66430 3290
rect 66442 3238 66494 3290
rect 66506 3238 66558 3290
rect 66570 3238 66622 3290
rect 31852 3179 31904 3188
rect 31852 3145 31861 3179
rect 31861 3145 31895 3179
rect 31895 3145 31904 3179
rect 31852 3136 31904 3145
rect 35992 3136 36044 3188
rect 31944 3000 31996 3052
rect 36268 3068 36320 3120
rect 44272 3136 44324 3188
rect 54300 3179 54352 3188
rect 39856 3068 39908 3120
rect 38660 3000 38712 3052
rect 44916 3068 44968 3120
rect 50804 3111 50856 3120
rect 54300 3145 54309 3179
rect 54309 3145 54343 3179
rect 54343 3145 54352 3179
rect 54300 3136 54352 3145
rect 50804 3077 50822 3111
rect 50822 3077 50856 3111
rect 50804 3068 50856 3077
rect 54024 3111 54076 3120
rect 54024 3077 54033 3111
rect 54033 3077 54067 3111
rect 54067 3077 54076 3111
rect 54024 3068 54076 3077
rect 55496 3068 55548 3120
rect 58256 3179 58308 3188
rect 58256 3145 58265 3179
rect 58265 3145 58299 3179
rect 58299 3145 58308 3179
rect 58256 3136 58308 3145
rect 56784 3068 56836 3120
rect 36176 2932 36228 2984
rect 37096 2975 37148 2984
rect 37096 2941 37105 2975
rect 37105 2941 37139 2975
rect 37139 2941 37148 2975
rect 37096 2932 37148 2941
rect 40040 3000 40092 3052
rect 44180 3000 44232 3052
rect 44824 3043 44876 3052
rect 44824 3009 44833 3043
rect 44833 3009 44867 3043
rect 44867 3009 44876 3043
rect 44824 3000 44876 3009
rect 45560 3043 45612 3052
rect 45560 3009 45569 3043
rect 45569 3009 45603 3043
rect 45603 3009 45612 3043
rect 45560 3000 45612 3009
rect 39488 2864 39540 2916
rect 51080 3043 51132 3052
rect 51080 3009 51089 3043
rect 51089 3009 51123 3043
rect 51123 3009 51132 3043
rect 51080 3000 51132 3009
rect 51448 3043 51500 3052
rect 51448 3009 51457 3043
rect 51457 3009 51491 3043
rect 51491 3009 51500 3043
rect 51448 3000 51500 3009
rect 32956 2796 33008 2848
rect 39396 2796 39448 2848
rect 41420 2839 41472 2848
rect 41420 2805 41429 2839
rect 41429 2805 41463 2839
rect 41463 2805 41472 2839
rect 41420 2796 41472 2805
rect 43352 2839 43404 2848
rect 43352 2805 43361 2839
rect 43361 2805 43395 2839
rect 43395 2805 43404 2839
rect 43352 2796 43404 2805
rect 43536 2796 43588 2848
rect 56048 2975 56100 2984
rect 56048 2941 56057 2975
rect 56057 2941 56091 2975
rect 56091 2941 56100 2975
rect 56048 2932 56100 2941
rect 49792 2864 49844 2916
rect 45008 2796 45060 2848
rect 45836 2796 45888 2848
rect 46480 2796 46532 2848
rect 47124 2796 47176 2848
rect 47768 2839 47820 2848
rect 47768 2805 47777 2839
rect 47777 2805 47811 2839
rect 47811 2805 47820 2839
rect 47768 2796 47820 2805
rect 49056 2796 49108 2848
rect 49700 2839 49752 2848
rect 49700 2805 49709 2839
rect 49709 2805 49743 2839
rect 49743 2805 49752 2839
rect 49700 2796 49752 2805
rect 51264 2796 51316 2848
rect 51632 2839 51684 2848
rect 51632 2805 51641 2839
rect 51641 2805 51675 2839
rect 51675 2805 51684 2839
rect 51632 2796 51684 2805
rect 53564 2796 53616 2848
rect 54116 2839 54168 2848
rect 54116 2805 54125 2839
rect 54125 2805 54159 2839
rect 54159 2805 54168 2839
rect 54116 2796 54168 2805
rect 55312 2796 55364 2848
rect 56324 3000 56376 3052
rect 57796 3000 57848 3052
rect 58716 3043 58768 3052
rect 58716 3009 58725 3043
rect 58725 3009 58759 3043
rect 58759 3009 58768 3043
rect 58716 3000 58768 3009
rect 68928 3179 68980 3188
rect 68928 3145 68937 3179
rect 68937 3145 68971 3179
rect 68971 3145 68980 3179
rect 68928 3136 68980 3145
rect 56600 2932 56652 2984
rect 58348 2975 58400 2984
rect 58348 2941 58357 2975
rect 58357 2941 58391 2975
rect 58391 2941 58400 2975
rect 58348 2932 58400 2941
rect 58440 2975 58492 2984
rect 58440 2941 58449 2975
rect 58449 2941 58483 2975
rect 58483 2941 58492 2975
rect 58440 2932 58492 2941
rect 58808 2975 58860 2984
rect 58808 2941 58817 2975
rect 58817 2941 58851 2975
rect 58851 2941 58860 2975
rect 58808 2932 58860 2941
rect 59820 3043 59872 3052
rect 59820 3009 59829 3043
rect 59829 3009 59863 3043
rect 59863 3009 59872 3043
rect 59820 3000 59872 3009
rect 66444 3068 66496 3120
rect 72424 3136 72476 3188
rect 72516 3179 72568 3188
rect 72516 3145 72525 3179
rect 72525 3145 72559 3179
rect 72559 3145 72568 3179
rect 72516 3136 72568 3145
rect 72608 3179 72660 3188
rect 72608 3145 72617 3179
rect 72617 3145 72651 3179
rect 72651 3145 72660 3179
rect 72608 3136 72660 3145
rect 73528 3179 73580 3188
rect 73528 3145 73537 3179
rect 73537 3145 73571 3179
rect 73571 3145 73580 3179
rect 73528 3136 73580 3145
rect 72148 3068 72200 3120
rect 77392 3068 77444 3120
rect 59636 2932 59688 2984
rect 59728 2975 59780 2984
rect 59728 2941 59737 2975
rect 59737 2941 59771 2975
rect 59771 2941 59780 2975
rect 59728 2932 59780 2941
rect 60004 2975 60056 2984
rect 60004 2941 60013 2975
rect 60013 2941 60047 2975
rect 60047 2941 60056 2975
rect 60004 2932 60056 2941
rect 66536 2975 66588 2984
rect 66536 2941 66545 2975
rect 66545 2941 66579 2975
rect 66579 2941 66588 2975
rect 66536 2932 66588 2941
rect 68192 3043 68244 3052
rect 68192 3009 68201 3043
rect 68201 3009 68235 3043
rect 68235 3009 68244 3043
rect 68192 3000 68244 3009
rect 68928 3000 68980 3052
rect 69020 3000 69072 3052
rect 71136 3043 71188 3052
rect 71136 3009 71145 3043
rect 71145 3009 71179 3043
rect 71179 3009 71188 3043
rect 71136 3000 71188 3009
rect 71228 3000 71280 3052
rect 72424 3000 72476 3052
rect 69756 2932 69808 2984
rect 72240 2975 72292 2984
rect 72240 2941 72249 2975
rect 72249 2941 72283 2975
rect 72283 2941 72292 2975
rect 72240 2932 72292 2941
rect 72516 2932 72568 2984
rect 73988 3000 74040 3052
rect 74172 3043 74224 3052
rect 74172 3009 74181 3043
rect 74181 3009 74215 3043
rect 74215 3009 74224 3043
rect 74172 3000 74224 3009
rect 76196 3043 76248 3052
rect 76196 3009 76205 3043
rect 76205 3009 76239 3043
rect 76239 3009 76248 3043
rect 76196 3000 76248 3009
rect 77852 3043 77904 3052
rect 77852 3009 77853 3043
rect 77853 3009 77887 3043
rect 77887 3009 77904 3043
rect 77852 3000 77904 3009
rect 78496 3000 78548 3052
rect 79232 3000 79284 3052
rect 57428 2839 57480 2848
rect 57428 2805 57437 2839
rect 57437 2805 57471 2839
rect 57471 2805 57480 2839
rect 57428 2796 57480 2805
rect 57980 2796 58032 2848
rect 68468 2864 68520 2916
rect 74448 2932 74500 2984
rect 61752 2839 61804 2848
rect 61752 2805 61761 2839
rect 61761 2805 61795 2839
rect 61795 2805 61804 2839
rect 61752 2796 61804 2805
rect 62396 2839 62448 2848
rect 62396 2805 62405 2839
rect 62405 2805 62439 2839
rect 62439 2805 62448 2839
rect 62396 2796 62448 2805
rect 63224 2839 63276 2848
rect 63224 2805 63233 2839
rect 63233 2805 63267 2839
rect 63267 2805 63276 2839
rect 63224 2796 63276 2805
rect 63684 2839 63736 2848
rect 63684 2805 63693 2839
rect 63693 2805 63727 2839
rect 63727 2805 63736 2839
rect 63684 2796 63736 2805
rect 64328 2839 64380 2848
rect 64328 2805 64337 2839
rect 64337 2805 64371 2839
rect 64371 2805 64380 2839
rect 64328 2796 64380 2805
rect 65984 2839 66036 2848
rect 65984 2805 65993 2839
rect 65993 2805 66027 2839
rect 66027 2805 66036 2839
rect 65984 2796 66036 2805
rect 66444 2796 66496 2848
rect 67640 2796 67692 2848
rect 68652 2796 68704 2848
rect 72976 2796 73028 2848
rect 74264 2864 74316 2916
rect 76104 2796 76156 2848
rect 76748 2796 76800 2848
rect 78036 2839 78088 2848
rect 78036 2805 78045 2839
rect 78045 2805 78079 2839
rect 78079 2805 78088 2839
rect 78036 2796 78088 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 38660 2635 38712 2644
rect 38660 2601 38669 2635
rect 38669 2601 38703 2635
rect 38703 2601 38712 2635
rect 38660 2592 38712 2601
rect 40040 2592 40092 2644
rect 44180 2592 44232 2644
rect 43168 2524 43220 2576
rect 39488 2499 39540 2508
rect 39488 2465 39497 2499
rect 39497 2465 39531 2499
rect 39531 2465 39540 2499
rect 39488 2456 39540 2465
rect 32956 2431 33008 2440
rect 32956 2397 32965 2431
rect 32965 2397 32999 2431
rect 32999 2397 33008 2431
rect 32956 2388 33008 2397
rect 38016 2431 38068 2440
rect 38016 2397 38025 2431
rect 38025 2397 38059 2431
rect 38059 2397 38068 2431
rect 38016 2388 38068 2397
rect 38200 2431 38252 2440
rect 38200 2397 38209 2431
rect 38209 2397 38243 2431
rect 38243 2397 38252 2431
rect 38200 2388 38252 2397
rect 40684 2456 40736 2508
rect 41420 2388 41472 2440
rect 43536 2456 43588 2508
rect 43076 2431 43128 2440
rect 43076 2397 43085 2431
rect 43085 2397 43119 2431
rect 43119 2397 43128 2431
rect 43076 2388 43128 2397
rect 43260 2431 43312 2440
rect 43260 2397 43269 2431
rect 43269 2397 43303 2431
rect 43303 2397 43312 2431
rect 43260 2388 43312 2397
rect 43352 2431 43404 2440
rect 43352 2397 43361 2431
rect 43361 2397 43395 2431
rect 43395 2397 43404 2431
rect 43352 2388 43404 2397
rect 45560 2592 45612 2644
rect 50988 2592 51040 2644
rect 54668 2592 54720 2644
rect 57980 2592 58032 2644
rect 58716 2592 58768 2644
rect 59820 2592 59872 2644
rect 66536 2592 66588 2644
rect 67640 2592 67692 2644
rect 69756 2592 69808 2644
rect 71136 2592 71188 2644
rect 72240 2635 72292 2644
rect 72240 2601 72249 2635
rect 72249 2601 72283 2635
rect 72283 2601 72292 2635
rect 72240 2592 72292 2601
rect 45100 2456 45152 2508
rect 45008 2431 45060 2440
rect 45008 2397 45017 2431
rect 45017 2397 45051 2431
rect 45051 2397 45060 2431
rect 45008 2388 45060 2397
rect 45192 2388 45244 2440
rect 45836 2431 45888 2440
rect 45836 2397 45845 2431
rect 45845 2397 45879 2431
rect 45879 2397 45888 2431
rect 45836 2388 45888 2397
rect 46480 2431 46532 2440
rect 46480 2397 46489 2431
rect 46489 2397 46523 2431
rect 46523 2397 46532 2431
rect 46480 2388 46532 2397
rect 47124 2431 47176 2440
rect 47124 2397 47133 2431
rect 47133 2397 47167 2431
rect 47167 2397 47176 2431
rect 47124 2388 47176 2397
rect 47768 2431 47820 2440
rect 47768 2397 47777 2431
rect 47777 2397 47811 2431
rect 47811 2397 47820 2431
rect 47768 2388 47820 2397
rect 49700 2524 49752 2576
rect 54300 2524 54352 2576
rect 49056 2431 49108 2440
rect 49056 2397 49065 2431
rect 49065 2397 49099 2431
rect 49099 2397 49108 2431
rect 49056 2388 49108 2397
rect 49792 2388 49844 2440
rect 32864 2252 32916 2304
rect 42524 2252 42576 2304
rect 43812 2252 43864 2304
rect 50160 2363 50212 2372
rect 50160 2329 50169 2363
rect 50169 2329 50203 2363
rect 50203 2329 50212 2363
rect 50160 2320 50212 2329
rect 50252 2320 50304 2372
rect 51264 2431 51316 2440
rect 51264 2397 51273 2431
rect 51273 2397 51307 2431
rect 51307 2397 51316 2431
rect 51264 2388 51316 2397
rect 51632 2431 51684 2440
rect 51632 2397 51641 2431
rect 51641 2397 51675 2431
rect 51675 2397 51684 2431
rect 51632 2388 51684 2397
rect 53564 2431 53616 2440
rect 53564 2397 53573 2431
rect 53573 2397 53607 2431
rect 53607 2397 53616 2431
rect 53564 2388 53616 2397
rect 54484 2456 54536 2508
rect 55496 2524 55548 2576
rect 57336 2524 57388 2576
rect 59728 2524 59780 2576
rect 54116 2388 54168 2440
rect 56048 2456 56100 2508
rect 56692 2456 56744 2508
rect 57428 2456 57480 2508
rect 54852 2431 54904 2440
rect 54852 2397 54861 2431
rect 54861 2397 54895 2431
rect 54895 2397 54904 2431
rect 54852 2388 54904 2397
rect 55312 2431 55364 2440
rect 55312 2397 55321 2431
rect 55321 2397 55355 2431
rect 55355 2397 55364 2431
rect 55312 2388 55364 2397
rect 58164 2456 58216 2508
rect 59636 2456 59688 2508
rect 69020 2524 69072 2576
rect 71228 2524 71280 2576
rect 74080 2592 74132 2644
rect 74264 2592 74316 2644
rect 76104 2635 76156 2644
rect 76104 2601 76113 2635
rect 76113 2601 76147 2635
rect 76147 2601 76156 2635
rect 76104 2592 76156 2601
rect 77392 2635 77444 2644
rect 77392 2601 77401 2635
rect 77401 2601 77435 2635
rect 77435 2601 77444 2635
rect 77392 2592 77444 2601
rect 77760 2635 77812 2644
rect 77760 2601 77769 2635
rect 77769 2601 77803 2635
rect 77803 2601 77812 2635
rect 77760 2592 77812 2601
rect 45560 2295 45612 2304
rect 45560 2261 45569 2295
rect 45569 2261 45603 2295
rect 45603 2261 45612 2295
rect 45560 2252 45612 2261
rect 45744 2252 45796 2304
rect 46388 2295 46440 2304
rect 46388 2261 46397 2295
rect 46397 2261 46431 2295
rect 46431 2261 46440 2295
rect 46388 2252 46440 2261
rect 46480 2252 46532 2304
rect 47032 2252 47084 2304
rect 47676 2252 47728 2304
rect 48320 2252 48372 2304
rect 48964 2252 49016 2304
rect 49608 2252 49660 2304
rect 50896 2252 50948 2304
rect 51540 2252 51592 2304
rect 52184 2295 52236 2304
rect 52184 2261 52193 2295
rect 52193 2261 52227 2295
rect 52227 2261 52236 2295
rect 52184 2252 52236 2261
rect 52460 2295 52512 2304
rect 52460 2261 52469 2295
rect 52469 2261 52503 2295
rect 52503 2261 52512 2295
rect 52460 2252 52512 2261
rect 52828 2295 52880 2304
rect 52828 2261 52837 2295
rect 52837 2261 52871 2295
rect 52871 2261 52880 2295
rect 52828 2252 52880 2261
rect 53472 2252 53524 2304
rect 54760 2252 54812 2304
rect 55036 2295 55088 2304
rect 55036 2261 55045 2295
rect 55045 2261 55079 2295
rect 55079 2261 55088 2295
rect 55036 2252 55088 2261
rect 56600 2320 56652 2372
rect 57980 2388 58032 2440
rect 56968 2252 57020 2304
rect 58624 2320 58676 2372
rect 61752 2388 61804 2440
rect 62396 2388 62448 2440
rect 63224 2431 63276 2440
rect 63224 2397 63233 2431
rect 63233 2397 63267 2431
rect 63267 2397 63276 2431
rect 63224 2388 63276 2397
rect 63684 2388 63736 2440
rect 64328 2388 64380 2440
rect 68652 2431 68704 2440
rect 68652 2397 68661 2431
rect 68661 2397 68695 2431
rect 68695 2397 68704 2431
rect 68652 2388 68704 2397
rect 72056 2388 72108 2440
rect 57704 2295 57756 2304
rect 57704 2261 57713 2295
rect 57713 2261 57747 2295
rect 57747 2261 57756 2295
rect 57704 2252 57756 2261
rect 58348 2252 58400 2304
rect 59268 2295 59320 2304
rect 59268 2261 59277 2295
rect 59277 2261 59311 2295
rect 59311 2261 59320 2295
rect 59268 2252 59320 2261
rect 59360 2295 59412 2304
rect 59360 2261 59369 2295
rect 59369 2261 59403 2295
rect 59403 2261 59412 2295
rect 59360 2252 59412 2261
rect 59912 2295 59964 2304
rect 59912 2261 59921 2295
rect 59921 2261 59955 2295
rect 59955 2261 59964 2295
rect 59912 2252 59964 2261
rect 60556 2295 60608 2304
rect 60556 2261 60565 2295
rect 60565 2261 60599 2295
rect 60599 2261 60608 2295
rect 60556 2252 60608 2261
rect 61200 2295 61252 2304
rect 61200 2261 61209 2295
rect 61209 2261 61243 2295
rect 61243 2261 61252 2295
rect 61200 2252 61252 2261
rect 61844 2252 61896 2304
rect 62488 2252 62540 2304
rect 63132 2252 63184 2304
rect 63776 2252 63828 2304
rect 64420 2252 64472 2304
rect 65064 2295 65116 2304
rect 65064 2261 65073 2295
rect 65073 2261 65107 2295
rect 65107 2261 65116 2295
rect 65064 2252 65116 2261
rect 65340 2295 65392 2304
rect 65340 2261 65349 2295
rect 65349 2261 65383 2295
rect 65383 2261 65392 2295
rect 65340 2252 65392 2261
rect 65708 2295 65760 2304
rect 65708 2261 65717 2295
rect 65717 2261 65751 2295
rect 65751 2261 65760 2295
rect 65708 2252 65760 2261
rect 66076 2252 66128 2304
rect 66260 2295 66312 2304
rect 66260 2261 66269 2295
rect 66269 2261 66303 2295
rect 66303 2261 66312 2295
rect 66260 2252 66312 2261
rect 66996 2295 67048 2304
rect 66996 2261 67005 2295
rect 67005 2261 67039 2295
rect 67039 2261 67048 2295
rect 66996 2252 67048 2261
rect 67640 2295 67692 2304
rect 67640 2261 67649 2295
rect 67649 2261 67683 2295
rect 67683 2261 67692 2295
rect 67640 2252 67692 2261
rect 68284 2252 68336 2304
rect 68928 2295 68980 2304
rect 68928 2261 68937 2295
rect 68937 2261 68971 2295
rect 68971 2261 68980 2295
rect 68928 2252 68980 2261
rect 69572 2295 69624 2304
rect 69572 2261 69581 2295
rect 69581 2261 69615 2295
rect 69615 2261 69624 2295
rect 69572 2252 69624 2261
rect 70216 2295 70268 2304
rect 70216 2261 70225 2295
rect 70225 2261 70259 2295
rect 70259 2261 70268 2295
rect 70216 2252 70268 2261
rect 70860 2295 70912 2304
rect 70860 2261 70869 2295
rect 70869 2261 70903 2295
rect 70903 2261 70912 2295
rect 70860 2252 70912 2261
rect 71136 2295 71188 2304
rect 71136 2261 71145 2295
rect 71145 2261 71179 2295
rect 71179 2261 71188 2295
rect 71136 2252 71188 2261
rect 71504 2295 71556 2304
rect 71504 2261 71513 2295
rect 71513 2261 71547 2295
rect 71547 2261 71556 2295
rect 71504 2252 71556 2261
rect 72884 2431 72936 2440
rect 72884 2397 72893 2431
rect 72893 2397 72927 2431
rect 72927 2397 72936 2431
rect 72884 2388 72936 2397
rect 72240 2320 72292 2372
rect 73436 2320 73488 2372
rect 76748 2431 76800 2440
rect 76748 2397 76757 2431
rect 76757 2397 76791 2431
rect 76791 2397 76800 2431
rect 76748 2388 76800 2397
rect 77944 2431 77996 2440
rect 77944 2397 77953 2431
rect 77953 2397 77987 2431
rect 77987 2397 77996 2431
rect 77944 2388 77996 2397
rect 78036 2431 78088 2440
rect 78036 2397 78045 2431
rect 78045 2397 78079 2431
rect 78079 2397 78088 2431
rect 78036 2388 78088 2397
rect 72792 2252 72844 2304
rect 74080 2295 74132 2304
rect 74080 2261 74089 2295
rect 74089 2261 74123 2295
rect 74123 2261 74132 2295
rect 74080 2252 74132 2261
rect 74724 2295 74776 2304
rect 74724 2261 74733 2295
rect 74733 2261 74767 2295
rect 74767 2261 74776 2295
rect 74724 2252 74776 2261
rect 75368 2295 75420 2304
rect 75368 2261 75377 2295
rect 75377 2261 75411 2295
rect 75411 2261 75420 2295
rect 75368 2252 75420 2261
rect 76012 2295 76064 2304
rect 76012 2261 76021 2295
rect 76021 2261 76055 2295
rect 76055 2261 76064 2295
rect 76012 2252 76064 2261
rect 76656 2252 76708 2304
rect 77300 2295 77352 2304
rect 77300 2261 77309 2295
rect 77309 2261 77343 2295
rect 77343 2261 77352 2295
rect 77300 2252 77352 2261
rect 78588 2252 78640 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 66314 2150 66366 2202
rect 66378 2150 66430 2202
rect 66442 2150 66494 2202
rect 66506 2150 66558 2202
rect 66570 2150 66622 2202
rect 44456 2048 44508 2100
rect 45192 2048 45244 2100
rect 45560 2048 45612 2100
rect 54852 2048 54904 2100
rect 55036 2048 55088 2100
rect 60004 2048 60056 2100
rect 65340 2048 65392 2100
rect 43352 1980 43404 2032
rect 46388 1980 46440 2032
rect 65984 1980 66036 2032
rect 72424 1980 72476 2032
rect 50160 1912 50212 1964
rect 54484 1912 54536 1964
rect 59360 1912 59412 1964
rect 66076 1912 66128 1964
rect 72516 1912 72568 1964
rect 52460 1844 52512 1896
rect 58808 1844 58860 1896
rect 50160 1776 50212 1828
rect 55220 1776 55272 1828
<< metal2 >>
rect 38658 39200 38714 40000
rect 39302 39200 39358 40000
rect 39946 39200 40002 40000
rect 40590 39200 40646 40000
rect 41234 39200 41290 40000
rect 41878 39200 41934 40000
rect 42522 39200 42578 40000
rect 43166 39200 43222 40000
rect 43810 39200 43866 40000
rect 44454 39200 44510 40000
rect 45098 39200 45154 40000
rect 45742 39200 45798 40000
rect 46386 39200 46442 40000
rect 47030 39200 47086 40000
rect 47674 39200 47730 40000
rect 48318 39200 48374 40000
rect 48962 39200 49018 40000
rect 49606 39200 49662 40000
rect 50250 39200 50306 40000
rect 50894 39200 50950 40000
rect 51538 39200 51594 40000
rect 52182 39200 52238 40000
rect 52826 39200 52882 40000
rect 53470 39200 53526 40000
rect 54114 39200 54170 40000
rect 54758 39200 54814 40000
rect 55402 39200 55458 40000
rect 56046 39200 56102 40000
rect 56690 39200 56746 40000
rect 57334 39200 57390 40000
rect 57978 39200 58034 40000
rect 58622 39200 58678 40000
rect 59266 39200 59322 40000
rect 59910 39200 59966 40000
rect 60554 39200 60610 40000
rect 61198 39200 61254 40000
rect 61842 39200 61898 40000
rect 62486 39200 62542 40000
rect 63130 39200 63186 40000
rect 63774 39200 63830 40000
rect 64418 39200 64474 40000
rect 65062 39200 65118 40000
rect 65706 39200 65762 40000
rect 66350 39200 66406 40000
rect 66994 39200 67050 40000
rect 67638 39200 67694 40000
rect 68282 39200 68338 40000
rect 68926 39200 68982 40000
rect 69570 39200 69626 40000
rect 70214 39200 70270 40000
rect 70858 39200 70914 40000
rect 71502 39200 71558 40000
rect 72146 39200 72202 40000
rect 72790 39200 72846 40000
rect 73434 39200 73490 40000
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 38672 37466 38700 39200
rect 38660 37460 38712 37466
rect 38660 37402 38712 37408
rect 36268 37256 36320 37262
rect 36268 37198 36320 37204
rect 35440 37120 35492 37126
rect 35440 37062 35492 37068
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 1306 36816 1362 36825
rect 35452 36786 35480 37062
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 36280 36922 36308 37198
rect 36268 36916 36320 36922
rect 36268 36858 36320 36864
rect 1306 36751 1362 36760
rect 35440 36780 35492 36786
rect 1320 36378 1348 36751
rect 35440 36722 35492 36728
rect 2136 36712 2188 36718
rect 2136 36654 2188 36660
rect 32220 36712 32272 36718
rect 32220 36654 32272 36660
rect 33232 36712 33284 36718
rect 33232 36654 33284 36660
rect 33876 36712 33928 36718
rect 33876 36654 33928 36660
rect 34152 36712 34204 36718
rect 34152 36654 34204 36660
rect 36176 36712 36228 36718
rect 36176 36654 36228 36660
rect 1308 36372 1360 36378
rect 1308 36314 1360 36320
rect 2148 36174 2176 36654
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 32232 36378 32260 36654
rect 32220 36372 32272 36378
rect 32220 36314 32272 36320
rect 2136 36168 2188 36174
rect 938 36136 994 36145
rect 2136 36110 2188 36116
rect 938 36071 994 36080
rect 952 36038 980 36071
rect 940 36032 992 36038
rect 940 35974 992 35980
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 940 35488 992 35494
rect 938 35456 940 35465
rect 31484 35488 31536 35494
rect 992 35456 994 35465
rect 31484 35430 31536 35436
rect 938 35391 994 35400
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 31496 35154 31524 35430
rect 28632 35148 28684 35154
rect 28632 35090 28684 35096
rect 28724 35148 28776 35154
rect 28724 35090 28776 35096
rect 31484 35148 31536 35154
rect 31484 35090 31536 35096
rect 2044 34944 2096 34950
rect 2044 34886 2096 34892
rect 1306 34776 1362 34785
rect 1306 34711 1308 34720
rect 1360 34711 1362 34720
rect 1308 34682 1360 34688
rect 2056 34610 2084 34886
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 2044 34604 2096 34610
rect 2044 34546 2096 34552
rect 2136 34536 2188 34542
rect 2136 34478 2188 34484
rect 940 34128 992 34134
rect 938 34096 940 34105
rect 992 34096 994 34105
rect 938 34031 994 34040
rect 2148 33998 2176 34478
rect 28356 34468 28408 34474
rect 28356 34410 28408 34416
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 28368 33998 28396 34410
rect 28448 34128 28500 34134
rect 28448 34070 28500 34076
rect 2136 33992 2188 33998
rect 2136 33934 2188 33940
rect 26976 33992 27028 33998
rect 26976 33934 27028 33940
rect 28356 33992 28408 33998
rect 28356 33934 28408 33940
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 938 33416 994 33425
rect 938 33351 940 33360
rect 992 33351 994 33360
rect 940 33322 992 33328
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 940 32768 992 32774
rect 938 32736 940 32745
rect 992 32736 994 32745
rect 938 32671 994 32680
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 17684 32496 17736 32502
rect 17684 32438 17736 32444
rect 18696 32496 18748 32502
rect 18696 32438 18748 32444
rect 2044 32360 2096 32366
rect 2044 32302 2096 32308
rect 17408 32360 17460 32366
rect 17408 32302 17460 32308
rect 1306 32056 1362 32065
rect 1306 31991 1308 32000
rect 1360 31991 1362 32000
rect 1308 31962 1360 31968
rect 2056 31822 2084 32302
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 17420 32026 17448 32302
rect 17408 32020 17460 32026
rect 17408 31962 17460 31968
rect 17696 31890 17724 32438
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 17684 31884 17736 31890
rect 17684 31826 17736 31832
rect 2044 31816 2096 31822
rect 2044 31758 2096 31764
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 15384 31816 15436 31822
rect 15384 31758 15436 31764
rect 2044 31680 2096 31686
rect 2044 31622 2096 31628
rect 940 31476 992 31482
rect 940 31418 992 31424
rect 952 31385 980 31418
rect 938 31376 994 31385
rect 2056 31346 2084 31622
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 11348 31362 11376 31758
rect 12348 31748 12400 31754
rect 12348 31690 12400 31696
rect 13636 31748 13688 31754
rect 13636 31690 13688 31696
rect 14740 31748 14792 31754
rect 14740 31690 14792 31696
rect 11612 31408 11664 31414
rect 11348 31346 11468 31362
rect 11612 31350 11664 31356
rect 938 31311 994 31320
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 11348 31340 11480 31346
rect 11348 31334 11428 31340
rect 9864 31272 9916 31278
rect 9864 31214 9916 31220
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 938 30696 994 30705
rect 938 30631 994 30640
rect 952 30598 980 30631
rect 940 30592 992 30598
rect 940 30534 992 30540
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 940 30048 992 30054
rect 938 30016 940 30025
rect 992 30016 994 30025
rect 938 29951 994 29960
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 9692 29714 9720 31078
rect 9876 30938 9904 31214
rect 11348 31142 11376 31334
rect 11428 31282 11480 31288
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 11428 31136 11480 31142
rect 11428 31078 11480 31084
rect 9864 30932 9916 30938
rect 9864 30874 9916 30880
rect 11440 30734 11468 31078
rect 11244 30728 11296 30734
rect 11244 30670 11296 30676
rect 11428 30728 11480 30734
rect 11428 30670 11480 30676
rect 11256 30394 11284 30670
rect 11244 30388 11296 30394
rect 11244 30330 11296 30336
rect 9680 29708 9732 29714
rect 9680 29650 9732 29656
rect 10232 29708 10284 29714
rect 10232 29650 10284 29656
rect 11152 29708 11204 29714
rect 11152 29650 11204 29656
rect 9220 29572 9272 29578
rect 9220 29514 9272 29520
rect 2044 29504 2096 29510
rect 2044 29446 2096 29452
rect 1306 29336 1362 29345
rect 1306 29271 1308 29280
rect 1360 29271 1362 29280
rect 1308 29242 1360 29248
rect 2056 29170 2084 29446
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 2044 29164 2096 29170
rect 2044 29106 2096 29112
rect 9232 29102 9260 29514
rect 2136 29096 2188 29102
rect 2136 29038 2188 29044
rect 9220 29096 9272 29102
rect 9220 29038 9272 29044
rect 940 28688 992 28694
rect 938 28656 940 28665
rect 992 28656 994 28665
rect 938 28591 994 28600
rect 2148 28558 2176 29038
rect 10244 29034 10272 29650
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10796 29170 10824 29446
rect 11164 29306 11192 29650
rect 11152 29300 11204 29306
rect 11152 29242 11204 29248
rect 10784 29164 10836 29170
rect 10784 29106 10836 29112
rect 10876 29164 10928 29170
rect 10876 29106 10928 29112
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 2136 28552 2188 28558
rect 2136 28494 2188 28500
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 9508 28218 9536 28494
rect 9496 28212 9548 28218
rect 9496 28154 9548 28160
rect 10244 28014 10272 28970
rect 10888 28778 10916 29106
rect 10796 28762 11008 28778
rect 10784 28756 11008 28762
rect 10836 28750 11008 28756
rect 10784 28698 10836 28704
rect 10876 28484 10928 28490
rect 10876 28426 10928 28432
rect 10508 28416 10560 28422
rect 10508 28358 10560 28364
rect 10520 28082 10548 28358
rect 10692 28212 10744 28218
rect 10692 28154 10744 28160
rect 10508 28076 10560 28082
rect 10508 28018 10560 28024
rect 10600 28076 10652 28082
rect 10600 28018 10652 28024
rect 10232 28008 10284 28014
rect 938 27976 994 27985
rect 10232 27950 10284 27956
rect 938 27911 940 27920
rect 992 27911 994 27920
rect 940 27882 992 27888
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 940 27328 992 27334
rect 938 27296 940 27305
rect 992 27296 994 27305
rect 938 27231 994 27240
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 10048 27056 10100 27062
rect 10048 26998 10100 27004
rect 2044 26920 2096 26926
rect 2044 26862 2096 26868
rect 1306 26616 1362 26625
rect 1306 26551 1308 26560
rect 1360 26551 1362 26560
rect 1308 26522 1360 26528
rect 2056 26382 2084 26862
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 2044 26376 2096 26382
rect 2044 26318 2096 26324
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 10060 26042 10088 26998
rect 10140 26784 10192 26790
rect 10140 26726 10192 26732
rect 10152 26314 10180 26726
rect 10244 26450 10272 27950
rect 10612 27674 10640 28018
rect 10600 27668 10652 27674
rect 10600 27610 10652 27616
rect 10612 26994 10640 27610
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 10704 26450 10732 28154
rect 10784 28076 10836 28082
rect 10784 28018 10836 28024
rect 10796 27130 10824 28018
rect 10888 27962 10916 28426
rect 10980 28082 11008 28750
rect 11164 28694 11192 29242
rect 11256 29170 11284 30330
rect 11624 29850 11652 31350
rect 11888 31272 11940 31278
rect 11888 31214 11940 31220
rect 12256 31272 12308 31278
rect 12256 31214 12308 31220
rect 11704 30796 11756 30802
rect 11704 30738 11756 30744
rect 11716 30666 11744 30738
rect 11704 30660 11756 30666
rect 11704 30602 11756 30608
rect 11716 30122 11744 30602
rect 11900 30258 11928 31214
rect 11888 30252 11940 30258
rect 11888 30194 11940 30200
rect 11704 30116 11756 30122
rect 11704 30058 11756 30064
rect 11612 29844 11664 29850
rect 11612 29786 11664 29792
rect 11624 29578 11652 29786
rect 11612 29572 11664 29578
rect 11612 29514 11664 29520
rect 11900 29170 11928 30194
rect 12268 30122 12296 31214
rect 12360 30938 12388 31690
rect 13648 31482 13676 31690
rect 13820 31680 13872 31686
rect 13820 31622 13872 31628
rect 13636 31476 13688 31482
rect 13636 31418 13688 31424
rect 13832 31278 13860 31622
rect 13820 31272 13872 31278
rect 13820 31214 13872 31220
rect 12808 31136 12860 31142
rect 12808 31078 12860 31084
rect 13544 31136 13596 31142
rect 13544 31078 13596 31084
rect 12348 30932 12400 30938
rect 12348 30874 12400 30880
rect 12820 30734 12848 31078
rect 12808 30728 12860 30734
rect 12808 30670 12860 30676
rect 13556 30394 13584 31078
rect 13544 30388 13596 30394
rect 13544 30330 13596 30336
rect 12532 30252 12584 30258
rect 13544 30252 13596 30258
rect 12532 30194 12584 30200
rect 13096 30212 13544 30240
rect 12544 30161 12572 30194
rect 12530 30152 12586 30161
rect 12256 30116 12308 30122
rect 13096 30122 13124 30212
rect 13544 30194 13596 30200
rect 14556 30184 14608 30190
rect 14554 30152 14556 30161
rect 14608 30152 14610 30161
rect 12530 30087 12586 30096
rect 13084 30116 13136 30122
rect 12256 30058 12308 30064
rect 13360 30116 13412 30122
rect 13084 30058 13136 30064
rect 13280 30076 13360 30104
rect 11244 29164 11296 29170
rect 11244 29106 11296 29112
rect 11336 29164 11388 29170
rect 11336 29106 11388 29112
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 11256 28762 11284 29106
rect 11244 28756 11296 28762
rect 11244 28698 11296 28704
rect 11152 28688 11204 28694
rect 11152 28630 11204 28636
rect 11348 28490 11376 29106
rect 12268 28966 12296 30058
rect 13280 29238 13308 30076
rect 14610 30110 14688 30138
rect 14554 30087 14610 30096
rect 13360 30058 13412 30064
rect 14660 29646 14688 30110
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 14556 29504 14608 29510
rect 14556 29446 14608 29452
rect 13360 29300 13412 29306
rect 13360 29242 13412 29248
rect 13268 29232 13320 29238
rect 13268 29174 13320 29180
rect 13268 29096 13320 29102
rect 13268 29038 13320 29044
rect 12256 28960 12308 28966
rect 12256 28902 12308 28908
rect 13280 28626 13308 29038
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 13268 28620 13320 28626
rect 13268 28562 13320 28568
rect 11336 28484 11388 28490
rect 11336 28426 11388 28432
rect 11440 28422 11468 28562
rect 11428 28416 11480 28422
rect 11428 28358 11480 28364
rect 10968 28076 11020 28082
rect 10968 28018 11020 28024
rect 10888 27934 11008 27962
rect 10980 27470 11008 27934
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 11336 27464 11388 27470
rect 11440 27418 11468 28358
rect 13280 28150 13308 28562
rect 13372 28558 13400 29242
rect 14568 28762 14596 29446
rect 14660 29102 14688 29582
rect 14752 29306 14780 31690
rect 15292 31680 15344 31686
rect 15292 31622 15344 31628
rect 15304 31414 15332 31622
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15396 30938 15424 31758
rect 16304 31748 16356 31754
rect 16304 31690 16356 31696
rect 17132 31748 17184 31754
rect 17132 31690 17184 31696
rect 16316 31414 16344 31690
rect 16304 31408 16356 31414
rect 16304 31350 16356 31356
rect 16488 31136 16540 31142
rect 16488 31078 16540 31084
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 15384 30932 15436 30938
rect 15384 30874 15436 30880
rect 15200 30728 15252 30734
rect 15200 30670 15252 30676
rect 15212 30394 15240 30670
rect 15292 30592 15344 30598
rect 15292 30534 15344 30540
rect 15200 30388 15252 30394
rect 15200 30330 15252 30336
rect 15212 30258 15240 30330
rect 15200 30252 15252 30258
rect 15200 30194 15252 30200
rect 14740 29300 14792 29306
rect 14740 29242 14792 29248
rect 15212 29170 15240 30194
rect 15304 30054 15332 30534
rect 15476 30320 15528 30326
rect 15476 30262 15528 30268
rect 15292 30048 15344 30054
rect 15292 29990 15344 29996
rect 15488 29850 15516 30262
rect 16500 30258 16528 31078
rect 16684 30734 16712 31078
rect 17144 30734 17172 31690
rect 17696 31346 17724 31826
rect 18524 31822 18552 32166
rect 18512 31816 18564 31822
rect 18512 31758 18564 31764
rect 18708 31482 18736 32438
rect 26988 31890 27016 33934
rect 27252 33924 27304 33930
rect 27252 33866 27304 33872
rect 27264 33658 27292 33866
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27988 32768 28040 32774
rect 27988 32710 28040 32716
rect 27344 32564 27396 32570
rect 27344 32506 27396 32512
rect 27252 32360 27304 32366
rect 27252 32302 27304 32308
rect 27264 32026 27292 32302
rect 27252 32020 27304 32026
rect 27252 31962 27304 31968
rect 21456 31884 21508 31890
rect 21456 31826 21508 31832
rect 26976 31884 27028 31890
rect 26976 31826 27028 31832
rect 18788 31816 18840 31822
rect 18788 31758 18840 31764
rect 18696 31476 18748 31482
rect 18616 31436 18696 31464
rect 17684 31340 17736 31346
rect 17684 31282 17736 31288
rect 18512 31272 18564 31278
rect 18512 31214 18564 31220
rect 18524 30938 18552 31214
rect 18512 30932 18564 30938
rect 18512 30874 18564 30880
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 17132 30728 17184 30734
rect 17132 30670 17184 30676
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 16488 30252 16540 30258
rect 16488 30194 16540 30200
rect 17144 30122 17172 30670
rect 17960 30592 18012 30598
rect 17960 30534 18012 30540
rect 17972 30394 18000 30534
rect 17960 30388 18012 30394
rect 17960 30330 18012 30336
rect 18432 30258 18460 30670
rect 17408 30252 17460 30258
rect 17408 30194 17460 30200
rect 18420 30252 18472 30258
rect 18420 30194 18472 30200
rect 17132 30116 17184 30122
rect 17132 30058 17184 30064
rect 15844 30048 15896 30054
rect 15844 29990 15896 29996
rect 15856 29850 15884 29990
rect 15476 29844 15528 29850
rect 15476 29786 15528 29792
rect 15844 29844 15896 29850
rect 15844 29786 15896 29792
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 15856 29646 15884 29786
rect 15844 29640 15896 29646
rect 15844 29582 15896 29588
rect 15856 29170 15884 29582
rect 16304 29572 16356 29578
rect 16304 29514 16356 29520
rect 15200 29164 15252 29170
rect 15200 29106 15252 29112
rect 15844 29164 15896 29170
rect 15844 29106 15896 29112
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 14556 28756 14608 28762
rect 14556 28698 14608 28704
rect 15212 28626 15240 29106
rect 16316 29034 16344 29514
rect 16500 29102 16528 29786
rect 17420 29714 17448 30194
rect 17684 30048 17736 30054
rect 17684 29990 17736 29996
rect 17408 29708 17460 29714
rect 17408 29650 17460 29656
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16488 29096 16540 29102
rect 16488 29038 16540 29044
rect 15292 29028 15344 29034
rect 15292 28970 15344 28976
rect 16304 29028 16356 29034
rect 16304 28970 16356 28976
rect 15200 28620 15252 28626
rect 15200 28562 15252 28568
rect 15304 28558 15332 28970
rect 15660 28960 15712 28966
rect 15660 28902 15712 28908
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 13360 28552 13412 28558
rect 13360 28494 13412 28500
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 13268 28144 13320 28150
rect 13268 28086 13320 28092
rect 13360 28008 13412 28014
rect 13360 27950 13412 27956
rect 13372 27606 13400 27950
rect 14660 27878 14688 28494
rect 15476 28484 15528 28490
rect 15476 28426 15528 28432
rect 15108 28416 15160 28422
rect 15108 28358 15160 28364
rect 14740 28212 14792 28218
rect 14740 28154 14792 28160
rect 14752 28014 14780 28154
rect 15016 28144 15068 28150
rect 15016 28086 15068 28092
rect 14740 28008 14792 28014
rect 14740 27950 14792 27956
rect 14648 27872 14700 27878
rect 14648 27814 14700 27820
rect 13360 27600 13412 27606
rect 13360 27542 13412 27548
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 11388 27412 11468 27418
rect 11336 27406 11468 27412
rect 10784 27124 10836 27130
rect 10784 27066 10836 27072
rect 10980 26586 11008 27406
rect 11348 27390 11468 27406
rect 11348 26994 11376 27390
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 12084 26994 12112 27066
rect 12452 26994 12480 27474
rect 14660 27470 14688 27814
rect 14752 27538 14780 27950
rect 14740 27532 14792 27538
rect 14740 27474 14792 27480
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 11336 26988 11388 26994
rect 11336 26930 11388 26936
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 13360 26988 13412 26994
rect 13360 26930 13412 26936
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 10232 26444 10284 26450
rect 10232 26386 10284 26392
rect 10692 26444 10744 26450
rect 10692 26386 10744 26392
rect 10704 26314 10732 26386
rect 10140 26308 10192 26314
rect 10140 26250 10192 26256
rect 10324 26308 10376 26314
rect 10324 26250 10376 26256
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 940 26036 992 26042
rect 940 25978 992 25984
rect 10048 26036 10100 26042
rect 10048 25978 10100 25984
rect 952 25945 980 25978
rect 938 25936 994 25945
rect 938 25871 994 25880
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 938 25256 994 25265
rect 938 25191 994 25200
rect 952 25158 980 25191
rect 940 25152 992 25158
rect 940 25094 992 25100
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 7748 24744 7800 24750
rect 7748 24686 7800 24692
rect 9036 24744 9088 24750
rect 9036 24686 9088 24692
rect 940 24608 992 24614
rect 938 24576 940 24585
rect 992 24576 994 24585
rect 938 24511 994 24520
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 2044 24064 2096 24070
rect 2044 24006 2096 24012
rect 1306 23896 1362 23905
rect 1306 23831 1308 23840
rect 1360 23831 1362 23840
rect 1308 23802 1360 23808
rect 2056 23730 2084 24006
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 7760 23730 7788 24686
rect 9048 24410 9076 24686
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9036 24404 9088 24410
rect 9036 24346 9088 24352
rect 9600 24206 9628 24550
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 10060 24138 10088 25978
rect 10048 24132 10100 24138
rect 10048 24074 10100 24080
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 9048 23798 9076 24006
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9036 23792 9088 23798
rect 9036 23734 9088 23740
rect 2044 23724 2096 23730
rect 2044 23666 2096 23672
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 2136 23656 2188 23662
rect 2136 23598 2188 23604
rect 1216 23248 1268 23254
rect 1214 23216 1216 23225
rect 1268 23216 1270 23225
rect 1214 23151 1270 23160
rect 2148 23118 2176 23598
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 2136 23112 2188 23118
rect 2136 23054 2188 23060
rect 940 22976 992 22982
rect 940 22918 992 22924
rect 952 22681 980 22918
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 938 22672 994 22681
rect 938 22607 994 22616
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 7012 22024 7064 22030
rect 846 21992 902 22001
rect 7012 21966 7064 21972
rect 846 21927 902 21936
rect 860 21894 888 21927
rect 848 21888 900 21894
rect 848 21830 900 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 848 21344 900 21350
rect 846 21312 848 21321
rect 900 21312 902 21321
rect 846 21247 902 21256
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 7024 21010 7052 21966
rect 7760 21622 7788 23666
rect 9692 22710 9720 23802
rect 10336 23798 10364 26250
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 10416 24676 10468 24682
rect 10416 24618 10468 24624
rect 10428 24138 10456 24618
rect 10888 24206 10916 24754
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 11152 24744 11204 24750
rect 11152 24686 11204 24692
rect 11072 24274 11100 24686
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 10416 24132 10468 24138
rect 10416 24074 10468 24080
rect 10612 23798 10640 24142
rect 10324 23792 10376 23798
rect 10324 23734 10376 23740
rect 10600 23792 10652 23798
rect 10600 23734 10652 23740
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9692 22098 9720 22646
rect 9680 22092 9732 22098
rect 10336 22094 10364 23734
rect 10888 23730 10916 24142
rect 10980 23866 11008 24142
rect 10968 23860 11020 23866
rect 10968 23802 11020 23808
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 11072 23594 11100 24210
rect 11164 24138 11192 24686
rect 11244 24676 11296 24682
rect 11244 24618 11296 24624
rect 11256 24138 11284 24618
rect 11348 24342 11376 26930
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11992 26586 12020 26726
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 12084 26382 12112 26930
rect 12164 26852 12216 26858
rect 12164 26794 12216 26800
rect 12072 26376 12124 26382
rect 12072 26318 12124 26324
rect 12176 26314 12204 26794
rect 12452 26586 12480 26930
rect 12532 26852 12584 26858
rect 12532 26794 12584 26800
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12544 26450 12572 26794
rect 13004 26790 13032 26930
rect 12992 26784 13044 26790
rect 12992 26726 13044 26732
rect 12532 26444 12584 26450
rect 12532 26386 12584 26392
rect 12900 26444 12952 26450
rect 12900 26386 12952 26392
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 12452 25362 12480 26318
rect 12440 25356 12492 25362
rect 12440 25298 12492 25304
rect 12912 25294 12940 26386
rect 13004 26382 13032 26726
rect 13372 26518 13400 26930
rect 14660 26790 14688 27406
rect 14752 26994 14780 27474
rect 15028 27402 15056 28086
rect 15016 27396 15068 27402
rect 15016 27338 15068 27344
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14648 26784 14700 26790
rect 14648 26726 14700 26732
rect 13360 26512 13412 26518
rect 13360 26454 13412 26460
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 12992 26036 13044 26042
rect 12992 25978 13044 25984
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 12900 24948 12952 24954
rect 12900 24890 12952 24896
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 11336 24336 11388 24342
rect 11336 24278 11388 24284
rect 11900 24274 11928 24550
rect 12544 24274 12572 24754
rect 11888 24268 11940 24274
rect 11888 24210 11940 24216
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 11152 24132 11204 24138
rect 11152 24074 11204 24080
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 11164 23730 11192 24074
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 10876 23520 10928 23526
rect 10876 23462 10928 23468
rect 10888 23186 10916 23462
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10704 22778 10732 23054
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 11072 22574 11100 23530
rect 11152 23180 11204 23186
rect 11152 23122 11204 23128
rect 11060 22568 11112 22574
rect 11060 22510 11112 22516
rect 9680 22034 9732 22040
rect 10060 22066 10364 22094
rect 10060 21962 10088 22066
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 10060 21622 10088 21898
rect 11072 21894 11100 22510
rect 11164 22234 11192 23122
rect 12912 22574 12940 24890
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 12452 22098 12480 22510
rect 13004 22166 13032 25978
rect 14556 25696 14608 25702
rect 14556 25638 14608 25644
rect 14568 25498 14596 25638
rect 13820 25492 13872 25498
rect 13820 25434 13872 25440
rect 14556 25492 14608 25498
rect 14556 25434 14608 25440
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 13188 24682 13216 25162
rect 13464 24750 13492 25230
rect 13740 24954 13768 25230
rect 13728 24948 13780 24954
rect 13728 24890 13780 24896
rect 13740 24818 13768 24890
rect 13832 24886 13860 25434
rect 15028 25378 15056 27338
rect 15120 25974 15148 28358
rect 15488 28082 15516 28426
rect 15672 28082 15700 28902
rect 15752 28552 15804 28558
rect 15752 28494 15804 28500
rect 15764 28082 15792 28494
rect 15948 28490 15976 28902
rect 16316 28490 16344 28970
rect 16500 28490 16528 29038
rect 16684 28626 16712 29106
rect 16672 28620 16724 28626
rect 16672 28562 16724 28568
rect 17420 28558 17448 29650
rect 17696 29578 17724 29990
rect 18432 29850 18460 30194
rect 17776 29844 17828 29850
rect 18420 29844 18472 29850
rect 17828 29804 17908 29832
rect 17776 29786 17828 29792
rect 17880 29730 17908 29804
rect 18420 29786 18472 29792
rect 17880 29702 18092 29730
rect 17684 29572 17736 29578
rect 17684 29514 17736 29520
rect 17960 29572 18012 29578
rect 17960 29514 18012 29520
rect 17408 28552 17460 28558
rect 17408 28494 17460 28500
rect 17592 28552 17644 28558
rect 17592 28494 17644 28500
rect 15936 28484 15988 28490
rect 15936 28426 15988 28432
rect 16304 28484 16356 28490
rect 16304 28426 16356 28432
rect 16488 28484 16540 28490
rect 16488 28426 16540 28432
rect 16028 28416 16080 28422
rect 16028 28358 16080 28364
rect 16120 28416 16172 28422
rect 16120 28358 16172 28364
rect 16040 28150 16068 28358
rect 16028 28144 16080 28150
rect 16028 28086 16080 28092
rect 16132 28082 16160 28358
rect 15476 28076 15528 28082
rect 15476 28018 15528 28024
rect 15660 28076 15712 28082
rect 15660 28018 15712 28024
rect 15752 28076 15804 28082
rect 15752 28018 15804 28024
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 15488 26042 15516 28018
rect 16120 27872 16172 27878
rect 16120 27814 16172 27820
rect 16132 27674 16160 27814
rect 17604 27674 17632 28494
rect 17972 28218 18000 29514
rect 18064 29510 18092 29702
rect 18052 29504 18104 29510
rect 18052 29446 18104 29452
rect 17960 28212 18012 28218
rect 17960 28154 18012 28160
rect 18616 28150 18644 31436
rect 18696 31418 18748 31424
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18708 30326 18736 31214
rect 18800 30394 18828 31758
rect 20168 31748 20220 31754
rect 20168 31690 20220 31696
rect 19524 31136 19576 31142
rect 19524 31078 19576 31084
rect 19536 30802 19564 31078
rect 19524 30796 19576 30802
rect 19524 30738 19576 30744
rect 18788 30388 18840 30394
rect 18788 30330 18840 30336
rect 18696 30320 18748 30326
rect 18696 30262 18748 30268
rect 18708 29646 18736 30262
rect 18800 29850 18828 30330
rect 19064 30184 19116 30190
rect 19064 30126 19116 30132
rect 18788 29844 18840 29850
rect 18788 29786 18840 29792
rect 19076 29646 19104 30126
rect 19248 30048 19300 30054
rect 19248 29990 19300 29996
rect 19260 29646 19288 29990
rect 19984 29708 20036 29714
rect 19984 29650 20036 29656
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 19064 29640 19116 29646
rect 19064 29582 19116 29588
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19076 29306 19104 29582
rect 19064 29300 19116 29306
rect 19064 29242 19116 29248
rect 19340 29164 19392 29170
rect 19168 29124 19340 29152
rect 18604 28144 18656 28150
rect 18604 28086 18656 28092
rect 18616 27878 18644 28086
rect 18604 27872 18656 27878
rect 18604 27814 18656 27820
rect 16120 27668 16172 27674
rect 16120 27610 16172 27616
rect 17592 27668 17644 27674
rect 17592 27610 17644 27616
rect 17960 27328 18012 27334
rect 17960 27270 18012 27276
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 17972 26058 18000 27270
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 18156 26790 18184 27066
rect 18524 27062 18552 27270
rect 18616 27130 18644 27814
rect 18604 27124 18656 27130
rect 18604 27066 18656 27072
rect 18512 27056 18564 27062
rect 18512 26998 18564 27004
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 18144 26784 18196 26790
rect 18144 26726 18196 26732
rect 17972 26042 18092 26058
rect 15476 26036 15528 26042
rect 15476 25978 15528 25984
rect 16948 26036 17000 26042
rect 16948 25978 17000 25984
rect 17960 26036 18092 26042
rect 18012 26030 18092 26036
rect 17960 25978 18012 25984
rect 15108 25968 15160 25974
rect 15108 25910 15160 25916
rect 14936 25350 15056 25378
rect 16580 25356 16632 25362
rect 14372 25288 14424 25294
rect 14372 25230 14424 25236
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14384 24954 14412 25230
rect 14372 24948 14424 24954
rect 14372 24890 14424 24896
rect 13820 24880 13872 24886
rect 13820 24822 13872 24828
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 13452 24744 13504 24750
rect 13452 24686 13504 24692
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 13464 24410 13492 24686
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13648 24206 13676 24550
rect 13820 24404 13872 24410
rect 13820 24346 13872 24352
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13832 24070 13860 24346
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 14292 23866 14320 24754
rect 14384 24682 14412 24890
rect 14476 24682 14504 25230
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 14384 24562 14412 24618
rect 14384 24534 14504 24562
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 13728 23044 13780 23050
rect 13728 22986 13780 22992
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 13096 22642 13124 22918
rect 13740 22710 13768 22986
rect 13728 22704 13780 22710
rect 13728 22646 13780 22652
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 14096 22500 14148 22506
rect 14096 22442 14148 22448
rect 12992 22160 13044 22166
rect 12992 22102 13044 22108
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 12452 21690 12480 22034
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 7748 21616 7800 21622
rect 9680 21616 9732 21622
rect 7800 21564 7880 21570
rect 7748 21558 7880 21564
rect 9680 21558 9732 21564
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 7380 21548 7432 21554
rect 7760 21542 7880 21558
rect 7380 21490 7432 21496
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1504 20505 1532 20742
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 1490 20496 1546 20505
rect 1490 20431 1546 20440
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 7024 19922 7052 20946
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7116 20602 7144 20878
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 7392 20466 7420 21490
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7576 21146 7604 21354
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 7484 20534 7512 20742
rect 7472 20528 7524 20534
rect 7472 20470 7524 20476
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7392 19990 7420 20402
rect 7668 20058 7696 20402
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7380 19984 7432 19990
rect 7380 19926 7432 19932
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 7760 19718 7788 20742
rect 7852 20466 7880 21542
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 7932 21072 7984 21078
rect 7932 21014 7984 21020
rect 7944 20602 7972 21014
rect 8220 21010 8248 21286
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7852 19922 7880 20402
rect 7944 20058 7972 20538
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 8220 19854 8248 20946
rect 8576 20868 8628 20874
rect 8576 20810 8628 20816
rect 8588 20398 8616 20810
rect 9692 20534 9720 21558
rect 13004 21010 13032 22102
rect 14108 22098 14136 22442
rect 14384 22438 14412 24142
rect 14476 23662 14504 24534
rect 14752 24274 14780 25094
rect 14936 24410 14964 25350
rect 16580 25298 16632 25304
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 16592 25242 16620 25298
rect 16960 25294 16988 25978
rect 17592 25900 17644 25906
rect 17592 25842 17644 25848
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17316 25832 17368 25838
rect 17316 25774 17368 25780
rect 16948 25288 17000 25294
rect 15028 24614 15056 25230
rect 16592 25214 16712 25242
rect 16948 25230 17000 25236
rect 15108 24812 15160 24818
rect 15108 24754 15160 24760
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14936 24070 14964 24346
rect 15028 24138 15056 24550
rect 15120 24410 15148 24754
rect 15108 24404 15160 24410
rect 15108 24346 15160 24352
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 14924 24064 14976 24070
rect 14924 24006 14976 24012
rect 14464 23656 14516 23662
rect 14464 23598 14516 23604
rect 14476 23118 14504 23598
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14476 22778 14504 23054
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14096 22092 14148 22098
rect 14384 22094 14412 22374
rect 14096 22034 14148 22040
rect 14292 22066 14412 22094
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 13924 21622 13952 21830
rect 13452 21616 13504 21622
rect 13452 21558 13504 21564
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 13464 21298 13492 21558
rect 14292 21486 14320 22066
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 13464 21270 13584 21298
rect 12992 21004 13044 21010
rect 12992 20946 13044 20952
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 10600 20800 10652 20806
rect 10600 20742 10652 20748
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 9680 20528 9732 20534
rect 10140 20528 10192 20534
rect 9680 20470 9732 20476
rect 10060 20476 10140 20482
rect 10060 20470 10192 20476
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9508 19854 9536 20334
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 848 19712 900 19718
rect 846 19680 848 19689
rect 7472 19712 7524 19718
rect 900 19680 902 19689
rect 7472 19654 7524 19660
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 846 19615 902 19624
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 7484 19378 7512 19654
rect 7760 19378 7788 19654
rect 7852 19378 7880 19722
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 7300 18698 7328 19110
rect 7852 18970 7880 19314
rect 9508 19310 9536 19790
rect 9692 19718 9720 20470
rect 10060 20454 10180 20470
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9876 20058 9904 20198
rect 10060 20058 10088 20454
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 10152 20058 10180 20334
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 10428 19786 10456 20198
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 10612 19378 10640 20742
rect 10704 20398 10732 20742
rect 11532 20534 11560 20878
rect 13556 20806 13584 21270
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20534 13584 20742
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 12072 20528 12124 20534
rect 12072 20470 12124 20476
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10980 19922 11008 20334
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 12084 19514 12112 20470
rect 14292 19922 14320 21422
rect 14936 21146 14964 24006
rect 16684 23662 16712 25214
rect 17328 25158 17356 25774
rect 17604 25378 17632 25842
rect 17684 25696 17736 25702
rect 17684 25638 17736 25644
rect 17696 25514 17724 25638
rect 17696 25486 17816 25514
rect 17684 25424 17736 25430
rect 17604 25372 17684 25378
rect 17604 25366 17736 25372
rect 17604 25350 17724 25366
rect 17696 25294 17724 25350
rect 17684 25288 17736 25294
rect 17684 25230 17736 25236
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 17316 25152 17368 25158
rect 17316 25094 17368 25100
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 16868 24818 16896 25094
rect 17328 24818 17356 25094
rect 17420 24954 17448 25094
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 16672 23656 16724 23662
rect 16672 23598 16724 23604
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 15488 22710 15516 23122
rect 16684 23050 16712 23598
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 16684 22574 16712 22986
rect 16960 22982 16988 23666
rect 17052 23254 17080 23666
rect 17236 23594 17264 24142
rect 17224 23588 17276 23594
rect 17224 23530 17276 23536
rect 17512 23322 17540 24142
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17604 23798 17632 24006
rect 17696 23866 17724 25230
rect 17788 25158 17816 25486
rect 17972 25294 18000 25842
rect 17960 25288 18012 25294
rect 17960 25230 18012 25236
rect 17868 25220 17920 25226
rect 17868 25162 17920 25168
rect 17776 25152 17828 25158
rect 17776 25094 17828 25100
rect 17788 24818 17816 25094
rect 17880 24954 17908 25162
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 17776 24812 17828 24818
rect 17776 24754 17828 24760
rect 17684 23860 17736 23866
rect 17684 23802 17736 23808
rect 17592 23792 17644 23798
rect 17592 23734 17644 23740
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 17500 23316 17552 23322
rect 17500 23258 17552 23264
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 16948 22976 17000 22982
rect 16948 22918 17000 22924
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 15108 22568 15160 22574
rect 15108 22510 15160 22516
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16948 22568 17000 22574
rect 16948 22510 17000 22516
rect 15120 22234 15148 22510
rect 16960 22234 16988 22510
rect 15108 22228 15160 22234
rect 15108 22170 15160 22176
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 17144 22030 17172 22714
rect 17512 22098 17540 23258
rect 17604 22982 17632 23598
rect 17696 23050 17724 23802
rect 17788 23322 17816 24754
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 17684 23044 17736 23050
rect 17684 22986 17736 22992
rect 17592 22976 17644 22982
rect 17592 22918 17644 22924
rect 17880 22778 17908 24686
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17972 22574 18000 25230
rect 18064 24954 18092 26030
rect 18156 25242 18184 26726
rect 18248 25362 18276 26862
rect 19064 25696 19116 25702
rect 19064 25638 19116 25644
rect 18236 25356 18288 25362
rect 18236 25298 18288 25304
rect 19076 25294 19104 25638
rect 18328 25288 18380 25294
rect 18156 25214 18276 25242
rect 18328 25230 18380 25236
rect 19064 25288 19116 25294
rect 19064 25230 19116 25236
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18052 24948 18104 24954
rect 18052 24890 18104 24896
rect 18064 23798 18092 24890
rect 18156 24682 18184 25094
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18052 23792 18104 23798
rect 18052 23734 18104 23740
rect 18064 22642 18092 23734
rect 18248 23186 18276 25214
rect 18340 25158 18368 25230
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 18512 25152 18564 25158
rect 18512 25094 18564 25100
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18340 24614 18368 25094
rect 18524 24818 18552 25094
rect 18616 24954 18644 25094
rect 18604 24948 18656 24954
rect 18604 24890 18656 24896
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18524 24206 18552 24754
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 18248 22710 18276 23122
rect 19168 23050 19196 29124
rect 19340 29106 19392 29112
rect 19340 28688 19392 28694
rect 19340 28630 19392 28636
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 19260 23662 19288 24550
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19352 23322 19380 28630
rect 19996 28558 20024 29650
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 20088 29306 20116 29582
rect 20076 29300 20128 29306
rect 20076 29242 20128 29248
rect 20180 28694 20208 31690
rect 20352 31408 20404 31414
rect 20352 31350 20404 31356
rect 20364 31142 20392 31350
rect 20352 31136 20404 31142
rect 20352 31078 20404 31084
rect 20260 29844 20312 29850
rect 20260 29786 20312 29792
rect 20168 28688 20220 28694
rect 20168 28630 20220 28636
rect 19984 28552 20036 28558
rect 20036 28500 20116 28506
rect 19984 28494 20116 28500
rect 19996 28478 20116 28494
rect 20272 28490 20300 29786
rect 20364 29102 20392 31078
rect 21468 29714 21496 31826
rect 27356 30802 27384 32506
rect 27712 32224 27764 32230
rect 27712 32166 27764 32172
rect 27724 31822 27752 32166
rect 28000 31822 28028 32710
rect 28368 32434 28396 33934
rect 28460 33522 28488 34070
rect 28644 33998 28672 35090
rect 28736 34678 28764 35090
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 30196 35080 30248 35086
rect 30196 35022 30248 35028
rect 28724 34672 28776 34678
rect 28724 34614 28776 34620
rect 29736 34468 29788 34474
rect 29736 34410 29788 34416
rect 29748 33998 29776 34410
rect 29932 34406 29960 35022
rect 30208 34746 30236 35022
rect 31576 35012 31628 35018
rect 31576 34954 31628 34960
rect 30196 34740 30248 34746
rect 30196 34682 30248 34688
rect 29920 34400 29972 34406
rect 29920 34342 29972 34348
rect 28632 33992 28684 33998
rect 28632 33934 28684 33940
rect 29736 33992 29788 33998
rect 29736 33934 29788 33940
rect 28644 33522 28672 33934
rect 29092 33924 29144 33930
rect 29092 33866 29144 33872
rect 29104 33658 29132 33866
rect 29460 33856 29512 33862
rect 29460 33798 29512 33804
rect 29092 33652 29144 33658
rect 29092 33594 29144 33600
rect 29000 33584 29052 33590
rect 29000 33526 29052 33532
rect 28448 33516 28500 33522
rect 28448 33458 28500 33464
rect 28632 33516 28684 33522
rect 28632 33458 28684 33464
rect 29012 32978 29040 33526
rect 29472 33454 29500 33798
rect 29932 33590 29960 34342
rect 30208 34066 30236 34682
rect 31588 34678 31616 34954
rect 31576 34672 31628 34678
rect 31576 34614 31628 34620
rect 30196 34060 30248 34066
rect 30196 34002 30248 34008
rect 29920 33584 29972 33590
rect 29920 33526 29972 33532
rect 29460 33448 29512 33454
rect 29460 33390 29512 33396
rect 29736 33312 29788 33318
rect 29736 33254 29788 33260
rect 29000 32972 29052 32978
rect 29000 32914 29052 32920
rect 29012 32434 29040 32914
rect 29184 32904 29236 32910
rect 29184 32846 29236 32852
rect 28356 32428 28408 32434
rect 28356 32370 28408 32376
rect 29000 32428 29052 32434
rect 29000 32370 29052 32376
rect 28368 31958 28396 32370
rect 29196 32366 29224 32846
rect 29368 32836 29420 32842
rect 29368 32778 29420 32784
rect 29184 32360 29236 32366
rect 29184 32302 29236 32308
rect 29380 32230 29408 32778
rect 29748 32434 29776 33254
rect 29736 32428 29788 32434
rect 29736 32370 29788 32376
rect 29932 32366 29960 33526
rect 30208 32978 30236 34002
rect 31588 33998 31616 34614
rect 32232 34610 32260 36314
rect 33244 35834 33272 36654
rect 33508 36576 33560 36582
rect 33508 36518 33560 36524
rect 33520 36242 33548 36518
rect 33888 36242 33916 36654
rect 34164 36378 34192 36654
rect 36084 36644 36136 36650
rect 36084 36586 36136 36592
rect 35716 36576 35768 36582
rect 35716 36518 35768 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34152 36372 34204 36378
rect 34152 36314 34204 36320
rect 34704 36304 34756 36310
rect 34704 36246 34756 36252
rect 33508 36236 33560 36242
rect 33508 36178 33560 36184
rect 33876 36236 33928 36242
rect 33876 36178 33928 36184
rect 32680 35828 32732 35834
rect 32680 35770 32732 35776
rect 33232 35828 33284 35834
rect 33232 35770 33284 35776
rect 32692 35714 32720 35770
rect 32692 35698 32812 35714
rect 32404 35692 32456 35698
rect 32692 35692 32824 35698
rect 32692 35686 32772 35692
rect 32404 35634 32456 35640
rect 32772 35634 32824 35640
rect 32416 35578 32444 35634
rect 32324 35550 32444 35578
rect 32220 34604 32272 34610
rect 32220 34546 32272 34552
rect 31944 34400 31996 34406
rect 31944 34342 31996 34348
rect 31576 33992 31628 33998
rect 31576 33934 31628 33940
rect 30380 33924 30432 33930
rect 30380 33866 30432 33872
rect 30392 33658 30420 33866
rect 30380 33652 30432 33658
rect 30380 33594 30432 33600
rect 31956 33386 31984 34342
rect 32232 33998 32260 34546
rect 32324 34542 32352 35550
rect 32784 34950 32812 35634
rect 32496 34944 32548 34950
rect 32496 34886 32548 34892
rect 32772 34944 32824 34950
rect 32772 34886 32824 34892
rect 32508 34542 32536 34886
rect 33888 34678 33916 36178
rect 34612 36032 34664 36038
rect 34612 35974 34664 35980
rect 34520 34944 34572 34950
rect 34520 34886 34572 34892
rect 33876 34672 33928 34678
rect 33876 34614 33928 34620
rect 32312 34536 32364 34542
rect 32496 34536 32548 34542
rect 32312 34478 32364 34484
rect 32416 34484 32496 34490
rect 32416 34478 32548 34484
rect 32588 34536 32640 34542
rect 32588 34478 32640 34484
rect 32220 33992 32272 33998
rect 32220 33934 32272 33940
rect 32036 33856 32088 33862
rect 32036 33798 32088 33804
rect 32048 33522 32076 33798
rect 32232 33590 32260 33934
rect 32324 33862 32352 34478
rect 32416 34462 32536 34478
rect 32416 33862 32444 34462
rect 32600 34066 32628 34478
rect 34532 34406 34560 34886
rect 34624 34746 34652 35974
rect 34716 35290 34744 36246
rect 35164 36168 35216 36174
rect 35164 36110 35216 36116
rect 35176 35834 35204 36110
rect 35728 36106 35756 36518
rect 36096 36174 36124 36586
rect 36188 36242 36216 36654
rect 36176 36236 36228 36242
rect 36176 36178 36228 36184
rect 36084 36168 36136 36174
rect 36084 36110 36136 36116
rect 35716 36100 35768 36106
rect 35716 36042 35768 36048
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 35164 35828 35216 35834
rect 35164 35770 35216 35776
rect 35348 35828 35400 35834
rect 35348 35770 35400 35776
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34704 35284 34756 35290
rect 34704 35226 34756 35232
rect 35256 34944 35308 34950
rect 35256 34886 35308 34892
rect 34612 34740 34664 34746
rect 34612 34682 34664 34688
rect 35268 34678 35296 34886
rect 35360 34678 35388 35770
rect 36188 35154 36216 36178
rect 36280 35834 36308 36858
rect 36360 36848 36412 36854
rect 36360 36790 36412 36796
rect 36820 36848 36872 36854
rect 36820 36790 36872 36796
rect 36372 36038 36400 36790
rect 36728 36100 36780 36106
rect 36728 36042 36780 36048
rect 36360 36032 36412 36038
rect 36360 35974 36412 35980
rect 36268 35828 36320 35834
rect 36268 35770 36320 35776
rect 36372 35698 36400 35974
rect 36360 35692 36412 35698
rect 36360 35634 36412 35640
rect 36740 35562 36768 36042
rect 36832 35834 36860 36790
rect 37464 36780 37516 36786
rect 37464 36722 37516 36728
rect 37280 36576 37332 36582
rect 37280 36518 37332 36524
rect 36820 35828 36872 35834
rect 36820 35770 36872 35776
rect 37292 35698 37320 36518
rect 37476 36106 37504 36722
rect 38476 36712 38528 36718
rect 38476 36654 38528 36660
rect 38488 36378 38516 36654
rect 38476 36372 38528 36378
rect 38476 36314 38528 36320
rect 39212 36372 39264 36378
rect 39212 36314 39264 36320
rect 39028 36304 39080 36310
rect 39028 36246 39080 36252
rect 38200 36236 38252 36242
rect 38200 36178 38252 36184
rect 37464 36100 37516 36106
rect 37464 36042 37516 36048
rect 37280 35692 37332 35698
rect 37280 35634 37332 35640
rect 36728 35556 36780 35562
rect 36728 35498 36780 35504
rect 36176 35148 36228 35154
rect 36176 35090 36228 35096
rect 35440 35080 35492 35086
rect 35440 35022 35492 35028
rect 35256 34672 35308 34678
rect 35256 34614 35308 34620
rect 35348 34672 35400 34678
rect 35348 34614 35400 34620
rect 35348 34536 35400 34542
rect 35348 34478 35400 34484
rect 34520 34400 34572 34406
rect 34520 34342 34572 34348
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 32588 34060 32640 34066
rect 32588 34002 32640 34008
rect 32312 33856 32364 33862
rect 32312 33798 32364 33804
rect 32404 33856 32456 33862
rect 32404 33798 32456 33804
rect 32220 33584 32272 33590
rect 32220 33526 32272 33532
rect 32416 33522 32444 33798
rect 32600 33522 32628 34002
rect 35360 33998 35388 34478
rect 35348 33992 35400 33998
rect 35348 33934 35400 33940
rect 33048 33924 33100 33930
rect 33048 33866 33100 33872
rect 35256 33924 35308 33930
rect 35256 33866 35308 33872
rect 32036 33516 32088 33522
rect 32036 33458 32088 33464
rect 32404 33516 32456 33522
rect 32404 33458 32456 33464
rect 32588 33516 32640 33522
rect 32588 33458 32640 33464
rect 31944 33380 31996 33386
rect 31944 33322 31996 33328
rect 33060 33318 33088 33866
rect 33692 33856 33744 33862
rect 33692 33798 33744 33804
rect 32036 33312 32088 33318
rect 32036 33254 32088 33260
rect 33048 33312 33100 33318
rect 33048 33254 33100 33260
rect 30288 33108 30340 33114
rect 30288 33050 30340 33056
rect 30196 32972 30248 32978
rect 30196 32914 30248 32920
rect 30208 32570 30236 32914
rect 30300 32570 30328 33050
rect 32048 32910 32076 33254
rect 33060 32978 33088 33254
rect 33048 32972 33100 32978
rect 33048 32914 33100 32920
rect 32036 32904 32088 32910
rect 32036 32846 32088 32852
rect 32128 32904 32180 32910
rect 32128 32846 32180 32852
rect 30196 32564 30248 32570
rect 30196 32506 30248 32512
rect 30288 32564 30340 32570
rect 30288 32506 30340 32512
rect 30012 32428 30064 32434
rect 30012 32370 30064 32376
rect 29920 32360 29972 32366
rect 29920 32302 29972 32308
rect 28816 32224 28868 32230
rect 28816 32166 28868 32172
rect 29368 32224 29420 32230
rect 29368 32166 29420 32172
rect 28356 31952 28408 31958
rect 28356 31894 28408 31900
rect 27712 31816 27764 31822
rect 27712 31758 27764 31764
rect 27988 31816 28040 31822
rect 27988 31758 28040 31764
rect 27724 31278 27752 31758
rect 27712 31272 27764 31278
rect 27712 31214 27764 31220
rect 27620 31136 27672 31142
rect 27620 31078 27672 31084
rect 27632 30802 27660 31078
rect 27344 30796 27396 30802
rect 27344 30738 27396 30744
rect 27620 30796 27672 30802
rect 27620 30738 27672 30744
rect 28368 30666 28396 31894
rect 28828 31822 28856 32166
rect 28816 31816 28868 31822
rect 28816 31758 28868 31764
rect 28828 31482 28856 31758
rect 28816 31476 28868 31482
rect 28816 31418 28868 31424
rect 29092 31340 29144 31346
rect 29092 31282 29144 31288
rect 29104 30938 29132 31282
rect 29092 30932 29144 30938
rect 29092 30874 29144 30880
rect 28356 30660 28408 30666
rect 28356 30602 28408 30608
rect 28368 30122 28396 30602
rect 28356 30116 28408 30122
rect 28356 30058 28408 30064
rect 22376 29844 22428 29850
rect 22376 29786 22428 29792
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 21456 29708 21508 29714
rect 21456 29650 21508 29656
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 20456 29238 20484 29446
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20824 29170 20852 29650
rect 22388 29170 22416 29786
rect 28368 29578 28396 30058
rect 28356 29572 28408 29578
rect 28356 29514 28408 29520
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 22376 29164 22428 29170
rect 22376 29106 22428 29112
rect 20352 29096 20404 29102
rect 20352 29038 20404 29044
rect 20444 28688 20496 28694
rect 20444 28630 20496 28636
rect 20628 28688 20680 28694
rect 20628 28630 20680 28636
rect 20352 28620 20404 28626
rect 20352 28562 20404 28568
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19996 28150 20024 28358
rect 20088 28150 20116 28478
rect 20260 28484 20312 28490
rect 20260 28426 20312 28432
rect 20364 28218 20392 28562
rect 20352 28212 20404 28218
rect 20352 28154 20404 28160
rect 19984 28144 20036 28150
rect 19984 28086 20036 28092
rect 20076 28144 20128 28150
rect 20076 28086 20128 28092
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19444 27470 19472 27814
rect 20180 27538 20208 28018
rect 20168 27532 20220 27538
rect 20168 27474 20220 27480
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19444 26330 19472 27406
rect 20180 27130 20208 27474
rect 20364 27334 20392 28154
rect 20352 27328 20404 27334
rect 20352 27270 20404 27276
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 20180 26382 20208 27066
rect 20364 26586 20392 27270
rect 20456 26994 20484 28630
rect 20536 28484 20588 28490
rect 20536 28426 20588 28432
rect 20548 28218 20576 28426
rect 20536 28212 20588 28218
rect 20536 28154 20588 28160
rect 20640 27402 20668 28630
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 21916 27396 21968 27402
rect 21916 27338 21968 27344
rect 20640 26994 20668 27338
rect 21928 27130 21956 27338
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 21916 27124 21968 27130
rect 21916 27066 21968 27072
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20168 26376 20220 26382
rect 19444 26302 19564 26330
rect 20168 26318 20220 26324
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19444 25974 19472 26182
rect 19432 25968 19484 25974
rect 19432 25910 19484 25916
rect 19536 25906 19564 26302
rect 20640 25906 20668 26386
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 19524 25900 19576 25906
rect 19524 25842 19576 25848
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20076 25832 20128 25838
rect 20076 25774 20128 25780
rect 20088 24954 20116 25774
rect 20640 25498 20668 25842
rect 20732 25770 20760 26250
rect 21364 26240 21416 26246
rect 21364 26182 21416 26188
rect 21376 25974 21404 26182
rect 22848 25974 22876 27270
rect 21364 25968 21416 25974
rect 21364 25910 21416 25916
rect 22836 25968 22888 25974
rect 22836 25910 22888 25916
rect 20720 25764 20772 25770
rect 20720 25706 20772 25712
rect 20628 25492 20680 25498
rect 20628 25434 20680 25440
rect 20076 24948 20128 24954
rect 20076 24890 20128 24896
rect 20640 24886 20668 25434
rect 20628 24880 20680 24886
rect 20628 24822 20680 24828
rect 20732 24614 20760 25706
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 21088 24200 21140 24206
rect 21088 24142 21140 24148
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19536 23730 19564 24006
rect 21100 23866 21128 24142
rect 22848 23866 22876 25910
rect 23584 25838 23612 27406
rect 29184 26036 29236 26042
rect 29184 25978 29236 25984
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 28448 25832 28500 25838
rect 28448 25774 28500 25780
rect 23584 25362 23612 25774
rect 27712 25492 27764 25498
rect 27712 25434 27764 25440
rect 23572 25356 23624 25362
rect 23572 25298 23624 25304
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 19524 23724 19576 23730
rect 19524 23666 19576 23672
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19156 23044 19208 23050
rect 19156 22986 19208 22992
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 18236 22704 18288 22710
rect 18236 22646 18288 22652
rect 18616 22642 18644 22918
rect 19260 22778 19288 22918
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 17960 22568 18012 22574
rect 17960 22510 18012 22516
rect 18616 22098 18644 22578
rect 17500 22092 17552 22098
rect 17500 22034 17552 22040
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 19352 20534 19380 23258
rect 27724 22094 27752 25434
rect 28460 25226 28488 25774
rect 29196 25770 29224 25978
rect 29184 25764 29236 25770
rect 29184 25706 29236 25712
rect 28448 25220 28500 25226
rect 28448 25162 28500 25168
rect 28460 24818 28488 25162
rect 29196 24886 29224 25706
rect 29380 25498 29408 32166
rect 30024 31754 30052 32370
rect 30208 31872 30236 32506
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 30392 32026 30420 32302
rect 30380 32020 30432 32026
rect 30380 31962 30432 31968
rect 30380 31884 30432 31890
rect 30208 31844 30380 31872
rect 30012 31748 30064 31754
rect 30012 31690 30064 31696
rect 29920 31680 29972 31686
rect 29920 31622 29972 31628
rect 29932 31278 29960 31622
rect 30024 31414 30052 31690
rect 30012 31408 30064 31414
rect 30012 31350 30064 31356
rect 29920 31272 29972 31278
rect 29920 31214 29972 31220
rect 29736 31204 29788 31210
rect 29736 31146 29788 31152
rect 29748 30258 29776 31146
rect 29932 31142 29960 31214
rect 29920 31136 29972 31142
rect 29920 31078 29972 31084
rect 29736 30252 29788 30258
rect 29736 30194 29788 30200
rect 29552 30048 29604 30054
rect 29552 29990 29604 29996
rect 29564 29170 29592 29990
rect 30208 29714 30236 31844
rect 30380 31826 30432 31832
rect 30748 31680 30800 31686
rect 30748 31622 30800 31628
rect 30760 31482 30788 31622
rect 30748 31476 30800 31482
rect 30748 31418 30800 31424
rect 31312 31210 31340 32370
rect 31392 32224 31444 32230
rect 31392 32166 31444 32172
rect 31404 32026 31432 32166
rect 31392 32020 31444 32026
rect 31392 31962 31444 31968
rect 31576 31272 31628 31278
rect 31576 31214 31628 31220
rect 31300 31204 31352 31210
rect 31300 31146 31352 31152
rect 31588 30938 31616 31214
rect 31576 30932 31628 30938
rect 31576 30874 31628 30880
rect 32140 30870 32168 32846
rect 33060 32570 33088 32914
rect 33704 32910 33732 33798
rect 35268 33590 35296 33866
rect 35452 33862 35480 35022
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 36188 34746 36216 35090
rect 36268 35012 36320 35018
rect 36268 34954 36320 34960
rect 36280 34746 36308 34954
rect 36176 34740 36228 34746
rect 36176 34682 36228 34688
rect 36268 34740 36320 34746
rect 36268 34682 36320 34688
rect 35532 34604 35584 34610
rect 35532 34546 35584 34552
rect 35544 34134 35572 34546
rect 35532 34128 35584 34134
rect 35532 34070 35584 34076
rect 35544 33998 35572 34070
rect 36188 33998 36216 34682
rect 37280 34400 37332 34406
rect 37280 34342 37332 34348
rect 37292 34066 37320 34342
rect 37476 34218 37504 36042
rect 38016 36032 38068 36038
rect 38016 35974 38068 35980
rect 38028 35766 38056 35974
rect 38016 35760 38068 35766
rect 38016 35702 38068 35708
rect 38212 35698 38240 36178
rect 39040 36174 39068 36246
rect 39224 36174 39252 36314
rect 39028 36168 39080 36174
rect 39028 36110 39080 36116
rect 39212 36168 39264 36174
rect 39212 36110 39264 36116
rect 38384 36100 38436 36106
rect 38384 36042 38436 36048
rect 38396 35698 38424 36042
rect 39040 35714 39068 36110
rect 39120 36032 39172 36038
rect 39120 35974 39172 35980
rect 39132 35834 39160 35974
rect 39120 35828 39172 35834
rect 39120 35770 39172 35776
rect 38200 35692 38252 35698
rect 38200 35634 38252 35640
rect 38384 35692 38436 35698
rect 39040 35686 39160 35714
rect 38384 35634 38436 35640
rect 38212 34610 38240 35634
rect 38568 35080 38620 35086
rect 38568 35022 38620 35028
rect 38200 34604 38252 34610
rect 38200 34546 38252 34552
rect 37384 34190 37504 34218
rect 38212 34202 38240 34546
rect 38200 34196 38252 34202
rect 37280 34060 37332 34066
rect 37280 34002 37332 34008
rect 35532 33992 35584 33998
rect 35532 33934 35584 33940
rect 36084 33992 36136 33998
rect 36084 33934 36136 33940
rect 36176 33992 36228 33998
rect 36176 33934 36228 33940
rect 35440 33856 35492 33862
rect 35440 33798 35492 33804
rect 35256 33584 35308 33590
rect 35256 33526 35308 33532
rect 35452 33522 35480 33798
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 35440 33516 35492 33522
rect 35440 33458 35492 33464
rect 35992 33516 36044 33522
rect 35992 33458 36044 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 33968 33108 34020 33114
rect 33968 33050 34020 33056
rect 33692 32904 33744 32910
rect 33692 32846 33744 32852
rect 33048 32564 33100 32570
rect 33048 32506 33100 32512
rect 33980 32502 34008 33050
rect 35348 32768 35400 32774
rect 35348 32710 35400 32716
rect 33968 32496 34020 32502
rect 33968 32438 34020 32444
rect 32864 32428 32916 32434
rect 32864 32370 32916 32376
rect 32876 31754 32904 32370
rect 34704 32360 34756 32366
rect 34704 32302 34756 32308
rect 34716 32026 34744 32302
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34704 32020 34756 32026
rect 34704 31962 34756 31968
rect 35360 31822 35388 32710
rect 35452 32026 35480 33458
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 36004 32366 36032 33458
rect 36096 33454 36124 33934
rect 36084 33448 36136 33454
rect 36084 33390 36136 33396
rect 36188 32978 36216 33934
rect 37384 33930 37412 34190
rect 38200 34138 38252 34144
rect 38580 34134 38608 35022
rect 38752 34944 38804 34950
rect 38752 34886 38804 34892
rect 38568 34128 38620 34134
rect 38568 34070 38620 34076
rect 37372 33924 37424 33930
rect 37372 33866 37424 33872
rect 36360 33856 36412 33862
rect 36360 33798 36412 33804
rect 36372 33522 36400 33798
rect 36360 33516 36412 33522
rect 36360 33458 36412 33464
rect 37004 33516 37056 33522
rect 37004 33458 37056 33464
rect 36372 33114 36400 33458
rect 37016 33114 37044 33458
rect 37280 33312 37332 33318
rect 37280 33254 37332 33260
rect 36360 33108 36412 33114
rect 36360 33050 36412 33056
rect 36912 33108 36964 33114
rect 36912 33050 36964 33056
rect 37004 33108 37056 33114
rect 37004 33050 37056 33056
rect 36924 32994 36952 33050
rect 36176 32972 36228 32978
rect 36924 32966 37136 32994
rect 36176 32914 36228 32920
rect 36188 32570 36216 32914
rect 37108 32910 37136 32966
rect 37096 32904 37148 32910
rect 37096 32846 37148 32852
rect 36176 32564 36228 32570
rect 36176 32506 36228 32512
rect 35992 32360 36044 32366
rect 35992 32302 36044 32308
rect 36176 32224 36228 32230
rect 36176 32166 36228 32172
rect 35440 32020 35492 32026
rect 35440 31962 35492 31968
rect 36188 31890 36216 32166
rect 36176 31884 36228 31890
rect 36176 31826 36228 31832
rect 37292 31822 37320 33254
rect 37384 32502 37412 33866
rect 38108 33516 38160 33522
rect 38108 33458 38160 33464
rect 37740 33312 37792 33318
rect 37740 33254 37792 33260
rect 37752 32978 37780 33254
rect 38120 33114 38148 33458
rect 38108 33108 38160 33114
rect 38108 33050 38160 33056
rect 37740 32972 37792 32978
rect 37740 32914 37792 32920
rect 37372 32496 37424 32502
rect 37372 32438 37424 32444
rect 35348 31816 35400 31822
rect 35348 31758 35400 31764
rect 37280 31816 37332 31822
rect 37280 31758 37332 31764
rect 32876 31726 32996 31754
rect 32128 30864 32180 30870
rect 32128 30806 32180 30812
rect 31300 30728 31352 30734
rect 31300 30670 31352 30676
rect 32128 30728 32180 30734
rect 32128 30670 32180 30676
rect 30380 30592 30432 30598
rect 30380 30534 30432 30540
rect 30392 30258 30420 30534
rect 30380 30252 30432 30258
rect 30380 30194 30432 30200
rect 30288 30048 30340 30054
rect 30288 29990 30340 29996
rect 30196 29708 30248 29714
rect 30196 29650 30248 29656
rect 30300 29578 30328 29990
rect 30104 29572 30156 29578
rect 30104 29514 30156 29520
rect 30288 29572 30340 29578
rect 30288 29514 30340 29520
rect 30116 29306 30144 29514
rect 30104 29300 30156 29306
rect 30104 29242 30156 29248
rect 29552 29164 29604 29170
rect 29552 29106 29604 29112
rect 30392 29034 30420 30194
rect 31312 30190 31340 30670
rect 32140 30258 32168 30670
rect 32968 30666 32996 31726
rect 36728 31680 36780 31686
rect 36728 31622 36780 31628
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 36740 31414 36768 31622
rect 37384 31498 37412 32438
rect 38580 31754 38608 34070
rect 38764 32978 38792 34886
rect 39132 34202 39160 35686
rect 39120 34196 39172 34202
rect 39120 34138 39172 34144
rect 38936 33992 38988 33998
rect 38936 33934 38988 33940
rect 38948 33658 38976 33934
rect 38936 33652 38988 33658
rect 38936 33594 38988 33600
rect 38948 33114 38976 33594
rect 38936 33108 38988 33114
rect 38936 33050 38988 33056
rect 38752 32972 38804 32978
rect 38752 32914 38804 32920
rect 37292 31470 37412 31498
rect 38488 31726 38608 31754
rect 35992 31408 36044 31414
rect 35992 31350 36044 31356
rect 36728 31408 36780 31414
rect 36728 31350 36780 31356
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34244 30728 34296 30734
rect 34244 30670 34296 30676
rect 32956 30660 33008 30666
rect 32956 30602 33008 30608
rect 33968 30660 34020 30666
rect 33968 30602 34020 30608
rect 32968 30326 32996 30602
rect 33140 30592 33192 30598
rect 33140 30534 33192 30540
rect 32956 30320 33008 30326
rect 32956 30262 33008 30268
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 31300 30184 31352 30190
rect 31300 30126 31352 30132
rect 31312 29850 31340 30126
rect 31760 30048 31812 30054
rect 31760 29990 31812 29996
rect 31300 29844 31352 29850
rect 31300 29786 31352 29792
rect 31576 29504 31628 29510
rect 31576 29446 31628 29452
rect 31588 29170 31616 29446
rect 31772 29170 31800 29990
rect 32140 29714 32168 30194
rect 32128 29708 32180 29714
rect 32128 29650 32180 29656
rect 32140 29306 32168 29650
rect 32968 29578 32996 30262
rect 33152 30258 33180 30534
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 33980 30054 34008 30602
rect 34256 30258 34284 30670
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 36004 30326 36032 31350
rect 37292 31346 37320 31470
rect 37372 31408 37424 31414
rect 37372 31350 37424 31356
rect 37280 31340 37332 31346
rect 37280 31282 37332 31288
rect 36912 31136 36964 31142
rect 36912 31078 36964 31084
rect 36924 30938 36952 31078
rect 36912 30932 36964 30938
rect 36912 30874 36964 30880
rect 36452 30660 36504 30666
rect 36452 30602 36504 30608
rect 36084 30592 36136 30598
rect 36084 30534 36136 30540
rect 35992 30320 36044 30326
rect 35992 30262 36044 30268
rect 34244 30252 34296 30258
rect 34244 30194 34296 30200
rect 33968 30048 34020 30054
rect 33968 29990 34020 29996
rect 34256 29646 34284 30194
rect 34520 30184 34572 30190
rect 34520 30126 34572 30132
rect 34532 29850 34560 30126
rect 35900 30048 35952 30054
rect 35900 29990 35952 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34520 29844 34572 29850
rect 34520 29786 34572 29792
rect 35912 29714 35940 29990
rect 36004 29782 36032 30262
rect 36096 30054 36124 30534
rect 36464 30190 36492 30602
rect 36544 30592 36596 30598
rect 36544 30534 36596 30540
rect 36556 30258 36584 30534
rect 36544 30252 36596 30258
rect 36544 30194 36596 30200
rect 36452 30184 36504 30190
rect 36452 30126 36504 30132
rect 37292 30054 37320 31282
rect 37384 30938 37412 31350
rect 37464 31136 37516 31142
rect 37464 31078 37516 31084
rect 37372 30932 37424 30938
rect 37372 30874 37424 30880
rect 37476 30734 37504 31078
rect 37464 30728 37516 30734
rect 37464 30670 37516 30676
rect 37740 30728 37792 30734
rect 37740 30670 37792 30676
rect 37832 30728 37884 30734
rect 37832 30670 37884 30676
rect 37752 30598 37780 30670
rect 37648 30592 37700 30598
rect 37648 30534 37700 30540
rect 37740 30592 37792 30598
rect 37740 30534 37792 30540
rect 37660 30410 37688 30534
rect 37844 30410 37872 30670
rect 37660 30382 37872 30410
rect 36084 30048 36136 30054
rect 36084 29990 36136 29996
rect 36360 30048 36412 30054
rect 36360 29990 36412 29996
rect 37280 30048 37332 30054
rect 37280 29990 37332 29996
rect 35992 29776 36044 29782
rect 35992 29718 36044 29724
rect 36372 29714 36400 29990
rect 35900 29708 35952 29714
rect 35900 29650 35952 29656
rect 36360 29708 36412 29714
rect 36360 29650 36412 29656
rect 34244 29640 34296 29646
rect 34244 29582 34296 29588
rect 35992 29640 36044 29646
rect 35992 29582 36044 29588
rect 32956 29572 33008 29578
rect 32956 29514 33008 29520
rect 32128 29300 32180 29306
rect 32128 29242 32180 29248
rect 32968 29238 32996 29514
rect 32956 29232 33008 29238
rect 32956 29174 33008 29180
rect 34256 29170 34284 29582
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 31576 29164 31628 29170
rect 31576 29106 31628 29112
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 34244 29164 34296 29170
rect 34244 29106 34296 29112
rect 36004 29102 36032 29582
rect 37292 29510 37320 29990
rect 37660 29850 37688 30382
rect 37648 29844 37700 29850
rect 37648 29786 37700 29792
rect 38488 29510 38516 31726
rect 39132 31686 39160 34138
rect 39212 33448 39264 33454
rect 39212 33390 39264 33396
rect 39224 33046 39252 33390
rect 39212 33040 39264 33046
rect 39212 32982 39264 32988
rect 39120 31680 39172 31686
rect 39120 31622 39172 31628
rect 38660 31136 38712 31142
rect 38660 31078 38712 31084
rect 38672 30054 38700 31078
rect 38660 30048 38712 30054
rect 38660 29990 38712 29996
rect 38672 29578 38700 29990
rect 38660 29572 38712 29578
rect 38660 29514 38712 29520
rect 37280 29504 37332 29510
rect 37280 29446 37332 29452
rect 38476 29504 38528 29510
rect 38476 29446 38528 29452
rect 38672 29238 38700 29514
rect 38844 29504 38896 29510
rect 38844 29446 38896 29452
rect 38660 29232 38712 29238
rect 38660 29174 38712 29180
rect 38292 29164 38344 29170
rect 38292 29106 38344 29112
rect 35992 29096 36044 29102
rect 35992 29038 36044 29044
rect 30380 29028 30432 29034
rect 30380 28970 30432 28976
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 36004 28626 36032 29038
rect 38304 28762 38332 29106
rect 38384 28960 38436 28966
rect 38384 28902 38436 28908
rect 38292 28756 38344 28762
rect 38292 28698 38344 28704
rect 35992 28620 36044 28626
rect 35992 28562 36044 28568
rect 38396 28558 38424 28902
rect 38672 28778 38700 29174
rect 38672 28750 38792 28778
rect 38764 28694 38792 28750
rect 38752 28688 38804 28694
rect 38752 28630 38804 28636
rect 36728 28552 36780 28558
rect 36728 28494 36780 28500
rect 38384 28552 38436 28558
rect 38384 28494 38436 28500
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 32036 28008 32088 28014
rect 32036 27950 32088 27956
rect 33232 28008 33284 28014
rect 33232 27950 33284 27956
rect 35348 28008 35400 28014
rect 35348 27950 35400 27956
rect 31668 27532 31720 27538
rect 31668 27474 31720 27480
rect 31392 27124 31444 27130
rect 31392 27066 31444 27072
rect 31116 26580 31168 26586
rect 31116 26522 31168 26528
rect 30380 26376 30432 26382
rect 30380 26318 30432 26324
rect 30840 26376 30892 26382
rect 30840 26318 30892 26324
rect 29368 25492 29420 25498
rect 29368 25434 29420 25440
rect 29184 24880 29236 24886
rect 29184 24822 29236 24828
rect 30392 24834 30420 26318
rect 30564 26240 30616 26246
rect 30564 26182 30616 26188
rect 30576 25838 30604 26182
rect 30564 25832 30616 25838
rect 30564 25774 30616 25780
rect 30852 25498 30880 26318
rect 30840 25492 30892 25498
rect 30840 25434 30892 25440
rect 30932 25220 30984 25226
rect 30932 25162 30984 25168
rect 30840 24948 30892 24954
rect 30840 24890 30892 24896
rect 30392 24818 30512 24834
rect 28448 24812 28500 24818
rect 30392 24812 30524 24818
rect 30392 24806 30472 24812
rect 28448 24754 28500 24760
rect 30472 24754 30524 24760
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 28460 23730 28488 24754
rect 30484 24290 30512 24754
rect 30668 24410 30696 24754
rect 30656 24404 30708 24410
rect 30656 24346 30708 24352
rect 30484 24262 30696 24290
rect 30104 23860 30156 23866
rect 30104 23802 30156 23808
rect 28448 23724 28500 23730
rect 28448 23666 28500 23672
rect 28460 22642 28488 23666
rect 30012 23316 30064 23322
rect 30012 23258 30064 23264
rect 29828 23112 29880 23118
rect 29826 23080 29828 23089
rect 29920 23112 29972 23118
rect 29880 23080 29882 23089
rect 29920 23054 29972 23060
rect 29826 23015 29882 23024
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 29932 22574 29960 23054
rect 29552 22568 29604 22574
rect 29920 22568 29972 22574
rect 29552 22510 29604 22516
rect 29840 22516 29920 22522
rect 29840 22510 29972 22516
rect 29564 22098 29592 22510
rect 29840 22494 29960 22510
rect 29840 22234 29868 22494
rect 29920 22432 29972 22438
rect 29920 22374 29972 22380
rect 29828 22228 29880 22234
rect 29828 22170 29880 22176
rect 27724 22066 27936 22094
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 14556 20256 14608 20262
rect 14556 20198 14608 20204
rect 14568 19922 14596 20198
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12636 19378 12664 19790
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 13004 19446 13032 19654
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 14004 19440 14056 19446
rect 14004 19382 14056 19388
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 9312 18692 9364 18698
rect 9312 18634 9364 18640
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 9324 17134 9352 18634
rect 9508 17678 9536 18770
rect 10060 18766 10088 19246
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10244 18766 10272 19110
rect 10796 18970 10824 19110
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 9784 18290 9812 18702
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 9876 18290 9904 18566
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9508 17338 9536 17614
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9508 17202 9536 17274
rect 9692 17270 9720 18022
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 9508 16250 9536 17138
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 1308 16108 1360 16114
rect 1308 16050 1360 16056
rect 1320 15745 1348 16050
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8116 15972 8168 15978
rect 8116 15914 8168 15920
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 1306 15736 1362 15745
rect 4214 15739 4522 15748
rect 1306 15671 1362 15680
rect 8128 15502 8156 15914
rect 8312 15706 8340 15982
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 1412 15065 1440 15438
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 1398 15056 1454 15065
rect 7944 15026 7972 15370
rect 8128 15162 8156 15438
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 9508 15026 9536 16186
rect 9784 15094 9812 18226
rect 10704 17746 10732 18566
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 12728 17678 12756 19314
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13280 17746 13308 18022
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11164 17202 11192 17546
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 12452 17134 12480 17478
rect 12728 17270 12756 17614
rect 14016 17270 14044 19382
rect 14936 18698 14964 19654
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 14924 18692 14976 18698
rect 14924 18634 14976 18640
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14188 17604 14240 17610
rect 14188 17546 14240 17552
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 1398 14991 1454 15000
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 8576 15020 8628 15026
rect 9496 15020 9548 15026
rect 8576 14962 8628 14968
rect 9416 14980 9496 15008
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 7668 14414 7696 14962
rect 8588 14618 8616 14962
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 1216 14408 1268 14414
rect 1214 14376 1216 14385
rect 7656 14408 7708 14414
rect 1268 14376 1270 14385
rect 7656 14350 7708 14356
rect 1214 14311 1270 14320
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 7668 14074 7696 14350
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7852 14006 7880 14214
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 8588 13326 8616 14554
rect 9416 13870 9444 14980
rect 10796 15008 10824 17070
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12176 16590 12204 16934
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 11520 16516 11572 16522
rect 11520 16458 11572 16464
rect 11532 16114 11560 16458
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11808 15706 11836 15982
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 12176 15502 12204 16526
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12268 16046 12296 16118
rect 12544 16046 12572 16390
rect 12636 16250 12664 16594
rect 12728 16522 12756 17206
rect 14016 16998 14044 17206
rect 14200 17202 14228 17546
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 14292 17134 14320 18158
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 14752 17338 14780 17546
rect 14936 17542 14964 18634
rect 15108 17740 15160 17746
rect 15028 17700 15108 17728
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 13636 16516 13688 16522
rect 13636 16458 13688 16464
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 13372 15570 13400 16186
rect 13648 16046 13676 16458
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 10876 15020 10928 15026
rect 10796 14980 10876 15008
rect 9496 14962 9548 14968
rect 10876 14962 10928 14968
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 10888 14006 10916 14962
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 14006 11836 14214
rect 12268 14006 12296 14962
rect 12360 14414 12388 14962
rect 12452 14482 12480 15506
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13464 14482 13492 14894
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 13464 14074 13492 14418
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9416 13394 9444 13806
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 10888 13258 10916 13942
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 12728 12306 12756 14010
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12986 13860 13126
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 12728 11762 12756 12242
rect 13004 11830 13032 12582
rect 14016 12442 14044 16934
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14108 14550 14136 16730
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14292 15706 14320 15982
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 14292 14414 14320 14758
rect 14476 14414 14504 16934
rect 14936 16454 14964 17478
rect 15028 17134 15056 17700
rect 15108 17682 15160 17688
rect 15488 17338 15516 19450
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16592 19258 16620 19314
rect 16500 19230 16620 19258
rect 16500 18834 16528 19230
rect 17880 18834 17908 19654
rect 17972 19446 18000 19654
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 18524 18970 18552 19790
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 17868 18828 17920 18834
rect 17868 18770 17920 18776
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 16212 17808 16264 17814
rect 16212 17750 16264 17756
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15580 17338 15608 17478
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 16224 17134 16252 17750
rect 16500 17746 16528 18770
rect 17880 18290 17908 18770
rect 18616 18698 18644 18770
rect 19076 18766 19104 19110
rect 19260 18834 19288 19246
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 18604 18692 18656 18698
rect 18604 18634 18656 18640
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16500 17134 16528 17682
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 17316 17128 17368 17134
rect 17316 17070 17368 17076
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14936 16182 14964 16390
rect 14924 16176 14976 16182
rect 14924 16118 14976 16124
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14660 15502 14688 15846
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14936 14278 14964 16118
rect 15028 15570 15056 17070
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 15638 15516 15846
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15764 15570 15792 15982
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 16132 15706 16160 15914
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 15028 14328 15056 15506
rect 16500 14482 16528 17070
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17052 16250 17080 16934
rect 17328 16250 17356 17070
rect 17512 16726 17540 17614
rect 17972 17270 18000 18634
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 17144 15162 17172 16050
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 15108 14340 15160 14346
rect 15028 14300 15108 14328
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14476 12986 14504 14214
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14016 11830 14044 12378
rect 14844 11898 14872 12718
rect 14936 12238 14964 14214
rect 15028 12714 15056 14300
rect 15108 14282 15160 14288
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15212 14074 15240 14282
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 14074 16804 14214
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16868 13938 16896 14962
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 14482 16988 14894
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 17420 13938 17448 15846
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16408 13326 16436 13806
rect 17420 13326 17448 13874
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 16408 12714 16436 13262
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16960 12782 16988 13194
rect 17328 12850 17356 13262
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15580 11898 15608 12174
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 16960 11762 16988 12718
rect 17328 12442 17356 12786
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 17144 11218 17172 12242
rect 17512 12170 17540 16662
rect 18064 16590 18092 18566
rect 19260 18290 19288 18770
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 18604 18148 18656 18154
rect 18604 18090 18656 18096
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17696 16114 17724 16390
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17972 13938 18000 14554
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17972 13326 18000 13874
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18064 12850 18092 13670
rect 18156 13190 18184 17546
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 18340 16522 18368 17070
rect 18432 16658 18460 17682
rect 18616 17678 18644 18090
rect 19352 17814 19380 20470
rect 27908 20466 27936 22066
rect 29552 22092 29604 22098
rect 29552 22034 29604 22040
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 29748 21554 29776 21830
rect 29840 21690 29868 22170
rect 29932 22030 29960 22374
rect 30024 22234 30052 23258
rect 30116 23118 30144 23802
rect 30472 23656 30524 23662
rect 30472 23598 30524 23604
rect 30380 23520 30432 23526
rect 30380 23462 30432 23468
rect 30392 23322 30420 23462
rect 30484 23322 30512 23598
rect 30380 23316 30432 23322
rect 30380 23258 30432 23264
rect 30472 23316 30524 23322
rect 30472 23258 30524 23264
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 30104 23112 30156 23118
rect 30104 23054 30156 23060
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 30116 22642 30144 22918
rect 30104 22636 30156 22642
rect 30104 22578 30156 22584
rect 30196 22636 30248 22642
rect 30196 22578 30248 22584
rect 30104 22500 30156 22506
rect 30104 22442 30156 22448
rect 30012 22228 30064 22234
rect 30012 22170 30064 22176
rect 30116 22030 30144 22442
rect 30208 22438 30236 22578
rect 30196 22432 30248 22438
rect 30196 22374 30248 22380
rect 30196 22160 30248 22166
rect 30196 22102 30248 22108
rect 29920 22024 29972 22030
rect 30104 22024 30156 22030
rect 29920 21966 29972 21972
rect 30024 21984 30104 22012
rect 29828 21684 29880 21690
rect 29828 21626 29880 21632
rect 29736 21548 29788 21554
rect 29736 21490 29788 21496
rect 29920 21548 29972 21554
rect 30024 21536 30052 21984
rect 30104 21966 30156 21972
rect 30104 21616 30156 21622
rect 30104 21558 30156 21564
rect 29972 21508 30052 21536
rect 29920 21490 29972 21496
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 25412 20256 25464 20262
rect 25412 20198 25464 20204
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24596 19378 24624 19790
rect 24952 19440 25004 19446
rect 24952 19382 25004 19388
rect 24584 19372 24636 19378
rect 24584 19314 24636 19320
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 19340 17808 19392 17814
rect 19340 17750 19392 17756
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18984 16658 19012 17070
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17500 12164 17552 12170
rect 17500 12106 17552 12112
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 11830 17448 12038
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17696 11762 17724 12582
rect 18064 12238 18092 12786
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17972 11558 18000 12174
rect 18156 11830 18184 13126
rect 18340 12374 18368 14214
rect 18432 13462 18460 16594
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18524 16182 18552 16390
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 19812 15745 19840 18566
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19996 17746 20024 18022
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19996 17066 20024 17682
rect 20088 17678 20116 18226
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 19996 16590 20024 17002
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20088 16590 20116 16934
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 20364 16114 20392 18362
rect 21284 18290 21312 18566
rect 23860 18426 23888 18702
rect 24872 18426 24900 19246
rect 23848 18420 23900 18426
rect 23848 18362 23900 18368
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 24964 18306 24992 19382
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 21272 18284 21324 18290
rect 24492 18284 24544 18290
rect 21272 18226 21324 18232
rect 24412 18244 24492 18272
rect 20456 17610 20484 18226
rect 20548 17814 20576 18226
rect 21456 18216 21508 18222
rect 21456 18158 21508 18164
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 21468 17814 21496 18158
rect 22112 17882 22140 18158
rect 23020 18080 23072 18086
rect 23020 18022 23072 18028
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 20444 17604 20496 17610
rect 20444 17546 20496 17552
rect 20456 17134 20484 17546
rect 20548 17338 20576 17750
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 20536 17332 20588 17338
rect 20536 17274 20588 17280
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20548 17066 20576 17274
rect 20536 17060 20588 17066
rect 20536 17002 20588 17008
rect 20640 16998 20668 17614
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20456 16794 20484 16934
rect 20640 16794 20668 16934
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20824 16522 20852 16934
rect 21008 16794 21036 17478
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20812 16516 20864 16522
rect 20812 16458 20864 16464
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20732 16114 20760 16390
rect 20824 16250 20852 16458
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 19798 15736 19854 15745
rect 19708 15700 19760 15706
rect 19798 15671 19854 15680
rect 19708 15642 19760 15648
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18616 15026 18644 15438
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18984 14822 19012 15438
rect 19536 14890 19564 15574
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19628 14958 19656 15438
rect 19720 14958 19748 15642
rect 19616 14952 19668 14958
rect 19616 14894 19668 14900
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 19064 14816 19116 14822
rect 19260 14770 19288 14826
rect 19116 14764 19288 14770
rect 19064 14758 19288 14764
rect 18984 14618 19012 14758
rect 19076 14742 19288 14758
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 19076 14414 19104 14742
rect 19628 14482 19656 14894
rect 19720 14618 19748 14894
rect 19708 14612 19760 14618
rect 19708 14554 19760 14560
rect 19812 14498 19840 15671
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20364 15094 20392 15438
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19720 14470 19840 14498
rect 20548 14482 20576 15846
rect 20640 15570 20668 16050
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20640 15094 20668 15506
rect 20732 15434 20760 16050
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20824 14618 20852 16050
rect 21008 16046 21036 16730
rect 22112 16658 22140 17614
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21468 16114 21496 16526
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 21008 15484 21036 15982
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21100 15609 21128 15846
rect 21086 15600 21142 15609
rect 21468 15570 21496 16050
rect 22112 15638 22140 16594
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 21086 15535 21142 15544
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21088 15496 21140 15502
rect 21008 15456 21088 15484
rect 21284 15473 21312 15506
rect 22756 15502 22784 16390
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 22744 15496 22796 15502
rect 21088 15438 21140 15444
rect 21270 15464 21326 15473
rect 21100 15366 21128 15438
rect 22744 15438 22796 15444
rect 21270 15399 21326 15408
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 21100 14890 21128 15302
rect 22480 14890 22508 15302
rect 22756 15026 22784 15438
rect 22940 15434 22968 15982
rect 23032 15586 23060 18022
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 23124 16658 23152 17138
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 23204 16584 23256 16590
rect 23204 16526 23256 16532
rect 23216 16250 23244 16526
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 23032 15558 23152 15586
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 22928 15428 22980 15434
rect 22928 15370 22980 15376
rect 22940 15026 22968 15370
rect 23032 15094 23060 15438
rect 23020 15088 23072 15094
rect 23020 15030 23072 15036
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 21088 14884 21140 14890
rect 21088 14826 21140 14832
rect 22468 14884 22520 14890
rect 22468 14826 22520 14832
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20536 14476 20588 14482
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 18420 13456 18472 13462
rect 18420 13398 18472 13404
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18432 12986 18460 13194
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18524 12918 18552 14350
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 18800 12850 18828 13262
rect 18892 12850 18920 13670
rect 19260 13394 19288 13874
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19076 12850 19104 13126
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 18432 12646 18460 12786
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18328 12368 18380 12374
rect 18328 12310 18380 12316
rect 18892 11898 18920 12786
rect 19168 12238 19196 12922
rect 19260 12646 19288 13330
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 17144 10674 17172 11154
rect 18708 11082 18736 11494
rect 19168 11354 19196 12174
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19260 11234 19288 12582
rect 19352 12306 19380 12650
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19444 12238 19472 13398
rect 19720 13326 19748 14470
rect 20536 14418 20588 14424
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19800 13252 19852 13258
rect 19800 13194 19852 13200
rect 19812 12850 19840 13194
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 20088 12442 20116 12786
rect 20732 12714 20760 13126
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19168 11206 19288 11234
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 19168 10810 19196 11206
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19260 10674 19288 11018
rect 19904 10810 19932 12174
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20548 11694 20576 12038
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 20548 11218 20576 11630
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20732 11014 20760 12650
rect 20916 11082 20944 14214
rect 21468 14074 21496 14350
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21468 13462 21496 14010
rect 22388 13938 22416 14350
rect 22480 13938 22508 14826
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22664 14618 22692 14758
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 22664 14278 22692 14554
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22572 14113 22600 14214
rect 22558 14104 22614 14113
rect 22558 14039 22614 14048
rect 22756 13938 22784 14758
rect 23124 14498 23152 15558
rect 23216 15502 23244 16186
rect 23308 16182 23336 17138
rect 23480 16720 23532 16726
rect 23480 16662 23532 16668
rect 23296 16176 23348 16182
rect 23296 16118 23348 16124
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23204 14612 23256 14618
rect 23204 14554 23256 14560
rect 23032 14470 23152 14498
rect 23032 13938 23060 14470
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23124 14074 23152 14350
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21456 13456 21508 13462
rect 21456 13398 21508 13404
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21468 12918 21496 13126
rect 21456 12912 21508 12918
rect 21456 12854 21508 12860
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21192 11762 21220 12582
rect 21468 12306 21496 12854
rect 21560 12850 21588 13466
rect 22388 13258 22416 13874
rect 22376 13252 22428 13258
rect 22376 13194 22428 13200
rect 22388 12986 22416 13194
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 22204 11830 22232 12922
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 19720 9926 19748 10610
rect 20732 10606 20760 10950
rect 21192 10606 21220 11698
rect 22480 11354 22508 13874
rect 23032 13530 23060 13874
rect 23216 13530 23244 14554
rect 23308 14482 23336 14758
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23400 14414 23428 15846
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23308 13326 23336 14282
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23400 14006 23428 14214
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 23492 13938 23520 16662
rect 24044 16590 24072 17138
rect 24032 16584 24084 16590
rect 24032 16526 24084 16532
rect 23572 16448 23624 16454
rect 23756 16448 23808 16454
rect 23572 16390 23624 16396
rect 23754 16416 23756 16425
rect 23848 16448 23900 16454
rect 23808 16416 23810 16425
rect 23584 14482 23612 16390
rect 23848 16390 23900 16396
rect 23754 16351 23810 16360
rect 23860 16182 23888 16390
rect 23848 16176 23900 16182
rect 23848 16118 23900 16124
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23492 13394 23520 13874
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23308 11762 23336 12038
rect 23400 11830 23428 12038
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 23296 11756 23348 11762
rect 23584 11744 23612 14418
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23676 13938 23704 14214
rect 23860 13938 23888 16118
rect 24044 15638 24072 16526
rect 24412 16114 24440 18244
rect 24492 18226 24544 18232
rect 24872 18278 24992 18306
rect 24872 18154 24900 18278
rect 24860 18148 24912 18154
rect 24860 18090 24912 18096
rect 24952 18148 25004 18154
rect 24952 18090 25004 18096
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24780 16250 24808 16594
rect 24584 16244 24636 16250
rect 24584 16186 24636 16192
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 24136 15706 24164 15982
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24032 15632 24084 15638
rect 24032 15574 24084 15580
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23952 14056 23980 15302
rect 24044 15094 24072 15574
rect 24214 15464 24270 15473
rect 24214 15399 24270 15408
rect 24032 15088 24084 15094
rect 24032 15030 24084 15036
rect 23952 14028 24072 14056
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 23952 12986 23980 13874
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 23952 11762 23980 12718
rect 24044 12238 24072 14028
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24136 13394 24164 13874
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24228 12442 24256 15399
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24320 13802 24348 14214
rect 24308 13796 24360 13802
rect 24308 13738 24360 13744
rect 24308 13388 24360 13394
rect 24308 13330 24360 13336
rect 24320 12442 24348 13330
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24308 12436 24360 12442
rect 24308 12378 24360 12384
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24044 12102 24072 12174
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24136 11898 24164 12174
rect 24228 12170 24256 12378
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24216 12164 24268 12170
rect 24216 12106 24268 12112
rect 24124 11892 24176 11898
rect 24044 11852 24124 11880
rect 23664 11756 23716 11762
rect 23584 11716 23664 11744
rect 23296 11698 23348 11704
rect 23664 11698 23716 11704
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 21468 10606 21496 11154
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22020 10742 22048 11086
rect 22664 11014 22692 11698
rect 22940 11626 22968 11698
rect 22928 11620 22980 11626
rect 22928 11562 22980 11568
rect 23296 11620 23348 11626
rect 23296 11562 23348 11568
rect 22940 11218 22968 11562
rect 22928 11212 22980 11218
rect 22928 11154 22980 11160
rect 23308 11082 23336 11562
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23400 11354 23428 11494
rect 23388 11348 23440 11354
rect 23388 11290 23440 11296
rect 24044 11286 24072 11852
rect 24124 11834 24176 11840
rect 24320 11762 24348 12174
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24032 11280 24084 11286
rect 24032 11222 24084 11228
rect 24136 11218 24164 11494
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 24228 11082 24256 11630
rect 24412 11354 24440 13126
rect 24596 12374 24624 16186
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24780 15638 24808 16050
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 24780 14550 24808 15574
rect 24768 14544 24820 14550
rect 24768 14486 24820 14492
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24766 14376 24822 14385
rect 24766 14311 24768 14320
rect 24820 14311 24822 14320
rect 24768 14282 24820 14288
rect 24872 13977 24900 14418
rect 24858 13968 24914 13977
rect 24858 13903 24860 13912
rect 24912 13903 24914 13912
rect 24860 13874 24912 13880
rect 24584 12368 24636 12374
rect 24584 12310 24636 12316
rect 24492 11756 24544 11762
rect 24492 11698 24544 11704
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24504 11150 24532 11698
rect 24596 11694 24624 12310
rect 24964 11830 24992 18090
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25148 15473 25176 15642
rect 25226 15600 25282 15609
rect 25226 15535 25282 15544
rect 25320 15564 25372 15570
rect 25240 15502 25268 15535
rect 25320 15506 25372 15512
rect 25228 15496 25280 15502
rect 25134 15464 25190 15473
rect 25228 15438 25280 15444
rect 25134 15399 25190 15408
rect 25148 14822 25176 15399
rect 25332 15026 25360 15506
rect 25320 15020 25372 15026
rect 25320 14962 25372 14968
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25044 13796 25096 13802
rect 25044 13738 25096 13744
rect 25056 13258 25084 13738
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25056 12306 25084 12922
rect 25228 12844 25280 12850
rect 25228 12786 25280 12792
rect 25240 12306 25268 12786
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 24952 11824 25004 11830
rect 24952 11766 25004 11772
rect 25240 11762 25268 12242
rect 25332 11762 25360 13874
rect 25228 11756 25280 11762
rect 25228 11698 25280 11704
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 24584 11688 24636 11694
rect 24584 11630 24636 11636
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 22652 11008 22704 11014
rect 22652 10950 22704 10956
rect 22008 10736 22060 10742
rect 22008 10678 22060 10684
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21468 10130 21496 10542
rect 22020 10470 22048 10678
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 19720 3942 19748 9862
rect 22020 8838 22048 10406
rect 25424 10266 25452 20198
rect 26620 19854 26648 20334
rect 27908 20262 27936 20402
rect 29564 20398 29592 20878
rect 29552 20392 29604 20398
rect 29552 20334 29604 20340
rect 27896 20256 27948 20262
rect 27896 20198 27948 20204
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 26608 19848 26660 19854
rect 26608 19790 26660 19796
rect 26884 19848 26936 19854
rect 26884 19790 26936 19796
rect 26620 19446 26648 19790
rect 26608 19440 26660 19446
rect 26608 19382 26660 19388
rect 26896 19378 26924 19790
rect 27264 19378 27292 19994
rect 28816 19712 28868 19718
rect 28816 19654 28868 19660
rect 28828 19446 28856 19654
rect 28816 19440 28868 19446
rect 28816 19382 28868 19388
rect 29564 19394 29592 20334
rect 29564 19378 29684 19394
rect 26884 19372 26936 19378
rect 26884 19314 26936 19320
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27528 19372 27580 19378
rect 29564 19372 29696 19378
rect 29564 19366 29644 19372
rect 27528 19314 27580 19320
rect 29644 19314 29696 19320
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25504 18148 25556 18154
rect 25504 18090 25556 18096
rect 25516 16794 25544 18090
rect 25608 17814 25636 18226
rect 25700 18086 25728 18226
rect 25688 18080 25740 18086
rect 25688 18022 25740 18028
rect 25596 17808 25648 17814
rect 25596 17750 25648 17756
rect 25976 17678 26004 18226
rect 26252 17678 26280 19110
rect 26332 18216 26384 18222
rect 26332 18158 26384 18164
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 25964 17672 26016 17678
rect 25964 17614 26016 17620
rect 26240 17672 26292 17678
rect 26240 17614 26292 17620
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 26240 16584 26292 16590
rect 26240 16526 26292 16532
rect 25596 16448 25648 16454
rect 25596 16390 25648 16396
rect 25608 16114 25636 16390
rect 26252 16130 26280 16526
rect 26344 16250 26372 18158
rect 26528 17882 26556 18158
rect 26516 17876 26568 17882
rect 26516 17818 26568 17824
rect 26988 17610 27016 19314
rect 27356 18766 27384 19314
rect 27344 18760 27396 18766
rect 27344 18702 27396 18708
rect 27356 18154 27384 18702
rect 27540 18426 27568 19314
rect 28356 19304 28408 19310
rect 28356 19246 28408 19252
rect 28368 18970 28396 19246
rect 28356 18964 28408 18970
rect 28356 18906 28408 18912
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 28080 18692 28132 18698
rect 28080 18634 28132 18640
rect 28632 18692 28684 18698
rect 28632 18634 28684 18640
rect 29184 18692 29236 18698
rect 29184 18634 29236 18640
rect 27528 18420 27580 18426
rect 27528 18362 27580 18368
rect 27436 18352 27488 18358
rect 27436 18294 27488 18300
rect 27344 18148 27396 18154
rect 27344 18090 27396 18096
rect 27448 17678 27476 18294
rect 28092 18290 28120 18634
rect 28356 18624 28408 18630
rect 28356 18566 28408 18572
rect 28368 18426 28396 18566
rect 28644 18426 28672 18634
rect 28356 18420 28408 18426
rect 28356 18362 28408 18368
rect 28632 18420 28684 18426
rect 28632 18362 28684 18368
rect 27804 18284 27856 18290
rect 27804 18226 27856 18232
rect 28080 18284 28132 18290
rect 28080 18226 28132 18232
rect 28172 18284 28224 18290
rect 28632 18284 28684 18290
rect 28172 18226 28224 18232
rect 28552 18244 28632 18272
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27252 17672 27304 17678
rect 27252 17614 27304 17620
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 26976 17604 27028 17610
rect 26976 17546 27028 17552
rect 26792 16584 26844 16590
rect 26792 16526 26844 16532
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26516 16516 26568 16522
rect 26516 16458 26568 16464
rect 26608 16516 26660 16522
rect 26608 16458 26660 16464
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 25596 16108 25648 16114
rect 25596 16050 25648 16056
rect 25964 16108 26016 16114
rect 26252 16102 26372 16130
rect 25964 16050 26016 16056
rect 25872 15904 25924 15910
rect 25872 15846 25924 15852
rect 25884 15570 25912 15846
rect 25872 15564 25924 15570
rect 25872 15506 25924 15512
rect 25976 15502 26004 16050
rect 26344 15910 26372 16102
rect 26528 16046 26556 16458
rect 26516 16040 26568 16046
rect 26516 15982 26568 15988
rect 26332 15904 26384 15910
rect 26332 15846 26384 15852
rect 26148 15564 26200 15570
rect 26148 15506 26200 15512
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25964 15496 26016 15502
rect 25964 15438 26016 15444
rect 25516 15366 25544 15438
rect 25504 15360 25556 15366
rect 25504 15302 25556 15308
rect 25516 15026 25544 15302
rect 25504 15020 25556 15026
rect 25504 14962 25556 14968
rect 25516 14074 25544 14962
rect 25976 14890 26004 15438
rect 25596 14884 25648 14890
rect 25596 14826 25648 14832
rect 25964 14884 26016 14890
rect 25964 14826 26016 14832
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25608 13938 25636 14826
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25516 12986 25544 13874
rect 25608 13841 25636 13874
rect 25976 13870 26004 14826
rect 26160 13938 26188 15506
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 26148 13932 26200 13938
rect 26148 13874 26200 13880
rect 25964 13864 26016 13870
rect 25594 13832 25650 13841
rect 25964 13806 26016 13812
rect 25594 13767 25650 13776
rect 25688 13796 25740 13802
rect 25688 13738 25740 13744
rect 25504 12980 25556 12986
rect 25504 12922 25556 12928
rect 25700 12850 25728 13738
rect 25976 13462 26004 13806
rect 26160 13462 26188 13874
rect 25964 13456 26016 13462
rect 25964 13398 26016 13404
rect 26148 13456 26200 13462
rect 26148 13398 26200 13404
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 25792 12442 25820 12786
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 26160 12374 26188 13398
rect 26148 12368 26200 12374
rect 26068 12316 26148 12322
rect 26068 12310 26200 12316
rect 26068 12294 26188 12310
rect 25780 12232 25832 12238
rect 25780 12174 25832 12180
rect 25792 10674 25820 12174
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25884 11830 25912 12038
rect 25872 11824 25924 11830
rect 25872 11766 25924 11772
rect 26068 11694 26096 12294
rect 26252 12238 26280 14214
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 25872 11688 25924 11694
rect 25872 11630 25924 11636
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 25884 11558 25912 11630
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 26068 11014 26096 11630
rect 26160 11354 26188 12174
rect 26240 11824 26292 11830
rect 26240 11766 26292 11772
rect 26148 11348 26200 11354
rect 26148 11290 26200 11296
rect 26252 11150 26280 11766
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26056 11008 26108 11014
rect 26056 10950 26108 10956
rect 26344 10674 26372 15846
rect 26424 15496 26476 15502
rect 26424 15438 26476 15444
rect 26436 15162 26464 15438
rect 26424 15156 26476 15162
rect 26424 15098 26476 15104
rect 26424 13864 26476 13870
rect 26422 13832 26424 13841
rect 26476 13832 26478 13841
rect 26422 13767 26478 13776
rect 26620 13734 26648 16458
rect 26698 16416 26754 16425
rect 26698 16351 26754 16360
rect 26608 13728 26660 13734
rect 26608 13670 26660 13676
rect 26712 13394 26740 16351
rect 26804 16182 26832 16526
rect 26792 16176 26844 16182
rect 26792 16118 26844 16124
rect 26896 14414 26924 16526
rect 26988 15366 27016 17546
rect 27264 17542 27292 17614
rect 27252 17536 27304 17542
rect 27252 17478 27304 17484
rect 27264 16250 27292 17478
rect 27448 17134 27476 17614
rect 27436 17128 27488 17134
rect 27436 17070 27488 17076
rect 27344 16516 27396 16522
rect 27344 16458 27396 16464
rect 27356 16425 27384 16458
rect 27342 16416 27398 16425
rect 27342 16351 27398 16360
rect 27252 16244 27304 16250
rect 27252 16186 27304 16192
rect 27344 16176 27396 16182
rect 27448 16130 27476 17070
rect 27528 16448 27580 16454
rect 27528 16390 27580 16396
rect 27540 16250 27568 16390
rect 27528 16244 27580 16250
rect 27528 16186 27580 16192
rect 27396 16124 27476 16130
rect 27344 16118 27476 16124
rect 27160 16108 27212 16114
rect 27356 16102 27476 16118
rect 27160 16050 27212 16056
rect 27068 15428 27120 15434
rect 27068 15370 27120 15376
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 27080 15026 27108 15370
rect 27172 15026 27200 16050
rect 27252 15972 27304 15978
rect 27252 15914 27304 15920
rect 27264 15502 27292 15914
rect 27448 15570 27476 16102
rect 27436 15564 27488 15570
rect 27436 15506 27488 15512
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27540 15434 27568 16186
rect 27528 15428 27580 15434
rect 27528 15370 27580 15376
rect 26976 15020 27028 15026
rect 26976 14962 27028 14968
rect 27068 15020 27120 15026
rect 27068 14962 27120 14968
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 26884 14408 26936 14414
rect 26884 14350 26936 14356
rect 26988 14346 27016 14962
rect 27172 14482 27200 14962
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27344 14408 27396 14414
rect 27528 14408 27580 14414
rect 27344 14350 27396 14356
rect 27526 14376 27528 14385
rect 27580 14376 27582 14385
rect 26976 14340 27028 14346
rect 26976 14282 27028 14288
rect 26792 13728 26844 13734
rect 26792 13670 26844 13676
rect 26804 13394 26832 13670
rect 26700 13388 26752 13394
rect 26700 13330 26752 13336
rect 26792 13388 26844 13394
rect 26792 13330 26844 13336
rect 26712 12918 26740 13330
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26700 12912 26752 12918
rect 26700 12854 26752 12860
rect 26712 12306 26740 12854
rect 26700 12300 26752 12306
rect 26700 12242 26752 12248
rect 26608 12096 26660 12102
rect 26608 12038 26660 12044
rect 26516 11688 26568 11694
rect 26516 11630 26568 11636
rect 26424 11552 26476 11558
rect 26424 11494 26476 11500
rect 26436 11150 26464 11494
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 26528 11082 26556 11630
rect 26620 11150 26648 12038
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26516 11076 26568 11082
rect 26516 11018 26568 11024
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 26332 10668 26384 10674
rect 26332 10610 26384 10616
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 25412 10260 25464 10266
rect 25412 10202 25464 10208
rect 25424 10062 25452 10202
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 26528 9586 26556 10066
rect 26620 10062 26648 10406
rect 26804 10062 26832 13126
rect 26988 12714 27016 14282
rect 27356 13977 27384 14350
rect 27526 14311 27582 14320
rect 27632 14226 27660 18158
rect 27712 17604 27764 17610
rect 27712 17546 27764 17552
rect 27724 16998 27752 17546
rect 27816 17202 27844 18226
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27712 16992 27764 16998
rect 27712 16934 27764 16940
rect 27816 16522 27844 17138
rect 28184 17066 28212 18226
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28276 17678 28304 18022
rect 28552 17746 28580 18244
rect 28632 18226 28684 18232
rect 28540 17740 28592 17746
rect 28540 17682 28592 17688
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28368 17270 28396 17614
rect 28356 17264 28408 17270
rect 28356 17206 28408 17212
rect 28264 17196 28316 17202
rect 28264 17138 28316 17144
rect 28172 17060 28224 17066
rect 28172 17002 28224 17008
rect 28184 16794 28212 17002
rect 28276 16794 28304 17138
rect 28172 16788 28224 16794
rect 28172 16730 28224 16736
rect 28264 16788 28316 16794
rect 28264 16730 28316 16736
rect 28368 16726 28396 17206
rect 28552 17202 28580 17682
rect 28908 17604 28960 17610
rect 28908 17546 28960 17552
rect 28816 17264 28868 17270
rect 28816 17206 28868 17212
rect 28540 17196 28592 17202
rect 28540 17138 28592 17144
rect 28552 16794 28580 17138
rect 28828 17066 28856 17206
rect 28920 17202 28948 17546
rect 29196 17338 29224 18634
rect 29276 18624 29328 18630
rect 29276 18566 29328 18572
rect 29288 18358 29316 18566
rect 29276 18352 29328 18358
rect 29276 18294 29328 18300
rect 29460 18216 29512 18222
rect 29458 18184 29460 18193
rect 29512 18184 29514 18193
rect 29458 18119 29514 18128
rect 29184 17332 29236 17338
rect 29184 17274 29236 17280
rect 28908 17196 28960 17202
rect 28908 17138 28960 17144
rect 29104 17190 29316 17218
rect 28816 17060 28868 17066
rect 28816 17002 28868 17008
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 28540 16788 28592 16794
rect 28540 16730 28592 16736
rect 28356 16720 28408 16726
rect 28356 16662 28408 16668
rect 28552 16590 28580 16730
rect 28540 16584 28592 16590
rect 28540 16526 28592 16532
rect 27804 16516 27856 16522
rect 27804 16458 27856 16464
rect 27712 15972 27764 15978
rect 27712 15914 27764 15920
rect 27724 15745 27752 15914
rect 27710 15736 27766 15745
rect 27816 15706 27844 16458
rect 27896 16448 27948 16454
rect 27896 16390 27948 16396
rect 27710 15671 27766 15680
rect 27804 15700 27856 15706
rect 27724 15502 27752 15671
rect 27804 15642 27856 15648
rect 27712 15496 27764 15502
rect 27712 15438 27764 15444
rect 27712 15020 27764 15026
rect 27712 14962 27764 14968
rect 27724 14550 27752 14962
rect 27804 14816 27856 14822
rect 27804 14758 27856 14764
rect 27712 14544 27764 14550
rect 27712 14486 27764 14492
rect 27540 14198 27660 14226
rect 27540 14006 27568 14198
rect 27618 14104 27674 14113
rect 27618 14039 27674 14048
rect 27528 14000 27580 14006
rect 27342 13968 27398 13977
rect 27528 13942 27580 13948
rect 27342 13903 27344 13912
rect 27396 13903 27398 13912
rect 27436 13932 27488 13938
rect 27344 13874 27396 13880
rect 27436 13874 27488 13880
rect 27068 13864 27120 13870
rect 27068 13806 27120 13812
rect 26976 12708 27028 12714
rect 26976 12650 27028 12656
rect 27080 12102 27108 13806
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 27172 13394 27200 13670
rect 27448 13530 27476 13874
rect 27540 13546 27568 13942
rect 27632 13734 27660 14039
rect 27816 13938 27844 14758
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27620 13728 27672 13734
rect 27620 13670 27672 13676
rect 27436 13524 27488 13530
rect 27540 13518 27660 13546
rect 27436 13466 27488 13472
rect 27160 13388 27212 13394
rect 27160 13330 27212 13336
rect 27528 13388 27580 13394
rect 27528 13330 27580 13336
rect 27344 12640 27396 12646
rect 27344 12582 27396 12588
rect 27068 12096 27120 12102
rect 27068 12038 27120 12044
rect 27252 11552 27304 11558
rect 27252 11494 27304 11500
rect 27264 11082 27292 11494
rect 27356 11150 27384 12582
rect 27540 11762 27568 13330
rect 27632 12186 27660 13518
rect 27724 13326 27752 13874
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27724 12374 27752 13262
rect 27908 13258 27936 16390
rect 27988 16108 28040 16114
rect 27988 16050 28040 16056
rect 28000 15638 28028 16050
rect 27988 15632 28040 15638
rect 27988 15574 28040 15580
rect 28356 15020 28408 15026
rect 28356 14962 28408 14968
rect 28170 14920 28226 14929
rect 28170 14855 28226 14864
rect 28184 14618 28212 14855
rect 28172 14612 28224 14618
rect 28172 14554 28224 14560
rect 28184 14498 28212 14554
rect 28092 14482 28212 14498
rect 28080 14476 28212 14482
rect 28132 14470 28212 14476
rect 28080 14418 28132 14424
rect 28080 14272 28132 14278
rect 28080 14214 28132 14220
rect 28092 13938 28120 14214
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 28368 13394 28396 14962
rect 28552 14362 28580 16526
rect 28644 15026 28672 16934
rect 28828 15586 28856 17002
rect 28920 16726 28948 17138
rect 29104 17066 29132 17190
rect 29288 17184 29316 17190
rect 29368 17196 29420 17202
rect 29288 17156 29368 17184
rect 29368 17138 29420 17144
rect 29184 17128 29236 17134
rect 29184 17070 29236 17076
rect 29092 17060 29144 17066
rect 29092 17002 29144 17008
rect 29196 16998 29224 17070
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 28908 16720 28960 16726
rect 28908 16662 28960 16668
rect 29184 16176 29236 16182
rect 29184 16118 29236 16124
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29012 15706 29040 16050
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 28828 15558 28948 15586
rect 28816 15496 28868 15502
rect 28816 15438 28868 15444
rect 28632 15020 28684 15026
rect 28632 14962 28684 14968
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 28736 14822 28764 14962
rect 28724 14816 28776 14822
rect 28724 14758 28776 14764
rect 28630 14376 28686 14385
rect 28552 14334 28630 14362
rect 28630 14311 28686 14320
rect 28356 13388 28408 13394
rect 28356 13330 28408 13336
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 27896 13252 27948 13258
rect 27896 13194 27948 13200
rect 28356 13252 28408 13258
rect 28356 13194 28408 13200
rect 27712 12368 27764 12374
rect 27712 12310 27764 12316
rect 27712 12232 27764 12238
rect 27632 12180 27712 12186
rect 27632 12174 27764 12180
rect 27632 12158 27752 12174
rect 27724 11762 27752 12158
rect 27528 11756 27580 11762
rect 27528 11698 27580 11704
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 27712 11756 27764 11762
rect 27712 11698 27764 11704
rect 27632 11218 27660 11698
rect 27816 11354 27844 13194
rect 27908 12986 27936 13194
rect 27896 12980 27948 12986
rect 27896 12922 27948 12928
rect 27896 12708 27948 12714
rect 27896 12650 27948 12656
rect 27908 12238 27936 12650
rect 28368 12434 28396 13194
rect 28540 12980 28592 12986
rect 28540 12922 28592 12928
rect 28552 12442 28580 12922
rect 28276 12406 28396 12434
rect 28540 12436 28592 12442
rect 28276 12238 28304 12406
rect 28540 12378 28592 12384
rect 27896 12232 27948 12238
rect 27896 12174 27948 12180
rect 27988 12232 28040 12238
rect 27988 12174 28040 12180
rect 28264 12232 28316 12238
rect 28264 12174 28316 12180
rect 27896 12096 27948 12102
rect 27896 12038 27948 12044
rect 27804 11348 27856 11354
rect 27804 11290 27856 11296
rect 27908 11218 27936 12038
rect 28000 11830 28028 12174
rect 28172 12164 28224 12170
rect 28172 12106 28224 12112
rect 27988 11824 28040 11830
rect 27988 11766 28040 11772
rect 27620 11212 27672 11218
rect 27620 11154 27672 11160
rect 27896 11212 27948 11218
rect 27896 11154 27948 11160
rect 28184 11150 28212 12106
rect 28276 11626 28304 12174
rect 28264 11620 28316 11626
rect 28264 11562 28316 11568
rect 27344 11144 27396 11150
rect 27344 11086 27396 11092
rect 28172 11144 28224 11150
rect 28552 11098 28580 12378
rect 28644 12306 28672 14311
rect 28736 13326 28764 14758
rect 28828 14074 28856 15438
rect 28920 15162 28948 15558
rect 28908 15156 28960 15162
rect 28908 15098 28960 15104
rect 29196 15026 29224 16118
rect 29564 16114 29592 18702
rect 29748 17882 29776 21490
rect 29826 20496 29882 20505
rect 29826 20431 29882 20440
rect 29840 19310 29868 20431
rect 30116 20058 30144 21558
rect 30208 20890 30236 22102
rect 30300 22030 30328 23122
rect 30668 23118 30696 24262
rect 30852 23798 30880 24890
rect 30944 24818 30972 25162
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30944 24682 30972 24754
rect 31128 24750 31156 26522
rect 31404 26042 31432 27066
rect 31680 26586 31708 27474
rect 32048 26926 32076 27950
rect 33244 27674 33272 27950
rect 34520 27872 34572 27878
rect 34520 27814 34572 27820
rect 33232 27668 33284 27674
rect 33232 27610 33284 27616
rect 34428 27600 34480 27606
rect 34428 27542 34480 27548
rect 34060 27464 34112 27470
rect 34060 27406 34112 27412
rect 34152 27464 34204 27470
rect 34152 27406 34204 27412
rect 32588 27396 32640 27402
rect 32588 27338 32640 27344
rect 32036 26920 32088 26926
rect 32036 26862 32088 26868
rect 32496 26920 32548 26926
rect 32496 26862 32548 26868
rect 31668 26580 31720 26586
rect 31668 26522 31720 26528
rect 31576 26376 31628 26382
rect 31576 26318 31628 26324
rect 31392 26036 31444 26042
rect 31392 25978 31444 25984
rect 31588 25974 31616 26318
rect 31576 25968 31628 25974
rect 31576 25910 31628 25916
rect 31392 25832 31444 25838
rect 31392 25774 31444 25780
rect 31300 25356 31352 25362
rect 31300 25298 31352 25304
rect 31116 24744 31168 24750
rect 31116 24686 31168 24692
rect 30932 24676 30984 24682
rect 30932 24618 30984 24624
rect 30944 23866 30972 24618
rect 30932 23860 30984 23866
rect 30932 23802 30984 23808
rect 30840 23792 30892 23798
rect 30840 23734 30892 23740
rect 30852 23662 30880 23734
rect 30840 23656 30892 23662
rect 30840 23598 30892 23604
rect 30656 23112 30708 23118
rect 30656 23054 30708 23060
rect 30380 23044 30432 23050
rect 30380 22986 30432 22992
rect 30392 22642 30420 22986
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30484 22166 30512 22714
rect 30668 22642 30696 23054
rect 30852 22778 30880 23598
rect 31024 23520 31076 23526
rect 31128 23474 31156 24686
rect 31312 24206 31340 25298
rect 31404 25294 31432 25774
rect 31392 25288 31444 25294
rect 31392 25230 31444 25236
rect 31404 24274 31432 25230
rect 31392 24268 31444 24274
rect 31392 24210 31444 24216
rect 31300 24200 31352 24206
rect 31076 23468 31156 23474
rect 31024 23462 31156 23468
rect 31036 23446 31156 23462
rect 31128 23322 31156 23446
rect 31220 24160 31300 24188
rect 31116 23316 31168 23322
rect 31116 23258 31168 23264
rect 31220 23186 31248 24160
rect 31300 24142 31352 24148
rect 31300 24064 31352 24070
rect 31300 24006 31352 24012
rect 31312 23730 31340 24006
rect 31300 23724 31352 23730
rect 31300 23666 31352 23672
rect 31208 23180 31260 23186
rect 31208 23122 31260 23128
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30656 22636 30708 22642
rect 30656 22578 30708 22584
rect 30472 22160 30524 22166
rect 30472 22102 30524 22108
rect 30564 22160 30616 22166
rect 30564 22102 30616 22108
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 30576 21554 30604 22102
rect 30668 21962 30696 22578
rect 31116 22432 31168 22438
rect 31116 22374 31168 22380
rect 31128 22234 31156 22374
rect 31116 22228 31168 22234
rect 31116 22170 31168 22176
rect 31128 22094 31156 22170
rect 31220 22166 31248 23122
rect 31312 23118 31340 23666
rect 31404 23254 31432 24210
rect 31588 24206 31616 25910
rect 31576 24200 31628 24206
rect 31576 24142 31628 24148
rect 31392 23248 31444 23254
rect 31392 23190 31444 23196
rect 31300 23112 31352 23118
rect 31300 23054 31352 23060
rect 31588 22982 31616 24142
rect 32048 23644 32076 26862
rect 32508 26586 32536 26862
rect 32496 26580 32548 26586
rect 32496 26522 32548 26528
rect 32600 26382 32628 27338
rect 33968 26784 34020 26790
rect 33968 26726 34020 26732
rect 32128 26376 32180 26382
rect 32128 26318 32180 26324
rect 32404 26376 32456 26382
rect 32404 26318 32456 26324
rect 32588 26376 32640 26382
rect 32588 26318 32640 26324
rect 32140 25294 32168 26318
rect 32416 26042 32444 26318
rect 32404 26036 32456 26042
rect 32404 25978 32456 25984
rect 32588 25900 32640 25906
rect 32588 25842 32640 25848
rect 32600 25401 32628 25842
rect 32586 25392 32642 25401
rect 32586 25327 32588 25336
rect 32640 25327 32642 25336
rect 32588 25298 32640 25304
rect 33980 25294 34008 26726
rect 34072 25906 34100 27406
rect 34164 26586 34192 27406
rect 34152 26580 34204 26586
rect 34152 26522 34204 26528
rect 34060 25900 34112 25906
rect 34060 25842 34112 25848
rect 34072 25294 34100 25842
rect 34244 25832 34296 25838
rect 34244 25774 34296 25780
rect 32128 25288 32180 25294
rect 32128 25230 32180 25236
rect 33968 25288 34020 25294
rect 33968 25230 34020 25236
rect 34060 25288 34112 25294
rect 34060 25230 34112 25236
rect 33784 25152 33836 25158
rect 33784 25094 33836 25100
rect 33796 24818 33824 25094
rect 33784 24812 33836 24818
rect 33784 24754 33836 24760
rect 33416 24744 33468 24750
rect 33416 24686 33468 24692
rect 33428 24138 33456 24686
rect 32772 24132 32824 24138
rect 32772 24074 32824 24080
rect 33416 24132 33468 24138
rect 33416 24074 33468 24080
rect 32784 23662 32812 24074
rect 32128 23656 32180 23662
rect 32048 23616 32128 23644
rect 32128 23598 32180 23604
rect 32772 23656 32824 23662
rect 32772 23598 32824 23604
rect 33140 23656 33192 23662
rect 33140 23598 33192 23604
rect 33324 23656 33376 23662
rect 33324 23598 33376 23604
rect 31852 23112 31904 23118
rect 31758 23080 31814 23089
rect 31852 23054 31904 23060
rect 31758 23015 31760 23024
rect 31812 23015 31814 23024
rect 31760 22986 31812 22992
rect 31576 22976 31628 22982
rect 31576 22918 31628 22924
rect 31864 22642 31892 23054
rect 32036 22772 32088 22778
rect 32036 22714 32088 22720
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 32048 22574 32076 22714
rect 32036 22568 32088 22574
rect 32036 22510 32088 22516
rect 31208 22160 31260 22166
rect 31208 22102 31260 22108
rect 31036 22066 31156 22094
rect 30656 21956 30708 21962
rect 30656 21898 30708 21904
rect 30748 21956 30800 21962
rect 30748 21898 30800 21904
rect 30668 21554 30696 21898
rect 30564 21548 30616 21554
rect 30564 21490 30616 21496
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 30472 21480 30524 21486
rect 30472 21422 30524 21428
rect 30484 21010 30512 21422
rect 30472 21004 30524 21010
rect 30472 20946 30524 20952
rect 30208 20874 30328 20890
rect 30208 20868 30340 20874
rect 30208 20862 30288 20868
rect 30288 20810 30340 20816
rect 30104 20052 30156 20058
rect 30104 19994 30156 20000
rect 30300 19786 30328 20810
rect 30288 19780 30340 19786
rect 30288 19722 30340 19728
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29840 18970 29868 19246
rect 29828 18964 29880 18970
rect 29828 18906 29880 18912
rect 30288 18624 30340 18630
rect 30288 18566 30340 18572
rect 29736 17876 29788 17882
rect 29736 17818 29788 17824
rect 29828 17536 29880 17542
rect 29828 17478 29880 17484
rect 29736 17332 29788 17338
rect 29736 17274 29788 17280
rect 29748 17134 29776 17274
rect 29840 17202 29868 17478
rect 30196 17264 30248 17270
rect 30194 17232 30196 17241
rect 30248 17232 30250 17241
rect 29828 17196 29880 17202
rect 29828 17138 29880 17144
rect 30012 17196 30064 17202
rect 30194 17167 30250 17176
rect 30012 17138 30064 17144
rect 29736 17128 29788 17134
rect 29736 17070 29788 17076
rect 29748 16794 29776 17070
rect 29736 16788 29788 16794
rect 29736 16730 29788 16736
rect 29552 16108 29604 16114
rect 29552 16050 29604 16056
rect 30024 15978 30052 17138
rect 30012 15972 30064 15978
rect 30012 15914 30064 15920
rect 29552 15904 29604 15910
rect 29552 15846 29604 15852
rect 29564 15502 29592 15846
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29184 15020 29236 15026
rect 29184 14962 29236 14968
rect 28816 14068 28868 14074
rect 28816 14010 28868 14016
rect 29196 13530 29224 14962
rect 29460 14476 29512 14482
rect 29460 14418 29512 14424
rect 29472 13870 29500 14418
rect 29564 14414 29592 15438
rect 29748 14482 29776 15438
rect 30012 14884 30064 14890
rect 30012 14826 30064 14832
rect 29736 14476 29788 14482
rect 29736 14418 29788 14424
rect 29552 14408 29604 14414
rect 29552 14350 29604 14356
rect 29460 13864 29512 13870
rect 29460 13806 29512 13812
rect 29184 13524 29236 13530
rect 29184 13466 29236 13472
rect 28724 13320 28776 13326
rect 28724 13262 28776 13268
rect 28632 12300 28684 12306
rect 28632 12242 28684 12248
rect 29472 12238 29500 13806
rect 29460 12232 29512 12238
rect 29460 12174 29512 12180
rect 29472 11762 29500 12174
rect 29460 11756 29512 11762
rect 29460 11698 29512 11704
rect 29460 11212 29512 11218
rect 29460 11154 29512 11160
rect 28172 11086 28224 11092
rect 28460 11082 28580 11098
rect 27252 11076 27304 11082
rect 27252 11018 27304 11024
rect 28448 11076 28580 11082
rect 28500 11070 28580 11076
rect 28448 11018 28500 11024
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 28632 11008 28684 11014
rect 28632 10950 28684 10956
rect 26976 10736 27028 10742
rect 26976 10678 27028 10684
rect 26988 10062 27016 10678
rect 28184 10606 28212 10950
rect 28644 10674 28672 10950
rect 29472 10674 29500 11154
rect 29564 10674 29592 14350
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29840 13530 29868 13806
rect 29828 13524 29880 13530
rect 29828 13466 29880 13472
rect 29828 12096 29880 12102
rect 29828 12038 29880 12044
rect 29736 11688 29788 11694
rect 29736 11630 29788 11636
rect 29748 11354 29776 11630
rect 29840 11354 29868 12038
rect 29736 11348 29788 11354
rect 29736 11290 29788 11296
rect 29828 11348 29880 11354
rect 29828 11290 29880 11296
rect 28632 10668 28684 10674
rect 28632 10610 28684 10616
rect 29460 10668 29512 10674
rect 29460 10610 29512 10616
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 28172 10600 28224 10606
rect 28172 10542 28224 10548
rect 29828 10600 29880 10606
rect 29828 10542 29880 10548
rect 28448 10464 28500 10470
rect 28448 10406 28500 10412
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 26792 10056 26844 10062
rect 26792 9998 26844 10004
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26884 9988 26936 9994
rect 26884 9930 26936 9936
rect 26896 9722 26924 9930
rect 27160 9920 27212 9926
rect 27160 9862 27212 9868
rect 26884 9716 26936 9722
rect 26884 9658 26936 9664
rect 26516 9580 26568 9586
rect 26516 9522 26568 9528
rect 26528 9042 26556 9522
rect 27172 9042 27200 9862
rect 28460 9654 28488 10406
rect 28448 9648 28500 9654
rect 28448 9590 28500 9596
rect 28816 9648 28868 9654
rect 28816 9590 28868 9596
rect 28828 9518 28856 9590
rect 27988 9512 28040 9518
rect 27986 9480 27988 9489
rect 28816 9512 28868 9518
rect 28040 9480 28042 9489
rect 27986 9415 28042 9424
rect 28262 9480 28318 9489
rect 28816 9454 28868 9460
rect 28262 9415 28318 9424
rect 28276 9178 28304 9415
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 27160 9036 27212 9042
rect 27160 8978 27212 8984
rect 28828 8838 28856 9454
rect 29840 9382 29868 10542
rect 29828 9376 29880 9382
rect 29828 9318 29880 9324
rect 29840 8945 29868 9318
rect 29826 8936 29882 8945
rect 29826 8871 29882 8880
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 28816 8832 28868 8838
rect 28816 8774 28868 8780
rect 29460 8560 29512 8566
rect 29460 8502 29512 8508
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 29196 8090 29224 8366
rect 29184 8084 29236 8090
rect 29184 8026 29236 8032
rect 29472 6866 29500 8502
rect 29460 6860 29512 6866
rect 29460 6802 29512 6808
rect 29472 6254 29500 6802
rect 29460 6248 29512 6254
rect 29460 6190 29512 6196
rect 29472 5778 29500 6190
rect 29460 5772 29512 5778
rect 29460 5714 29512 5720
rect 30024 4826 30052 14826
rect 30300 13258 30328 18566
rect 30760 18426 30788 21898
rect 31036 21554 31064 22066
rect 32140 22030 32168 23598
rect 32956 23520 33008 23526
rect 32956 23462 33008 23468
rect 32588 23316 32640 23322
rect 32588 23258 32640 23264
rect 32600 23186 32628 23258
rect 32864 23248 32916 23254
rect 32864 23190 32916 23196
rect 32588 23180 32640 23186
rect 32588 23122 32640 23128
rect 32312 23112 32364 23118
rect 32312 23054 32364 23060
rect 32324 22642 32352 23054
rect 32312 22636 32364 22642
rect 32312 22578 32364 22584
rect 32600 22438 32628 23122
rect 32680 22772 32732 22778
rect 32680 22714 32732 22720
rect 32692 22642 32720 22714
rect 32876 22710 32904 23190
rect 32864 22704 32916 22710
rect 32864 22646 32916 22652
rect 32968 22642 32996 23462
rect 33152 23322 33180 23598
rect 33140 23316 33192 23322
rect 33140 23258 33192 23264
rect 33232 23044 33284 23050
rect 33232 22986 33284 22992
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32956 22636 33008 22642
rect 32956 22578 33008 22584
rect 33048 22636 33100 22642
rect 33048 22578 33100 22584
rect 32692 22438 32720 22578
rect 32404 22432 32456 22438
rect 32404 22374 32456 22380
rect 32588 22432 32640 22438
rect 32588 22374 32640 22380
rect 32680 22432 32732 22438
rect 32680 22374 32732 22380
rect 32416 22098 32444 22374
rect 32404 22092 32456 22098
rect 32404 22034 32456 22040
rect 31116 22024 31168 22030
rect 31116 21966 31168 21972
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 31128 21690 31156 21966
rect 31944 21956 31996 21962
rect 31944 21898 31996 21904
rect 31116 21684 31168 21690
rect 31116 21626 31168 21632
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 30748 18284 30800 18290
rect 30748 18226 30800 18232
rect 30760 18086 30788 18226
rect 30656 18080 30708 18086
rect 30656 18022 30708 18028
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30668 17746 30696 18022
rect 30760 17882 30788 18022
rect 30748 17876 30800 17882
rect 30748 17818 30800 17824
rect 30656 17740 30708 17746
rect 30656 17682 30708 17688
rect 30668 17202 30696 17682
rect 30748 17536 30800 17542
rect 30748 17478 30800 17484
rect 30760 17338 30788 17478
rect 30748 17332 30800 17338
rect 30748 17274 30800 17280
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30668 14618 30696 17138
rect 30656 14612 30708 14618
rect 30656 14554 30708 14560
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30392 13326 30420 14214
rect 30380 13320 30432 13326
rect 30380 13262 30432 13268
rect 30288 13252 30340 13258
rect 30288 13194 30340 13200
rect 30300 11218 30328 13194
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 30104 10260 30156 10266
rect 30104 10202 30156 10208
rect 30116 6458 30144 10202
rect 30380 8288 30432 8294
rect 30380 8230 30432 8236
rect 30392 7886 30420 8230
rect 30380 7880 30432 7886
rect 30380 7822 30432 7828
rect 30564 7880 30616 7886
rect 30564 7822 30616 7828
rect 30576 7342 30604 7822
rect 30564 7336 30616 7342
rect 30564 7278 30616 7284
rect 30748 7200 30800 7206
rect 30748 7142 30800 7148
rect 30760 7002 30788 7142
rect 30748 6996 30800 7002
rect 30748 6938 30800 6944
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 30288 5772 30340 5778
rect 30288 5714 30340 5720
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 30024 4622 30052 4762
rect 30300 4690 30328 5714
rect 30656 5636 30708 5642
rect 30656 5578 30708 5584
rect 30668 5370 30696 5578
rect 30656 5364 30708 5370
rect 30656 5306 30708 5312
rect 30288 4684 30340 4690
rect 30288 4626 30340 4632
rect 30012 4616 30064 4622
rect 30300 4570 30328 4626
rect 30012 4558 30064 4564
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 30024 3738 30052 4558
rect 30208 4542 30328 4570
rect 30012 3732 30064 3738
rect 30012 3674 30064 3680
rect 30208 3602 30236 4542
rect 30852 4146 30880 21286
rect 31036 20754 31064 21490
rect 31404 21350 31432 21490
rect 31392 21344 31444 21350
rect 31392 21286 31444 21292
rect 31956 21146 31984 21898
rect 32140 21554 32168 21966
rect 32128 21548 32180 21554
rect 32128 21490 32180 21496
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 31116 20800 31168 20806
rect 31036 20748 31116 20754
rect 31036 20742 31168 20748
rect 31036 20726 31156 20742
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 30944 19446 30972 19654
rect 30932 19440 30984 19446
rect 30932 19382 30984 19388
rect 30944 17678 30972 19382
rect 31036 17814 31064 20726
rect 32140 20466 32168 21490
rect 32128 20460 32180 20466
rect 32128 20402 32180 20408
rect 32404 20392 32456 20398
rect 32404 20334 32456 20340
rect 31760 20324 31812 20330
rect 31760 20266 31812 20272
rect 31772 20058 31800 20266
rect 32416 20058 32444 20334
rect 31760 20052 31812 20058
rect 31760 19994 31812 20000
rect 32404 20052 32456 20058
rect 32404 19994 32456 20000
rect 31116 19304 31168 19310
rect 31772 19281 31800 19994
rect 32968 19378 32996 22578
rect 33060 22506 33088 22578
rect 33048 22500 33100 22506
rect 33048 22442 33100 22448
rect 32956 19372 33008 19378
rect 32784 19320 32956 19334
rect 32784 19314 33008 19320
rect 32680 19304 32732 19310
rect 31116 19246 31168 19252
rect 31758 19272 31814 19281
rect 31128 18970 31156 19246
rect 32680 19246 32732 19252
rect 32784 19306 32996 19314
rect 31758 19207 31814 19216
rect 32128 19168 32180 19174
rect 32128 19110 32180 19116
rect 31116 18964 31168 18970
rect 31116 18906 31168 18912
rect 32140 18766 32168 19110
rect 32404 18964 32456 18970
rect 32404 18906 32456 18912
rect 32128 18760 32180 18766
rect 32128 18702 32180 18708
rect 32036 18692 32088 18698
rect 32036 18634 32088 18640
rect 32048 18290 32076 18634
rect 32220 18352 32272 18358
rect 32220 18294 32272 18300
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 31392 17876 31444 17882
rect 31392 17818 31444 17824
rect 31024 17808 31076 17814
rect 31024 17750 31076 17756
rect 31116 17740 31168 17746
rect 31168 17700 31248 17728
rect 31116 17682 31168 17688
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 31024 17604 31076 17610
rect 31024 17546 31076 17552
rect 31116 17604 31168 17610
rect 31116 17546 31168 17552
rect 31036 17338 31064 17546
rect 31024 17332 31076 17338
rect 31024 17274 31076 17280
rect 31024 17128 31076 17134
rect 31024 17070 31076 17076
rect 30932 14408 30984 14414
rect 30932 14350 30984 14356
rect 30944 13802 30972 14350
rect 30932 13796 30984 13802
rect 30932 13738 30984 13744
rect 31036 12646 31064 17070
rect 31128 15502 31156 17546
rect 31220 16590 31248 17700
rect 31404 17649 31432 17818
rect 31390 17640 31446 17649
rect 31390 17575 31446 17584
rect 31208 16584 31260 16590
rect 31208 16526 31260 16532
rect 31116 15496 31168 15502
rect 31116 15438 31168 15444
rect 31128 14498 31156 15438
rect 31128 14470 31248 14498
rect 31220 14006 31248 14470
rect 31208 14000 31260 14006
rect 31208 13942 31260 13948
rect 31024 12640 31076 12646
rect 31024 12582 31076 12588
rect 31404 11694 31432 17575
rect 32048 17338 32076 18226
rect 32128 18080 32180 18086
rect 32128 18022 32180 18028
rect 32140 17746 32168 18022
rect 32128 17740 32180 17746
rect 32128 17682 32180 17688
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 31758 17096 31814 17105
rect 31758 17031 31814 17040
rect 31772 16998 31800 17031
rect 31760 16992 31812 16998
rect 31760 16934 31812 16940
rect 31576 16584 31628 16590
rect 31576 16526 31628 16532
rect 31588 15434 31616 16526
rect 31852 16516 31904 16522
rect 31852 16458 31904 16464
rect 31864 16250 31892 16458
rect 31852 16244 31904 16250
rect 31852 16186 31904 16192
rect 32048 16114 32076 17274
rect 32036 16108 32088 16114
rect 32036 16050 32088 16056
rect 31576 15428 31628 15434
rect 31576 15370 31628 15376
rect 31484 15088 31536 15094
rect 31484 15030 31536 15036
rect 31496 13682 31524 15030
rect 31588 14482 31616 15370
rect 32232 15026 32260 18294
rect 32416 18086 32444 18906
rect 32588 18760 32640 18766
rect 32588 18702 32640 18708
rect 32496 18624 32548 18630
rect 32496 18566 32548 18572
rect 32508 18290 32536 18566
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 32404 18080 32456 18086
rect 32404 18022 32456 18028
rect 32600 17202 32628 18702
rect 32692 18290 32720 19246
rect 32784 18766 32812 19306
rect 32864 19168 32916 19174
rect 32864 19110 32916 19116
rect 32956 19168 33008 19174
rect 32956 19110 33008 19116
rect 32876 18902 32904 19110
rect 32864 18896 32916 18902
rect 32864 18838 32916 18844
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32968 18698 32996 19110
rect 32956 18692 33008 18698
rect 32956 18634 33008 18640
rect 32680 18284 32732 18290
rect 32680 18226 32732 18232
rect 32692 17882 32720 18226
rect 32968 18034 32996 18634
rect 32876 18006 33088 18034
rect 32680 17876 32732 17882
rect 32680 17818 32732 17824
rect 32876 17202 32904 18006
rect 33060 17882 33088 18006
rect 32956 17876 33008 17882
rect 32956 17818 33008 17824
rect 33048 17876 33100 17882
rect 33048 17818 33100 17824
rect 32968 17202 32996 17818
rect 33140 17536 33192 17542
rect 33140 17478 33192 17484
rect 33152 17338 33180 17478
rect 33140 17332 33192 17338
rect 33140 17274 33192 17280
rect 33244 17202 33272 22986
rect 33336 22642 33364 23598
rect 33980 23594 34008 25230
rect 34152 24608 34204 24614
rect 34152 24550 34204 24556
rect 34164 23798 34192 24550
rect 34152 23792 34204 23798
rect 34152 23734 34204 23740
rect 33968 23588 34020 23594
rect 33968 23530 34020 23536
rect 33324 22636 33376 22642
rect 33324 22578 33376 22584
rect 33784 22636 33836 22642
rect 33784 22578 33836 22584
rect 33796 22438 33824 22578
rect 33784 22432 33836 22438
rect 33784 22374 33836 22380
rect 33796 22098 33824 22374
rect 33784 22092 33836 22098
rect 33784 22034 33836 22040
rect 33416 21956 33468 21962
rect 33416 21898 33468 21904
rect 33428 21622 33456 21898
rect 34256 21894 34284 25774
rect 34440 25362 34468 27542
rect 34532 27470 34560 27814
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35360 27674 35388 27950
rect 36544 27872 36596 27878
rect 36544 27814 36596 27820
rect 35348 27668 35400 27674
rect 35348 27610 35400 27616
rect 36556 27470 36584 27814
rect 36740 27674 36768 28494
rect 37096 28484 37148 28490
rect 37096 28426 37148 28432
rect 37108 28150 37136 28426
rect 37924 28416 37976 28422
rect 37924 28358 37976 28364
rect 37096 28144 37148 28150
rect 37096 28086 37148 28092
rect 36728 27668 36780 27674
rect 36728 27610 36780 27616
rect 34520 27464 34572 27470
rect 34520 27406 34572 27412
rect 35440 27464 35492 27470
rect 35440 27406 35492 27412
rect 36544 27464 36596 27470
rect 36544 27406 36596 27412
rect 36912 27464 36964 27470
rect 36912 27406 36964 27412
rect 34532 27062 34560 27406
rect 35452 27130 35480 27406
rect 36360 27328 36412 27334
rect 36360 27270 36412 27276
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35440 27124 35492 27130
rect 35440 27066 35492 27072
rect 34520 27056 34572 27062
rect 34520 26998 34572 27004
rect 35532 26988 35584 26994
rect 35532 26930 35584 26936
rect 35624 26988 35676 26994
rect 35624 26930 35676 26936
rect 34612 26784 34664 26790
rect 34612 26726 34664 26732
rect 34624 26382 34652 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34612 26376 34664 26382
rect 35544 26330 35572 26930
rect 34612 26318 34664 26324
rect 34520 26308 34572 26314
rect 34520 26250 34572 26256
rect 34428 25356 34480 25362
rect 34428 25298 34480 25304
rect 34244 21888 34296 21894
rect 34244 21830 34296 21836
rect 33416 21616 33468 21622
rect 33416 21558 33468 21564
rect 33428 20534 33456 21558
rect 34336 21344 34388 21350
rect 34440 21298 34468 25298
rect 34532 25294 34560 26250
rect 34520 25288 34572 25294
rect 34520 25230 34572 25236
rect 34532 24954 34560 25230
rect 34520 24948 34572 24954
rect 34520 24890 34572 24896
rect 34624 24834 34652 26318
rect 35072 26308 35124 26314
rect 35072 26250 35124 26256
rect 35452 26302 35572 26330
rect 35636 26314 35664 26930
rect 35624 26308 35676 26314
rect 35084 25974 35112 26250
rect 34796 25968 34848 25974
rect 34796 25910 34848 25916
rect 35072 25968 35124 25974
rect 35072 25910 35124 25916
rect 34704 25696 34756 25702
rect 34704 25638 34756 25644
rect 34716 25208 34744 25638
rect 34808 25362 34836 25910
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34886 25392 34942 25401
rect 34796 25356 34848 25362
rect 34886 25327 34942 25336
rect 34796 25298 34848 25304
rect 34900 25294 34928 25327
rect 35452 25294 35480 26302
rect 35624 26250 35676 26256
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 34888 25288 34940 25294
rect 34888 25230 34940 25236
rect 35440 25288 35492 25294
rect 35440 25230 35492 25236
rect 36084 25288 36136 25294
rect 36084 25230 36136 25236
rect 34796 25220 34848 25226
rect 34716 25180 34796 25208
rect 34796 25162 34848 25168
rect 34388 21292 34468 21298
rect 34336 21286 34468 21292
rect 34348 21270 34468 21286
rect 33416 20528 33468 20534
rect 33416 20470 33468 20476
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33704 19922 33732 20402
rect 34058 20360 34114 20369
rect 34058 20295 34114 20304
rect 33968 20256 34020 20262
rect 33968 20198 34020 20204
rect 33692 19916 33744 19922
rect 33692 19858 33744 19864
rect 33416 19168 33468 19174
rect 33416 19110 33468 19116
rect 33428 18766 33456 19110
rect 33508 18896 33560 18902
rect 33508 18838 33560 18844
rect 33704 18850 33732 19858
rect 33980 19854 34008 20198
rect 34072 20058 34100 20295
rect 34440 20262 34468 21270
rect 34532 24806 34652 24834
rect 34532 21146 34560 24806
rect 34808 24342 34836 25162
rect 34888 25152 34940 25158
rect 34888 25094 34940 25100
rect 34900 24750 34928 25094
rect 35348 24948 35400 24954
rect 35348 24890 35400 24896
rect 34888 24744 34940 24750
rect 34888 24686 34940 24692
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24426 35388 24890
rect 35268 24398 35388 24426
rect 34796 24336 34848 24342
rect 34796 24278 34848 24284
rect 34704 23792 34756 23798
rect 34704 23734 34756 23740
rect 34716 23610 34744 23734
rect 34808 23730 34836 24278
rect 35268 23730 35296 24398
rect 35452 24324 35480 25230
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 36096 24954 36124 25230
rect 36084 24948 36136 24954
rect 36084 24890 36136 24896
rect 36176 24880 36228 24886
rect 36176 24822 36228 24828
rect 35360 24296 35480 24324
rect 35360 23730 35388 24296
rect 35992 24132 36044 24138
rect 35992 24074 36044 24080
rect 35440 24064 35492 24070
rect 35440 24006 35492 24012
rect 35452 23798 35480 24006
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 36004 23798 36032 24074
rect 35440 23792 35492 23798
rect 35440 23734 35492 23740
rect 35992 23792 36044 23798
rect 35992 23734 36044 23740
rect 34796 23724 34848 23730
rect 34796 23666 34848 23672
rect 35256 23724 35308 23730
rect 35256 23666 35308 23672
rect 35348 23724 35400 23730
rect 35348 23666 35400 23672
rect 34624 23582 34744 23610
rect 34624 22030 34652 23582
rect 34704 23520 34756 23526
rect 34704 23462 34756 23468
rect 34716 23050 34744 23462
rect 34808 23118 34836 23666
rect 35268 23474 35296 23666
rect 36084 23588 36136 23594
rect 36084 23530 36136 23536
rect 35268 23446 35388 23474
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35360 23118 35388 23446
rect 35992 23316 36044 23322
rect 35992 23258 36044 23264
rect 34796 23112 34848 23118
rect 34796 23054 34848 23060
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 34704 23044 34756 23050
rect 34704 22986 34756 22992
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 35624 22636 35676 22642
rect 35624 22578 35676 22584
rect 35636 22438 35664 22578
rect 35624 22432 35676 22438
rect 35624 22374 35676 22380
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35636 22166 35664 22374
rect 35624 22160 35676 22166
rect 35624 22102 35676 22108
rect 34612 22024 34664 22030
rect 34612 21966 34664 21972
rect 34520 21140 34572 21146
rect 34520 21082 34572 21088
rect 34520 20936 34572 20942
rect 34520 20878 34572 20884
rect 34532 20398 34560 20878
rect 34624 20874 34652 21966
rect 36004 21962 36032 23258
rect 35992 21956 36044 21962
rect 35992 21898 36044 21904
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 34704 21480 34756 21486
rect 34704 21422 34756 21428
rect 35440 21480 35492 21486
rect 35440 21422 35492 21428
rect 34612 20868 34664 20874
rect 34612 20810 34664 20816
rect 34520 20392 34572 20398
rect 34520 20334 34572 20340
rect 34428 20256 34480 20262
rect 34428 20198 34480 20204
rect 34060 20052 34112 20058
rect 34060 19994 34112 20000
rect 34440 19922 34468 20198
rect 34428 19916 34480 19922
rect 34428 19858 34480 19864
rect 33968 19848 34020 19854
rect 33968 19790 34020 19796
rect 34440 18850 34468 19858
rect 34532 18902 34560 20334
rect 34624 19854 34652 20810
rect 34716 20602 34744 21422
rect 35348 21412 35400 21418
rect 35348 21354 35400 21360
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 21140 34848 21146
rect 34796 21082 34848 21088
rect 34704 20596 34756 20602
rect 34704 20538 34756 20544
rect 34612 19848 34664 19854
rect 34612 19790 34664 19796
rect 34624 19174 34652 19790
rect 34612 19168 34664 19174
rect 34612 19110 34664 19116
rect 33520 18766 33548 18838
rect 33704 18822 33824 18850
rect 34348 18834 34468 18850
rect 34520 18896 34572 18902
rect 34520 18838 34572 18844
rect 34808 18850 34836 21082
rect 34980 20800 35032 20806
rect 34980 20742 35032 20748
rect 34992 20466 35020 20742
rect 35360 20466 35388 21354
rect 34980 20460 35032 20466
rect 34980 20402 35032 20408
rect 35348 20460 35400 20466
rect 35348 20402 35400 20408
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35452 19922 35480 21422
rect 36004 20942 36032 21898
rect 35992 20936 36044 20942
rect 35992 20878 36044 20884
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35440 19916 35492 19922
rect 35440 19858 35492 19864
rect 34888 19848 34940 19854
rect 34888 19790 34940 19796
rect 35348 19848 35400 19854
rect 35348 19790 35400 19796
rect 34900 19378 34928 19790
rect 35164 19780 35216 19786
rect 35164 19722 35216 19728
rect 35176 19446 35204 19722
rect 35164 19440 35216 19446
rect 35164 19382 35216 19388
rect 35360 19378 35388 19790
rect 35452 19446 35480 19858
rect 35992 19712 36044 19718
rect 35992 19654 36044 19660
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35440 19440 35492 19446
rect 35440 19382 35492 19388
rect 36004 19378 36032 19654
rect 34888 19372 34940 19378
rect 34888 19314 34940 19320
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 35992 19372 36044 19378
rect 35992 19314 36044 19320
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 33796 18766 33824 18822
rect 34336 18828 34468 18834
rect 34388 18822 34468 18828
rect 34808 18822 34928 18850
rect 34336 18770 34388 18776
rect 33324 18760 33376 18766
rect 33324 18702 33376 18708
rect 33416 18760 33468 18766
rect 33416 18702 33468 18708
rect 33508 18760 33560 18766
rect 33508 18702 33560 18708
rect 33600 18760 33652 18766
rect 33600 18702 33652 18708
rect 33784 18760 33836 18766
rect 33784 18702 33836 18708
rect 34060 18760 34112 18766
rect 34060 18702 34112 18708
rect 33336 18426 33364 18702
rect 33324 18420 33376 18426
rect 33324 18362 33376 18368
rect 33416 18080 33468 18086
rect 33416 18022 33468 18028
rect 33324 17536 33376 17542
rect 33324 17478 33376 17484
rect 32588 17196 32640 17202
rect 32588 17138 32640 17144
rect 32864 17196 32916 17202
rect 32864 17138 32916 17144
rect 32956 17196 33008 17202
rect 32956 17138 33008 17144
rect 33232 17196 33284 17202
rect 33232 17138 33284 17144
rect 32404 16992 32456 16998
rect 32404 16934 32456 16940
rect 32416 16114 32444 16934
rect 32600 16794 32628 17138
rect 32954 17096 33010 17105
rect 32954 17031 33010 17040
rect 32588 16788 32640 16794
rect 32588 16730 32640 16736
rect 32680 16448 32732 16454
rect 32680 16390 32732 16396
rect 32692 16114 32720 16390
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32680 16108 32732 16114
rect 32680 16050 32732 16056
rect 32220 15020 32272 15026
rect 32220 14962 32272 14968
rect 32036 14612 32088 14618
rect 32036 14554 32088 14560
rect 31576 14476 31628 14482
rect 31576 14418 31628 14424
rect 31576 14340 31628 14346
rect 31576 14282 31628 14288
rect 31588 14074 31616 14282
rect 31944 14272 31996 14278
rect 31944 14214 31996 14220
rect 31576 14068 31628 14074
rect 31576 14010 31628 14016
rect 31956 13870 31984 14214
rect 31944 13864 31996 13870
rect 31944 13806 31996 13812
rect 31496 13654 31616 13682
rect 31484 12640 31536 12646
rect 31484 12582 31536 12588
rect 31496 12306 31524 12582
rect 31484 12300 31536 12306
rect 31484 12242 31536 12248
rect 31392 11688 31444 11694
rect 31392 11630 31444 11636
rect 31208 11552 31260 11558
rect 31208 11494 31260 11500
rect 31220 11150 31248 11494
rect 31208 11144 31260 11150
rect 31206 11112 31208 11121
rect 31260 11112 31262 11121
rect 31206 11047 31262 11056
rect 30932 10056 30984 10062
rect 30932 9998 30984 10004
rect 30944 9450 30972 9998
rect 31208 9988 31260 9994
rect 31208 9930 31260 9936
rect 31220 9722 31248 9930
rect 31208 9716 31260 9722
rect 31208 9658 31260 9664
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 30932 9444 30984 9450
rect 30932 9386 30984 9392
rect 31036 9330 31064 9522
rect 30944 9302 31064 9330
rect 30944 7410 30972 9302
rect 31300 9172 31352 9178
rect 31300 9114 31352 9120
rect 31208 8968 31260 8974
rect 31208 8910 31260 8916
rect 31024 8492 31076 8498
rect 31024 8434 31076 8440
rect 31116 8492 31168 8498
rect 31220 8480 31248 8910
rect 31312 8566 31340 9114
rect 31404 8906 31432 11630
rect 31588 9625 31616 13654
rect 31956 13326 31984 13806
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31944 13184 31996 13190
rect 31944 13126 31996 13132
rect 31668 12980 31720 12986
rect 31668 12922 31720 12928
rect 31680 11558 31708 12922
rect 31852 12164 31904 12170
rect 31852 12106 31904 12112
rect 31864 11830 31892 12106
rect 31852 11824 31904 11830
rect 31852 11766 31904 11772
rect 31668 11552 31720 11558
rect 31668 11494 31720 11500
rect 31574 9616 31630 9625
rect 31574 9551 31630 9560
rect 31852 9580 31904 9586
rect 31484 9172 31536 9178
rect 31484 9114 31536 9120
rect 31496 8974 31524 9114
rect 31484 8968 31536 8974
rect 31484 8910 31536 8916
rect 31588 8906 31616 9551
rect 31852 9522 31904 9528
rect 31760 9444 31812 9450
rect 31760 9386 31812 9392
rect 31666 9344 31722 9353
rect 31666 9279 31722 9288
rect 31680 8974 31708 9279
rect 31668 8968 31720 8974
rect 31668 8910 31720 8916
rect 31392 8900 31444 8906
rect 31392 8842 31444 8848
rect 31576 8900 31628 8906
rect 31576 8842 31628 8848
rect 31484 8832 31536 8838
rect 31484 8774 31536 8780
rect 31300 8560 31352 8566
rect 31300 8502 31352 8508
rect 31496 8498 31524 8774
rect 31168 8452 31248 8480
rect 31392 8492 31444 8498
rect 31116 8434 31168 8440
rect 31392 8434 31444 8440
rect 31484 8492 31536 8498
rect 31484 8434 31536 8440
rect 31036 7886 31064 8434
rect 31404 8362 31432 8434
rect 31116 8356 31168 8362
rect 31116 8298 31168 8304
rect 31392 8356 31444 8362
rect 31392 8298 31444 8304
rect 31128 7954 31156 8298
rect 31116 7948 31168 7954
rect 31116 7890 31168 7896
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 31024 7744 31076 7750
rect 31024 7686 31076 7692
rect 31036 7410 31064 7686
rect 30932 7404 30984 7410
rect 30932 7346 30984 7352
rect 31024 7404 31076 7410
rect 31024 7346 31076 7352
rect 30944 5234 30972 7346
rect 31404 6866 31432 8298
rect 31680 7886 31708 8910
rect 31772 8634 31800 9386
rect 31864 9178 31892 9522
rect 31852 9172 31904 9178
rect 31852 9114 31904 9120
rect 31760 8628 31812 8634
rect 31812 8588 31892 8616
rect 31760 8570 31812 8576
rect 31484 7880 31536 7886
rect 31484 7822 31536 7828
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 31392 6860 31444 6866
rect 31392 6802 31444 6808
rect 31404 6390 31432 6802
rect 31496 6458 31524 7822
rect 31760 7744 31812 7750
rect 31760 7686 31812 7692
rect 31772 7002 31800 7686
rect 31864 7546 31892 8588
rect 31852 7540 31904 7546
rect 31852 7482 31904 7488
rect 31760 6996 31812 7002
rect 31760 6938 31812 6944
rect 31668 6792 31720 6798
rect 31668 6734 31720 6740
rect 31484 6452 31536 6458
rect 31484 6394 31536 6400
rect 31392 6384 31444 6390
rect 31392 6326 31444 6332
rect 31496 6322 31524 6394
rect 31484 6316 31536 6322
rect 31484 6258 31536 6264
rect 31208 6112 31260 6118
rect 31208 6054 31260 6060
rect 31220 5234 31248 6054
rect 30932 5228 30984 5234
rect 30932 5170 30984 5176
rect 31208 5228 31260 5234
rect 31208 5170 31260 5176
rect 31496 4622 31524 6258
rect 31484 4616 31536 4622
rect 31484 4558 31536 4564
rect 31680 4486 31708 6734
rect 31772 6390 31800 6938
rect 31864 6798 31892 7482
rect 31852 6792 31904 6798
rect 31852 6734 31904 6740
rect 31760 6384 31812 6390
rect 31760 6326 31812 6332
rect 31864 5914 31892 6734
rect 31852 5908 31904 5914
rect 31852 5850 31904 5856
rect 31760 5704 31812 5710
rect 31864 5692 31892 5850
rect 31812 5664 31892 5692
rect 31760 5646 31812 5652
rect 31668 4480 31720 4486
rect 31668 4422 31720 4428
rect 30840 4140 30892 4146
rect 30840 4082 30892 4088
rect 31772 3670 31800 5646
rect 31956 4162 31984 13126
rect 32048 12850 32076 14554
rect 32864 14340 32916 14346
rect 32864 14282 32916 14288
rect 32876 14074 32904 14282
rect 32588 14068 32640 14074
rect 32864 14068 32916 14074
rect 32588 14010 32640 14016
rect 32692 14028 32864 14056
rect 32128 14000 32180 14006
rect 32128 13942 32180 13948
rect 32402 13968 32458 13977
rect 32140 13530 32168 13942
rect 32402 13903 32404 13912
rect 32456 13903 32458 13912
rect 32404 13874 32456 13880
rect 32128 13524 32180 13530
rect 32128 13466 32180 13472
rect 32036 12844 32088 12850
rect 32036 12786 32088 12792
rect 32140 11830 32168 13466
rect 32312 12980 32364 12986
rect 32416 12968 32444 13874
rect 32600 13462 32628 14010
rect 32588 13456 32640 13462
rect 32588 13398 32640 13404
rect 32364 12940 32444 12968
rect 32312 12922 32364 12928
rect 32128 11824 32180 11830
rect 32128 11766 32180 11772
rect 32128 10600 32180 10606
rect 32128 10542 32180 10548
rect 32140 8566 32168 10542
rect 32404 10464 32456 10470
rect 32404 10406 32456 10412
rect 32416 9654 32444 10406
rect 32692 10266 32720 14028
rect 32864 14010 32916 14016
rect 32772 12844 32824 12850
rect 32772 12786 32824 12792
rect 32784 12374 32812 12786
rect 32864 12708 32916 12714
rect 32864 12650 32916 12656
rect 32876 12442 32904 12650
rect 32864 12436 32916 12442
rect 32864 12378 32916 12384
rect 32772 12368 32824 12374
rect 32772 12310 32824 12316
rect 32876 12170 32904 12378
rect 32864 12164 32916 12170
rect 32864 12106 32916 12112
rect 32968 10810 32996 17031
rect 33232 16108 33284 16114
rect 33232 16050 33284 16056
rect 33244 15434 33272 16050
rect 33232 15428 33284 15434
rect 33232 15370 33284 15376
rect 33244 15162 33272 15370
rect 33232 15156 33284 15162
rect 33232 15098 33284 15104
rect 33138 15056 33194 15065
rect 33244 15026 33272 15098
rect 33138 14991 33140 15000
rect 33192 14991 33194 15000
rect 33232 15020 33284 15026
rect 33140 14962 33192 14968
rect 33232 14962 33284 14968
rect 33048 14612 33100 14618
rect 33048 14554 33100 14560
rect 33060 13938 33088 14554
rect 33152 14414 33180 14962
rect 33232 14884 33284 14890
rect 33232 14826 33284 14832
rect 33244 14618 33272 14826
rect 33232 14612 33284 14618
rect 33232 14554 33284 14560
rect 33140 14408 33192 14414
rect 33140 14350 33192 14356
rect 33048 13932 33100 13938
rect 33048 13874 33100 13880
rect 33152 13734 33180 14350
rect 33140 13728 33192 13734
rect 33140 13670 33192 13676
rect 33336 12986 33364 17478
rect 33428 17134 33456 18022
rect 33612 17678 33640 18702
rect 33796 18358 33824 18702
rect 33876 18624 33928 18630
rect 33876 18566 33928 18572
rect 33888 18358 33916 18566
rect 33784 18352 33836 18358
rect 33784 18294 33836 18300
rect 33876 18352 33928 18358
rect 33876 18294 33928 18300
rect 33876 18216 33928 18222
rect 33876 18158 33928 18164
rect 33784 17876 33836 17882
rect 33784 17818 33836 17824
rect 33600 17672 33652 17678
rect 33600 17614 33652 17620
rect 33796 17542 33824 17818
rect 33784 17536 33836 17542
rect 33784 17478 33836 17484
rect 33598 17232 33654 17241
rect 33598 17167 33600 17176
rect 33652 17167 33654 17176
rect 33600 17138 33652 17144
rect 33416 17128 33468 17134
rect 33416 17070 33468 17076
rect 33428 16046 33456 17070
rect 33888 16590 33916 18158
rect 34072 17202 34100 18702
rect 34060 17196 34112 17202
rect 34060 17138 34112 17144
rect 34072 17066 34100 17138
rect 34348 17134 34376 18770
rect 34900 18426 34928 18822
rect 35360 18766 35388 19314
rect 35440 18964 35492 18970
rect 35440 18906 35492 18912
rect 35348 18760 35400 18766
rect 35348 18702 35400 18708
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 34888 18420 34940 18426
rect 34888 18362 34940 18368
rect 34808 18204 34836 18362
rect 34888 18216 34940 18222
rect 34808 18176 34888 18204
rect 34520 18080 34572 18086
rect 34520 18022 34572 18028
rect 34428 17876 34480 17882
rect 34532 17864 34560 18022
rect 34480 17836 34560 17864
rect 34428 17818 34480 17824
rect 34520 17536 34572 17542
rect 34520 17478 34572 17484
rect 34532 17202 34560 17478
rect 34808 17202 34836 18176
rect 34888 18158 34940 18164
rect 35360 18086 35388 18702
rect 35452 18358 35480 18906
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35440 18352 35492 18358
rect 35440 18294 35492 18300
rect 35348 18080 35400 18086
rect 35348 18022 35400 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17746 35388 18022
rect 35348 17740 35400 17746
rect 35348 17682 35400 17688
rect 35452 17678 35480 18294
rect 36096 18290 36124 23530
rect 36188 23322 36216 24822
rect 36176 23316 36228 23322
rect 36176 23258 36228 23264
rect 36176 23180 36228 23186
rect 36176 23122 36228 23128
rect 36188 22982 36216 23122
rect 36176 22976 36228 22982
rect 36174 22944 36176 22953
rect 36228 22944 36230 22953
rect 36174 22879 36230 22888
rect 36176 20800 36228 20806
rect 36176 20742 36228 20748
rect 36188 20330 36216 20742
rect 36176 20324 36228 20330
rect 36176 20266 36228 20272
rect 36188 19378 36216 20266
rect 36268 20052 36320 20058
rect 36268 19994 36320 20000
rect 36280 19378 36308 19994
rect 36176 19372 36228 19378
rect 36176 19314 36228 19320
rect 36268 19372 36320 19378
rect 36268 19314 36320 19320
rect 36176 18760 36228 18766
rect 36176 18702 36228 18708
rect 36188 18426 36216 18702
rect 36176 18420 36228 18426
rect 36176 18362 36228 18368
rect 35532 18284 35584 18290
rect 35532 18226 35584 18232
rect 36084 18284 36136 18290
rect 36084 18226 36136 18232
rect 35440 17672 35492 17678
rect 35440 17614 35492 17620
rect 35348 17536 35400 17542
rect 35348 17478 35400 17484
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34796 17196 34848 17202
rect 34796 17138 34848 17144
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34060 17060 34112 17066
rect 34060 17002 34112 17008
rect 34152 16992 34204 16998
rect 34152 16934 34204 16940
rect 34244 16992 34296 16998
rect 34244 16934 34296 16940
rect 33508 16584 33560 16590
rect 33508 16526 33560 16532
rect 33876 16584 33928 16590
rect 33876 16526 33928 16532
rect 33520 16454 33548 16526
rect 33508 16448 33560 16454
rect 33508 16390 33560 16396
rect 33888 16114 33916 16526
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33416 16040 33468 16046
rect 33416 15982 33468 15988
rect 34164 15620 34192 16934
rect 34256 16182 34284 16934
rect 34808 16250 34836 17138
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35256 16448 35308 16454
rect 35360 16436 35388 17478
rect 35452 16522 35480 17614
rect 35544 17542 35572 18226
rect 36096 18086 36124 18226
rect 36268 18216 36320 18222
rect 36268 18158 36320 18164
rect 36084 18080 36136 18086
rect 36084 18022 36136 18028
rect 35532 17536 35584 17542
rect 35532 17478 35584 17484
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 35440 16516 35492 16522
rect 35440 16458 35492 16464
rect 36084 16516 36136 16522
rect 36084 16458 36136 16464
rect 35308 16408 35388 16436
rect 35256 16390 35308 16396
rect 34796 16244 34848 16250
rect 34796 16186 34848 16192
rect 34244 16176 34296 16182
rect 34244 16118 34296 16124
rect 35268 16114 35296 16390
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35256 16108 35308 16114
rect 35256 16050 35308 16056
rect 35268 15978 35296 16050
rect 36096 15978 36124 16458
rect 35256 15972 35308 15978
rect 35256 15914 35308 15920
rect 36084 15972 36136 15978
rect 36084 15914 36136 15920
rect 35992 15904 36044 15910
rect 35992 15846 36044 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 36004 15638 36032 15846
rect 34428 15632 34480 15638
rect 34164 15592 34428 15620
rect 34428 15574 34480 15580
rect 35992 15632 36044 15638
rect 35992 15574 36044 15580
rect 33692 15496 33744 15502
rect 33692 15438 33744 15444
rect 33508 15360 33560 15366
rect 33508 15302 33560 15308
rect 33520 14958 33548 15302
rect 33508 14952 33560 14958
rect 33508 14894 33560 14900
rect 33416 14408 33468 14414
rect 33416 14350 33468 14356
rect 33428 13977 33456 14350
rect 33508 14340 33560 14346
rect 33508 14282 33560 14288
rect 33520 14006 33548 14282
rect 33508 14000 33560 14006
rect 33414 13968 33470 13977
rect 33508 13942 33560 13948
rect 33414 13903 33470 13912
rect 33324 12980 33376 12986
rect 33324 12922 33376 12928
rect 33428 12730 33456 13903
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33612 12850 33640 13806
rect 33704 13734 33732 15438
rect 34244 15428 34296 15434
rect 34244 15370 34296 15376
rect 34336 15428 34388 15434
rect 34336 15370 34388 15376
rect 34256 14822 34284 15370
rect 34244 14816 34296 14822
rect 34244 14758 34296 14764
rect 33876 14544 33928 14550
rect 33876 14486 33928 14492
rect 33888 13954 33916 14486
rect 33968 14272 34020 14278
rect 33968 14214 34020 14220
rect 34152 14272 34204 14278
rect 34152 14214 34204 14220
rect 33796 13938 33916 13954
rect 33784 13932 33916 13938
rect 33836 13926 33916 13932
rect 33980 13954 34008 14214
rect 34058 13968 34114 13977
rect 33980 13926 34058 13954
rect 34164 13938 34192 14214
rect 34058 13903 34060 13912
rect 33784 13874 33836 13880
rect 34112 13903 34114 13912
rect 34152 13932 34204 13938
rect 34060 13874 34112 13880
rect 34152 13874 34204 13880
rect 33692 13728 33744 13734
rect 33692 13670 33744 13676
rect 33600 12844 33652 12850
rect 33600 12786 33652 12792
rect 33428 12702 33548 12730
rect 33416 12640 33468 12646
rect 33416 12582 33468 12588
rect 33232 12368 33284 12374
rect 33232 12310 33284 12316
rect 33244 11558 33272 12310
rect 33428 12238 33456 12582
rect 33520 12238 33548 12702
rect 33612 12306 33640 12786
rect 33600 12300 33652 12306
rect 33600 12242 33652 12248
rect 33416 12232 33468 12238
rect 33416 12174 33468 12180
rect 33508 12232 33560 12238
rect 33508 12174 33560 12180
rect 33232 11552 33284 11558
rect 33232 11494 33284 11500
rect 33600 11552 33652 11558
rect 33600 11494 33652 11500
rect 32956 10804 33008 10810
rect 32956 10746 33008 10752
rect 32956 10668 33008 10674
rect 32956 10610 33008 10616
rect 33232 10668 33284 10674
rect 33232 10610 33284 10616
rect 33324 10668 33376 10674
rect 33324 10610 33376 10616
rect 32968 10266 32996 10610
rect 32680 10260 32732 10266
rect 32680 10202 32732 10208
rect 32956 10260 33008 10266
rect 32956 10202 33008 10208
rect 32496 10056 32548 10062
rect 32496 9998 32548 10004
rect 32404 9648 32456 9654
rect 32404 9590 32456 9596
rect 32218 9072 32274 9081
rect 32218 9007 32274 9016
rect 32232 8974 32260 9007
rect 32220 8968 32272 8974
rect 32404 8968 32456 8974
rect 32272 8928 32352 8956
rect 32220 8910 32272 8916
rect 32220 8832 32272 8838
rect 32220 8774 32272 8780
rect 32128 8560 32180 8566
rect 32128 8502 32180 8508
rect 32232 8430 32260 8774
rect 32220 8424 32272 8430
rect 32220 8366 32272 8372
rect 32324 7954 32352 8928
rect 32508 8956 32536 9998
rect 32692 9994 32720 10202
rect 33048 10056 33100 10062
rect 33048 9998 33100 10004
rect 32680 9988 32732 9994
rect 32680 9930 32732 9936
rect 32692 9450 32720 9930
rect 33060 9518 33088 9998
rect 33048 9512 33100 9518
rect 33244 9489 33272 10610
rect 33048 9454 33100 9460
rect 33230 9480 33286 9489
rect 32680 9444 32732 9450
rect 33230 9415 33286 9424
rect 32680 9386 32732 9392
rect 33232 9376 33284 9382
rect 32770 9344 32826 9353
rect 33336 9353 33364 10610
rect 33612 10606 33640 11494
rect 33796 10742 33824 13874
rect 34256 13802 34284 14758
rect 34244 13796 34296 13802
rect 34244 13738 34296 13744
rect 34152 13388 34204 13394
rect 34256 13376 34284 13738
rect 34204 13348 34284 13376
rect 34152 13330 34204 13336
rect 33876 12912 33928 12918
rect 33876 12854 33928 12860
rect 33888 12434 33916 12854
rect 33888 12406 34100 12434
rect 33968 12096 34020 12102
rect 33968 12038 34020 12044
rect 33980 11830 34008 12038
rect 33968 11824 34020 11830
rect 33968 11766 34020 11772
rect 33784 10736 33836 10742
rect 33784 10678 33836 10684
rect 33600 10600 33652 10606
rect 33600 10542 33652 10548
rect 33876 10600 33928 10606
rect 33876 10542 33928 10548
rect 33416 9512 33468 9518
rect 33416 9454 33468 9460
rect 33232 9318 33284 9324
rect 33322 9344 33378 9353
rect 32770 9279 32826 9288
rect 32456 8928 32536 8956
rect 32404 8910 32456 8916
rect 32784 8906 32812 9279
rect 32772 8900 32824 8906
rect 32772 8842 32824 8848
rect 33048 8900 33100 8906
rect 33048 8842 33100 8848
rect 32588 8832 32640 8838
rect 32588 8774 32640 8780
rect 32680 8832 32732 8838
rect 32680 8774 32732 8780
rect 32600 8566 32628 8774
rect 32588 8560 32640 8566
rect 32588 8502 32640 8508
rect 32312 7948 32364 7954
rect 32312 7890 32364 7896
rect 32036 7880 32088 7886
rect 32036 7822 32088 7828
rect 32048 5846 32076 7822
rect 32600 7818 32628 8502
rect 32692 8498 32720 8774
rect 33060 8634 33088 8842
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 32772 8560 32824 8566
rect 32772 8502 32824 8508
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32784 8362 32812 8502
rect 33244 8430 33272 9318
rect 33322 9279 33378 9288
rect 33428 8537 33456 9454
rect 33612 9042 33640 10542
rect 33888 10266 33916 10542
rect 33876 10260 33928 10266
rect 33876 10202 33928 10208
rect 33876 9920 33928 9926
rect 33876 9862 33928 9868
rect 33784 9444 33836 9450
rect 33784 9386 33836 9392
rect 33796 9353 33824 9386
rect 33782 9344 33838 9353
rect 33782 9279 33838 9288
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 33414 8528 33470 8537
rect 33414 8463 33470 8472
rect 33888 8430 33916 9862
rect 34072 9330 34100 12406
rect 34164 12238 34192 13330
rect 34244 12368 34296 12374
rect 34244 12310 34296 12316
rect 34256 12238 34284 12310
rect 34152 12232 34204 12238
rect 34152 12174 34204 12180
rect 34244 12232 34296 12238
rect 34244 12174 34296 12180
rect 34164 9500 34192 12174
rect 34348 9926 34376 15370
rect 34440 14618 34468 15574
rect 35440 15564 35492 15570
rect 35440 15506 35492 15512
rect 34796 15496 34848 15502
rect 34796 15438 34848 15444
rect 35348 15496 35400 15502
rect 35348 15438 35400 15444
rect 34704 14884 34756 14890
rect 34704 14826 34756 14832
rect 34428 14612 34480 14618
rect 34428 14554 34480 14560
rect 34716 14226 34744 14826
rect 34808 14822 34836 15438
rect 34796 14816 34848 14822
rect 34796 14758 34848 14764
rect 34808 14346 34836 14758
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14618 35388 15438
rect 35452 15094 35480 15506
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35440 15088 35492 15094
rect 35440 15030 35492 15036
rect 36096 14958 36124 15914
rect 36084 14952 36136 14958
rect 36084 14894 36136 14900
rect 35348 14612 35400 14618
rect 35348 14554 35400 14560
rect 35808 14476 35860 14482
rect 35808 14418 35860 14424
rect 35820 14346 35848 14418
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 34796 14340 34848 14346
rect 34796 14282 34848 14288
rect 35808 14340 35860 14346
rect 35808 14282 35860 14288
rect 35348 14272 35400 14278
rect 34716 14198 34836 14226
rect 35348 14214 35400 14220
rect 34704 13184 34756 13190
rect 34704 13126 34756 13132
rect 34716 12918 34744 13126
rect 34808 12918 34836 14198
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34704 12912 34756 12918
rect 34704 12854 34756 12860
rect 34796 12912 34848 12918
rect 34796 12854 34848 12860
rect 34428 12776 34480 12782
rect 34428 12718 34480 12724
rect 34440 11778 34468 12718
rect 34520 12436 34572 12442
rect 34520 12378 34572 12384
rect 34532 12170 34560 12378
rect 34520 12164 34572 12170
rect 34520 12106 34572 12112
rect 34808 11898 34836 12854
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35360 12306 35388 14214
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 36188 14074 36216 14350
rect 36176 14068 36228 14074
rect 36176 14010 36228 14016
rect 36280 14006 36308 18158
rect 36372 17542 36400 27270
rect 36556 26926 36584 27406
rect 36924 27130 36952 27406
rect 36728 27124 36780 27130
rect 36728 27066 36780 27072
rect 36912 27124 36964 27130
rect 36912 27066 36964 27072
rect 36740 26994 36768 27066
rect 37004 27056 37056 27062
rect 37004 26998 37056 27004
rect 36728 26988 36780 26994
rect 36728 26930 36780 26936
rect 36544 26920 36596 26926
rect 36544 26862 36596 26868
rect 36556 26382 36584 26862
rect 36544 26376 36596 26382
rect 36544 26318 36596 26324
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 36464 18766 36492 24006
rect 36556 23118 36584 26318
rect 36636 25900 36688 25906
rect 36636 25842 36688 25848
rect 36648 24818 36676 25842
rect 36636 24812 36688 24818
rect 36636 24754 36688 24760
rect 36912 24064 36964 24070
rect 36912 24006 36964 24012
rect 36728 23520 36780 23526
rect 36728 23462 36780 23468
rect 36544 23112 36596 23118
rect 36544 23054 36596 23060
rect 36544 22976 36596 22982
rect 36544 22918 36596 22924
rect 36556 22642 36584 22918
rect 36544 22636 36596 22642
rect 36544 22578 36596 22584
rect 36740 22438 36768 23462
rect 36820 23112 36872 23118
rect 36820 23054 36872 23060
rect 36728 22432 36780 22438
rect 36728 22374 36780 22380
rect 36832 22250 36860 23054
rect 36740 22222 36860 22250
rect 36636 20800 36688 20806
rect 36636 20742 36688 20748
rect 36648 20466 36676 20742
rect 36636 20460 36688 20466
rect 36636 20402 36688 20408
rect 36740 19718 36768 22222
rect 36924 22094 36952 24006
rect 36832 22066 36952 22094
rect 37016 22094 37044 26998
rect 37108 25226 37136 28086
rect 37832 27532 37884 27538
rect 37832 27474 37884 27480
rect 37280 26988 37332 26994
rect 37280 26930 37332 26936
rect 37372 26988 37424 26994
rect 37372 26930 37424 26936
rect 37188 26852 37240 26858
rect 37188 26794 37240 26800
rect 37096 25220 37148 25226
rect 37096 25162 37148 25168
rect 37108 24954 37136 25162
rect 37096 24948 37148 24954
rect 37096 24890 37148 24896
rect 37200 24682 37228 26794
rect 37292 26042 37320 26930
rect 37280 26036 37332 26042
rect 37280 25978 37332 25984
rect 37384 25906 37412 26930
rect 37740 26036 37792 26042
rect 37740 25978 37792 25984
rect 37752 25906 37780 25978
rect 37372 25900 37424 25906
rect 37372 25842 37424 25848
rect 37740 25900 37792 25906
rect 37740 25842 37792 25848
rect 37648 25764 37700 25770
rect 37648 25706 37700 25712
rect 37280 25696 37332 25702
rect 37280 25638 37332 25644
rect 37292 24750 37320 25638
rect 37556 25152 37608 25158
rect 37556 25094 37608 25100
rect 37568 24818 37596 25094
rect 37660 24818 37688 25706
rect 37844 25362 37872 27474
rect 37936 27470 37964 28358
rect 38764 27538 38792 28630
rect 38752 27532 38804 27538
rect 38752 27474 38804 27480
rect 37924 27464 37976 27470
rect 37924 27406 37976 27412
rect 38108 27464 38160 27470
rect 38108 27406 38160 27412
rect 37936 27010 37964 27406
rect 38120 27130 38148 27406
rect 38660 27328 38712 27334
rect 38660 27270 38712 27276
rect 38108 27124 38160 27130
rect 38108 27066 38160 27072
rect 37936 26982 38148 27010
rect 38672 26994 38700 27270
rect 38764 26994 38792 27474
rect 38120 26790 38148 26982
rect 38384 26988 38436 26994
rect 38384 26930 38436 26936
rect 38660 26988 38712 26994
rect 38660 26930 38712 26936
rect 38752 26988 38804 26994
rect 38752 26930 38804 26936
rect 38108 26784 38160 26790
rect 38108 26726 38160 26732
rect 38120 25906 38148 26726
rect 38396 26042 38424 26930
rect 38384 26036 38436 26042
rect 38384 25978 38436 25984
rect 38108 25900 38160 25906
rect 38108 25842 38160 25848
rect 37924 25832 37976 25838
rect 37924 25774 37976 25780
rect 37832 25356 37884 25362
rect 37832 25298 37884 25304
rect 37936 24818 37964 25774
rect 37556 24812 37608 24818
rect 37556 24754 37608 24760
rect 37648 24812 37700 24818
rect 37648 24754 37700 24760
rect 37924 24812 37976 24818
rect 37924 24754 37976 24760
rect 37280 24744 37332 24750
rect 37280 24686 37332 24692
rect 37188 24676 37240 24682
rect 37188 24618 37240 24624
rect 37096 24268 37148 24274
rect 37096 24210 37148 24216
rect 37108 23866 37136 24210
rect 37096 23860 37148 23866
rect 37096 23802 37148 23808
rect 37200 23798 37228 24618
rect 37464 24132 37516 24138
rect 37464 24074 37516 24080
rect 37188 23792 37240 23798
rect 37188 23734 37240 23740
rect 37372 23656 37424 23662
rect 37372 23598 37424 23604
rect 37280 23520 37332 23526
rect 37280 23462 37332 23468
rect 37292 23186 37320 23462
rect 37280 23180 37332 23186
rect 37280 23122 37332 23128
rect 37188 23044 37240 23050
rect 37188 22986 37240 22992
rect 37200 22098 37228 22986
rect 37384 22506 37412 23598
rect 37372 22500 37424 22506
rect 37372 22442 37424 22448
rect 37016 22066 37136 22094
rect 36832 20058 36860 22066
rect 36912 20256 36964 20262
rect 36912 20198 36964 20204
rect 37004 20256 37056 20262
rect 37004 20198 37056 20204
rect 36924 20058 36952 20198
rect 36820 20052 36872 20058
rect 36820 19994 36872 20000
rect 36912 20052 36964 20058
rect 36912 19994 36964 20000
rect 37016 19938 37044 20198
rect 36832 19910 37044 19938
rect 36728 19712 36780 19718
rect 36648 19672 36728 19700
rect 36544 19236 36596 19242
rect 36544 19178 36596 19184
rect 36556 18766 36584 19178
rect 36452 18760 36504 18766
rect 36452 18702 36504 18708
rect 36544 18760 36596 18766
rect 36544 18702 36596 18708
rect 36452 18420 36504 18426
rect 36452 18362 36504 18368
rect 36464 18222 36492 18362
rect 36452 18216 36504 18222
rect 36452 18158 36504 18164
rect 36452 17808 36504 17814
rect 36452 17750 36504 17756
rect 36360 17536 36412 17542
rect 36360 17478 36412 17484
rect 36464 17270 36492 17750
rect 36556 17610 36584 18702
rect 36544 17604 36596 17610
rect 36544 17546 36596 17552
rect 36452 17264 36504 17270
rect 36452 17206 36504 17212
rect 36452 16992 36504 16998
rect 36452 16934 36504 16940
rect 36464 16658 36492 16934
rect 36544 16788 36596 16794
rect 36544 16730 36596 16736
rect 36452 16652 36504 16658
rect 36452 16594 36504 16600
rect 36556 16522 36584 16730
rect 36544 16516 36596 16522
rect 36544 16458 36596 16464
rect 36544 14816 36596 14822
rect 36544 14758 36596 14764
rect 36556 14346 36584 14758
rect 36648 14498 36676 19672
rect 36728 19654 36780 19660
rect 36726 19408 36782 19417
rect 36832 19378 36860 19910
rect 36912 19712 36964 19718
rect 36910 19680 36912 19689
rect 36964 19680 36966 19689
rect 36910 19615 36966 19624
rect 37108 19530 37136 22066
rect 37188 22092 37240 22098
rect 37476 22094 37504 24074
rect 37568 23798 37596 24754
rect 37556 23792 37608 23798
rect 37556 23734 37608 23740
rect 37476 22066 37596 22094
rect 37188 22034 37240 22040
rect 36924 19502 37136 19530
rect 36726 19343 36728 19352
rect 36780 19343 36782 19352
rect 36820 19372 36872 19378
rect 36728 19314 36780 19320
rect 36820 19314 36872 19320
rect 36924 18986 36952 19502
rect 37200 19394 37228 22034
rect 37464 21888 37516 21894
rect 37464 21830 37516 21836
rect 37476 21554 37504 21830
rect 37464 21548 37516 21554
rect 37464 21490 37516 21496
rect 37280 21344 37332 21350
rect 37280 21286 37332 21292
rect 37292 20602 37320 21286
rect 37372 21140 37424 21146
rect 37372 21082 37424 21088
rect 37280 20596 37332 20602
rect 37280 20538 37332 20544
rect 37384 19394 37412 21082
rect 37476 21010 37504 21490
rect 37568 21350 37596 22066
rect 37660 21554 37688 24754
rect 37832 24336 37884 24342
rect 37832 24278 37884 24284
rect 37844 23730 37872 24278
rect 37832 23724 37884 23730
rect 37832 23666 37884 23672
rect 37740 22704 37792 22710
rect 37740 22646 37792 22652
rect 37648 21548 37700 21554
rect 37648 21490 37700 21496
rect 37556 21344 37608 21350
rect 37556 21286 37608 21292
rect 37464 21004 37516 21010
rect 37516 20964 37596 20992
rect 37464 20946 37516 20952
rect 37464 20868 37516 20874
rect 37464 20810 37516 20816
rect 37476 20398 37504 20810
rect 37568 20602 37596 20964
rect 37556 20596 37608 20602
rect 37556 20538 37608 20544
rect 37464 20392 37516 20398
rect 37464 20334 37516 20340
rect 37200 19378 37320 19394
rect 37188 19372 37320 19378
rect 37240 19366 37320 19372
rect 37384 19366 37504 19394
rect 37188 19314 37240 19320
rect 37188 19168 37240 19174
rect 37188 19110 37240 19116
rect 36832 18958 36952 18986
rect 36728 18624 36780 18630
rect 36728 18566 36780 18572
rect 36740 18426 36768 18566
rect 36728 18420 36780 18426
rect 36728 18362 36780 18368
rect 36832 18290 36860 18958
rect 36912 18896 36964 18902
rect 36912 18838 36964 18844
rect 36820 18284 36872 18290
rect 36820 18226 36872 18232
rect 36924 16674 36952 18838
rect 37200 18766 37228 19110
rect 37292 18970 37320 19366
rect 37372 19304 37424 19310
rect 37372 19246 37424 19252
rect 37384 19145 37412 19246
rect 37370 19136 37426 19145
rect 37370 19071 37426 19080
rect 37280 18964 37332 18970
rect 37280 18906 37332 18912
rect 37476 18850 37504 19366
rect 37292 18822 37504 18850
rect 37188 18760 37240 18766
rect 37188 18702 37240 18708
rect 37004 18692 37056 18698
rect 37004 18634 37056 18640
rect 37016 18222 37044 18634
rect 37292 18630 37320 18822
rect 37464 18760 37516 18766
rect 37464 18702 37516 18708
rect 37280 18624 37332 18630
rect 37280 18566 37332 18572
rect 37372 18624 37424 18630
rect 37372 18566 37424 18572
rect 37280 18420 37332 18426
rect 37280 18362 37332 18368
rect 37004 18216 37056 18222
rect 37004 18158 37056 18164
rect 37292 17814 37320 18362
rect 37384 18154 37412 18566
rect 37476 18222 37504 18702
rect 37568 18426 37596 20538
rect 37660 20534 37688 21490
rect 37648 20528 37700 20534
rect 37648 20470 37700 20476
rect 37648 19508 37700 19514
rect 37648 19450 37700 19456
rect 37660 19417 37688 19450
rect 37646 19408 37702 19417
rect 37646 19343 37702 19352
rect 37752 18970 37780 22646
rect 37832 22500 37884 22506
rect 37832 22442 37884 22448
rect 37844 21434 37872 22442
rect 37936 21894 37964 24754
rect 38120 22710 38148 25842
rect 38752 25764 38804 25770
rect 38752 25706 38804 25712
rect 38200 25288 38252 25294
rect 38200 25230 38252 25236
rect 38212 24954 38240 25230
rect 38200 24948 38252 24954
rect 38200 24890 38252 24896
rect 38764 24818 38792 25706
rect 38752 24812 38804 24818
rect 38752 24754 38804 24760
rect 38200 24336 38252 24342
rect 38200 24278 38252 24284
rect 38212 24070 38240 24278
rect 38856 24206 38884 29446
rect 39028 28552 39080 28558
rect 39028 28494 39080 28500
rect 38936 26784 38988 26790
rect 38936 26726 38988 26732
rect 38948 24614 38976 26726
rect 38936 24608 38988 24614
rect 38936 24550 38988 24556
rect 38844 24200 38896 24206
rect 38844 24142 38896 24148
rect 38200 24064 38252 24070
rect 38200 24006 38252 24012
rect 38212 23866 38240 24006
rect 38200 23860 38252 23866
rect 38200 23802 38252 23808
rect 38476 23588 38528 23594
rect 38476 23530 38528 23536
rect 38384 22772 38436 22778
rect 38384 22714 38436 22720
rect 38108 22704 38160 22710
rect 38108 22646 38160 22652
rect 38200 22704 38252 22710
rect 38396 22681 38424 22714
rect 38200 22646 38252 22652
rect 38382 22672 38438 22681
rect 38212 22234 38240 22646
rect 38292 22636 38344 22642
rect 38382 22607 38438 22616
rect 38292 22578 38344 22584
rect 38200 22228 38252 22234
rect 38200 22170 38252 22176
rect 38304 21894 38332 22578
rect 38382 22536 38438 22545
rect 38488 22522 38516 23530
rect 38752 22636 38804 22642
rect 38752 22578 38804 22584
rect 38438 22494 38516 22522
rect 38660 22568 38712 22574
rect 38660 22510 38712 22516
rect 38382 22471 38438 22480
rect 37924 21888 37976 21894
rect 37924 21830 37976 21836
rect 38292 21888 38344 21894
rect 38292 21830 38344 21836
rect 37844 21406 38056 21434
rect 37832 21344 37884 21350
rect 37832 21286 37884 21292
rect 37740 18964 37792 18970
rect 37740 18906 37792 18912
rect 37752 18850 37780 18906
rect 37660 18822 37780 18850
rect 37660 18766 37688 18822
rect 37844 18766 37872 21286
rect 37924 19780 37976 19786
rect 37924 19722 37976 19728
rect 37936 19446 37964 19722
rect 38028 19514 38056 21406
rect 38304 21078 38332 21830
rect 38292 21072 38344 21078
rect 38292 21014 38344 21020
rect 38200 20528 38252 20534
rect 38200 20470 38252 20476
rect 38212 19718 38240 20470
rect 38200 19712 38252 19718
rect 38200 19654 38252 19660
rect 38290 19544 38346 19553
rect 38016 19508 38068 19514
rect 38396 19514 38424 22471
rect 38672 21894 38700 22510
rect 38660 21888 38712 21894
rect 38660 21830 38712 21836
rect 38764 21690 38792 22578
rect 38948 22409 38976 24550
rect 38934 22400 38990 22409
rect 38934 22335 38990 22344
rect 38752 21684 38804 21690
rect 38752 21626 38804 21632
rect 38660 21344 38712 21350
rect 38660 21286 38712 21292
rect 38568 21004 38620 21010
rect 38568 20946 38620 20952
rect 38476 19712 38528 19718
rect 38476 19654 38528 19660
rect 38488 19514 38516 19654
rect 38290 19479 38292 19488
rect 38016 19450 38068 19456
rect 38344 19479 38346 19488
rect 38384 19508 38436 19514
rect 38292 19450 38344 19456
rect 38384 19450 38436 19456
rect 38476 19508 38528 19514
rect 38476 19450 38528 19456
rect 37924 19440 37976 19446
rect 37924 19382 37976 19388
rect 38016 19372 38068 19378
rect 38016 19314 38068 19320
rect 37648 18760 37700 18766
rect 37648 18702 37700 18708
rect 37832 18760 37884 18766
rect 37832 18702 37884 18708
rect 37556 18420 37608 18426
rect 37556 18362 37608 18368
rect 37464 18216 37516 18222
rect 37464 18158 37516 18164
rect 37372 18148 37424 18154
rect 37372 18090 37424 18096
rect 37280 17808 37332 17814
rect 37280 17750 37332 17756
rect 37476 17746 37504 18158
rect 37568 17882 37596 18362
rect 37844 18358 37872 18702
rect 37832 18352 37884 18358
rect 37832 18294 37884 18300
rect 37740 18284 37792 18290
rect 37740 18226 37792 18232
rect 37556 17876 37608 17882
rect 37556 17818 37608 17824
rect 37464 17740 37516 17746
rect 37464 17682 37516 17688
rect 37372 17672 37424 17678
rect 37372 17614 37424 17620
rect 37384 17542 37412 17614
rect 37280 17536 37332 17542
rect 37280 17478 37332 17484
rect 37372 17536 37424 17542
rect 37372 17478 37424 17484
rect 37004 17196 37056 17202
rect 37004 17138 37056 17144
rect 36832 16646 36952 16674
rect 36648 14470 36768 14498
rect 36832 14482 36860 16646
rect 37016 16402 37044 17138
rect 37292 16998 37320 17478
rect 37280 16992 37332 16998
rect 37280 16934 37332 16940
rect 37096 16448 37148 16454
rect 37016 16396 37096 16402
rect 37016 16390 37148 16396
rect 37016 16374 37136 16390
rect 37016 16046 37044 16374
rect 37004 16040 37056 16046
rect 37004 15982 37056 15988
rect 37384 15638 37412 17478
rect 37568 16726 37596 17818
rect 37556 16720 37608 16726
rect 37556 16662 37608 16668
rect 37372 15632 37424 15638
rect 37372 15574 37424 15580
rect 37004 15496 37056 15502
rect 37004 15438 37056 15444
rect 37752 15450 37780 18226
rect 37924 15496 37976 15502
rect 37016 14822 37044 15438
rect 37280 15428 37332 15434
rect 37280 15370 37332 15376
rect 37648 15428 37700 15434
rect 37752 15422 37872 15450
rect 37924 15438 37976 15444
rect 37648 15370 37700 15376
rect 37004 14816 37056 14822
rect 37004 14758 37056 14764
rect 36636 14408 36688 14414
rect 36634 14376 36636 14385
rect 36688 14376 36690 14385
rect 36360 14340 36412 14346
rect 36360 14282 36412 14288
rect 36544 14340 36596 14346
rect 36634 14311 36690 14320
rect 36544 14282 36596 14288
rect 36372 14006 36400 14282
rect 36268 14000 36320 14006
rect 36268 13942 36320 13948
rect 36360 14000 36412 14006
rect 36360 13942 36412 13948
rect 35992 13932 36044 13938
rect 35992 13874 36044 13880
rect 35440 13252 35492 13258
rect 35440 13194 35492 13200
rect 35452 12442 35480 13194
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 35716 12708 35768 12714
rect 35716 12650 35768 12656
rect 35440 12436 35492 12442
rect 35440 12378 35492 12384
rect 35728 12374 35756 12650
rect 36004 12442 36032 13874
rect 36280 13802 36308 13942
rect 36452 13932 36504 13938
rect 36452 13874 36504 13880
rect 36268 13796 36320 13802
rect 36268 13738 36320 13744
rect 35992 12436 36044 12442
rect 35992 12378 36044 12384
rect 35716 12368 35768 12374
rect 35716 12310 35768 12316
rect 35348 12300 35400 12306
rect 35348 12242 35400 12248
rect 36004 12170 36032 12378
rect 35992 12164 36044 12170
rect 35992 12106 36044 12112
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 34796 11892 34848 11898
rect 34796 11834 34848 11840
rect 34440 11762 34560 11778
rect 34440 11756 34572 11762
rect 34440 11750 34520 11756
rect 34440 11558 34468 11750
rect 34520 11698 34572 11704
rect 34428 11552 34480 11558
rect 34428 11494 34480 11500
rect 34440 11218 34468 11494
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34428 11212 34480 11218
rect 34428 11154 34480 11160
rect 35992 11076 36044 11082
rect 35992 11018 36044 11024
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 36004 10810 36032 11018
rect 35992 10804 36044 10810
rect 35992 10746 36044 10752
rect 34428 10736 34480 10742
rect 34428 10678 34480 10684
rect 34336 9920 34388 9926
rect 34336 9862 34388 9868
rect 34334 9616 34390 9625
rect 34334 9551 34336 9560
rect 34388 9551 34390 9560
rect 34336 9522 34388 9528
rect 34244 9512 34296 9518
rect 34164 9472 34244 9500
rect 34244 9454 34296 9460
rect 34072 9302 34192 9330
rect 33968 8832 34020 8838
rect 33968 8774 34020 8780
rect 32956 8424 33008 8430
rect 32956 8366 33008 8372
rect 33232 8424 33284 8430
rect 33232 8366 33284 8372
rect 33692 8424 33744 8430
rect 33692 8366 33744 8372
rect 33876 8424 33928 8430
rect 33876 8366 33928 8372
rect 32772 8356 32824 8362
rect 32772 8298 32824 8304
rect 32588 7812 32640 7818
rect 32588 7754 32640 7760
rect 32784 7410 32812 8298
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 32968 6322 32996 8366
rect 33704 7410 33732 8366
rect 33692 7404 33744 7410
rect 33692 7346 33744 7352
rect 33876 7404 33928 7410
rect 33876 7346 33928 7352
rect 33048 7336 33100 7342
rect 33048 7278 33100 7284
rect 33060 6662 33088 7278
rect 33416 6996 33468 7002
rect 33416 6938 33468 6944
rect 33324 6860 33376 6866
rect 33324 6802 33376 6808
rect 33336 6662 33364 6802
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 32956 6316 33008 6322
rect 32956 6258 33008 6264
rect 32968 6118 32996 6258
rect 32956 6112 33008 6118
rect 32956 6054 33008 6060
rect 32036 5840 32088 5846
rect 32036 5782 32088 5788
rect 32048 5234 32076 5782
rect 33060 5778 33088 6598
rect 33324 6316 33376 6322
rect 33428 6304 33456 6938
rect 33704 6866 33732 7346
rect 33692 6860 33744 6866
rect 33692 6802 33744 6808
rect 33600 6724 33652 6730
rect 33600 6666 33652 6672
rect 33508 6452 33560 6458
rect 33508 6394 33560 6400
rect 33520 6322 33548 6394
rect 33376 6276 33456 6304
rect 33508 6316 33560 6322
rect 33324 6258 33376 6264
rect 33508 6258 33560 6264
rect 33048 5772 33100 5778
rect 33048 5714 33100 5720
rect 33336 5642 33364 6258
rect 33520 5710 33548 6258
rect 33508 5704 33560 5710
rect 33508 5646 33560 5652
rect 33324 5636 33376 5642
rect 33324 5578 33376 5584
rect 33140 5568 33192 5574
rect 33140 5510 33192 5516
rect 33152 5234 33180 5510
rect 32036 5228 32088 5234
rect 32036 5170 32088 5176
rect 33140 5228 33192 5234
rect 33140 5170 33192 5176
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 32324 4690 32352 4966
rect 32312 4684 32364 4690
rect 32312 4626 32364 4632
rect 33612 4554 33640 6666
rect 33704 5302 33732 6802
rect 33888 6458 33916 7346
rect 33980 6730 34008 8774
rect 34060 7200 34112 7206
rect 34060 7142 34112 7148
rect 34072 7002 34100 7142
rect 34060 6996 34112 7002
rect 34060 6938 34112 6944
rect 33968 6724 34020 6730
rect 33968 6666 34020 6672
rect 34164 6644 34192 9302
rect 34440 8906 34468 10678
rect 34888 10600 34940 10606
rect 34808 10548 34888 10554
rect 34808 10542 34940 10548
rect 34808 10526 34928 10542
rect 34612 10464 34664 10470
rect 34612 10406 34664 10412
rect 34624 10130 34652 10406
rect 34612 10124 34664 10130
rect 34612 10066 34664 10072
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34532 9353 34560 9998
rect 34808 9994 34836 10526
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 9988 34848 9994
rect 34796 9930 34848 9936
rect 34704 9920 34756 9926
rect 34704 9862 34756 9868
rect 34716 9654 34744 9862
rect 34704 9648 34756 9654
rect 34704 9590 34756 9596
rect 34808 9586 34836 9930
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 35716 9648 35768 9654
rect 35714 9616 35716 9625
rect 35768 9616 35770 9625
rect 34796 9580 34848 9586
rect 34796 9522 34848 9528
rect 35256 9580 35308 9586
rect 35714 9551 35770 9560
rect 35256 9522 35308 9528
rect 34612 9512 34664 9518
rect 34612 9454 34664 9460
rect 35268 9466 35296 9522
rect 35900 9512 35952 9518
rect 34518 9344 34574 9353
rect 34518 9279 34574 9288
rect 34624 9081 34652 9454
rect 35268 9438 35388 9466
rect 35900 9454 35952 9460
rect 35990 9480 36046 9489
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34610 9072 34666 9081
rect 34610 9007 34666 9016
rect 35164 9036 35216 9042
rect 35164 8978 35216 8984
rect 34428 8900 34480 8906
rect 34428 8842 34480 8848
rect 34704 8832 34756 8838
rect 34704 8774 34756 8780
rect 34716 8498 34744 8774
rect 35176 8498 35204 8978
rect 35360 8634 35388 9438
rect 35912 9382 35940 9454
rect 35990 9415 36046 9424
rect 36176 9444 36228 9450
rect 35440 9376 35492 9382
rect 35900 9376 35952 9382
rect 35440 9318 35492 9324
rect 35898 9344 35900 9353
rect 35952 9344 35954 9353
rect 35452 8634 35480 9318
rect 35898 9279 35954 9288
rect 36004 9110 36032 9415
rect 36176 9386 36228 9392
rect 35992 9104 36044 9110
rect 35992 9046 36044 9052
rect 35900 8968 35952 8974
rect 35952 8928 36032 8956
rect 35900 8910 35952 8916
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 35348 8628 35400 8634
rect 35348 8570 35400 8576
rect 35440 8628 35492 8634
rect 35440 8570 35492 8576
rect 35532 8628 35584 8634
rect 35532 8570 35584 8576
rect 35544 8537 35572 8570
rect 35530 8528 35586 8537
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 35164 8492 35216 8498
rect 35440 8492 35492 8498
rect 35164 8434 35216 8440
rect 35360 8452 35440 8480
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34428 7880 34480 7886
rect 34428 7822 34480 7828
rect 34244 6656 34296 6662
rect 34164 6616 34244 6644
rect 34244 6598 34296 6604
rect 33876 6452 33928 6458
rect 33876 6394 33928 6400
rect 34152 6112 34204 6118
rect 34152 6054 34204 6060
rect 34164 5710 34192 6054
rect 34256 5914 34284 6598
rect 34440 6254 34468 7822
rect 34704 7812 34756 7818
rect 34704 7754 34756 7760
rect 34428 6248 34480 6254
rect 34428 6190 34480 6196
rect 34244 5908 34296 5914
rect 34244 5850 34296 5856
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 34152 5704 34204 5710
rect 34152 5646 34204 5652
rect 33692 5296 33744 5302
rect 33692 5238 33744 5244
rect 33704 4604 33732 5238
rect 34072 4690 34100 5646
rect 34440 5302 34468 6190
rect 34612 5704 34664 5710
rect 34716 5692 34744 7754
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35360 6882 35388 8452
rect 35530 8463 35586 8472
rect 35716 8492 35768 8498
rect 35440 8434 35492 8440
rect 35768 8452 35940 8480
rect 35716 8434 35768 8440
rect 35440 8356 35492 8362
rect 35440 8298 35492 8304
rect 35452 8090 35480 8298
rect 35440 8084 35492 8090
rect 35440 8026 35492 8032
rect 35912 7954 35940 8452
rect 35900 7948 35952 7954
rect 35900 7890 35952 7896
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 35360 6854 35480 6882
rect 34796 6792 34848 6798
rect 34796 6734 34848 6740
rect 35348 6792 35400 6798
rect 35348 6734 35400 6740
rect 34808 6322 34836 6734
rect 35164 6724 35216 6730
rect 35164 6666 35216 6672
rect 35072 6656 35124 6662
rect 35072 6598 35124 6604
rect 35084 6390 35112 6598
rect 35176 6390 35204 6666
rect 35072 6384 35124 6390
rect 35072 6326 35124 6332
rect 35164 6384 35216 6390
rect 35164 6326 35216 6332
rect 34796 6316 34848 6322
rect 34796 6258 34848 6264
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35360 5914 35388 6734
rect 35348 5908 35400 5914
rect 35348 5850 35400 5856
rect 34796 5704 34848 5710
rect 34716 5664 34796 5692
rect 34612 5646 34664 5652
rect 34796 5646 34848 5652
rect 35164 5704 35216 5710
rect 35164 5646 35216 5652
rect 34520 5636 34572 5642
rect 34520 5578 34572 5584
rect 34532 5386 34560 5578
rect 34624 5574 34652 5646
rect 34888 5636 34940 5642
rect 34888 5578 34940 5584
rect 34612 5568 34664 5574
rect 34612 5510 34664 5516
rect 34900 5386 34928 5578
rect 34532 5358 34928 5386
rect 34428 5296 34480 5302
rect 34428 5238 34480 5244
rect 34440 4758 34468 5238
rect 34900 5234 34928 5358
rect 35176 5234 35204 5646
rect 35452 5642 35480 6854
rect 36004 6662 36032 8928
rect 36188 8906 36216 9386
rect 36280 9382 36308 13738
rect 36360 13320 36412 13326
rect 36360 13262 36412 13268
rect 36372 12918 36400 13262
rect 36360 12912 36412 12918
rect 36360 12854 36412 12860
rect 36372 12646 36400 12854
rect 36360 12640 36412 12646
rect 36360 12582 36412 12588
rect 36464 12434 36492 13874
rect 36556 13870 36584 14282
rect 36544 13864 36596 13870
rect 36544 13806 36596 13812
rect 36636 13728 36688 13734
rect 36636 13670 36688 13676
rect 36648 13530 36676 13670
rect 36636 13524 36688 13530
rect 36636 13466 36688 13472
rect 36740 13326 36768 14470
rect 36820 14476 36872 14482
rect 36820 14418 36872 14424
rect 36910 14376 36966 14385
rect 37016 14346 37044 14758
rect 37292 14482 37320 15370
rect 37660 15162 37688 15370
rect 37740 15360 37792 15366
rect 37740 15302 37792 15308
rect 37648 15156 37700 15162
rect 37648 15098 37700 15104
rect 37660 14498 37688 15098
rect 37752 15094 37780 15302
rect 37740 15088 37792 15094
rect 37740 15030 37792 15036
rect 37568 14482 37688 14498
rect 37188 14476 37240 14482
rect 37188 14418 37240 14424
rect 37280 14476 37332 14482
rect 37280 14418 37332 14424
rect 37556 14476 37688 14482
rect 37608 14470 37688 14476
rect 37556 14418 37608 14424
rect 36910 14311 36966 14320
rect 37004 14340 37056 14346
rect 36924 14278 36952 14311
rect 37004 14282 37056 14288
rect 36820 14272 36872 14278
rect 36820 14214 36872 14220
rect 36912 14272 36964 14278
rect 36912 14214 36964 14220
rect 36832 13462 36860 14214
rect 36820 13456 36872 13462
rect 36820 13398 36872 13404
rect 36728 13320 36780 13326
rect 36728 13262 36780 13268
rect 37004 13320 37056 13326
rect 37004 13262 37056 13268
rect 36544 13184 36596 13190
rect 36544 13126 36596 13132
rect 36372 12406 36492 12434
rect 36268 9376 36320 9382
rect 36372 9353 36400 12406
rect 36556 11898 36584 13126
rect 36636 12368 36688 12374
rect 36636 12310 36688 12316
rect 36544 11892 36596 11898
rect 36544 11834 36596 11840
rect 36556 11694 36584 11834
rect 36648 11762 36676 12310
rect 36636 11756 36688 11762
rect 36636 11698 36688 11704
rect 36544 11688 36596 11694
rect 36544 11630 36596 11636
rect 36544 11552 36596 11558
rect 36544 11494 36596 11500
rect 36556 10674 36584 11494
rect 36544 10668 36596 10674
rect 36544 10610 36596 10616
rect 36636 9512 36688 9518
rect 36636 9454 36688 9460
rect 36268 9318 36320 9324
rect 36358 9344 36414 9353
rect 36176 8900 36228 8906
rect 36176 8842 36228 8848
rect 36280 8498 36308 9318
rect 36358 9279 36414 9288
rect 36648 8974 36676 9454
rect 36360 8968 36412 8974
rect 36360 8910 36412 8916
rect 36636 8968 36688 8974
rect 36636 8910 36688 8916
rect 36740 8922 36768 13262
rect 37016 12986 37044 13262
rect 37096 13252 37148 13258
rect 37096 13194 37148 13200
rect 36912 12980 36964 12986
rect 36912 12922 36964 12928
rect 37004 12980 37056 12986
rect 37004 12922 37056 12928
rect 36820 12844 36872 12850
rect 36820 12786 36872 12792
rect 36832 9042 36860 12786
rect 36924 11762 36952 12922
rect 37108 12850 37136 13194
rect 37096 12844 37148 12850
rect 37096 12786 37148 12792
rect 37096 11892 37148 11898
rect 37096 11834 37148 11840
rect 36912 11756 36964 11762
rect 36912 11698 36964 11704
rect 37108 11626 37136 11834
rect 37096 11620 37148 11626
rect 37096 11562 37148 11568
rect 37004 9104 37056 9110
rect 37004 9046 37056 9052
rect 36820 9036 36872 9042
rect 36820 8978 36872 8984
rect 36372 8673 36400 8910
rect 36740 8894 36860 8922
rect 36544 8832 36596 8838
rect 36544 8774 36596 8780
rect 36636 8832 36688 8838
rect 36636 8774 36688 8780
rect 36358 8664 36414 8673
rect 36556 8634 36584 8774
rect 36358 8599 36414 8608
rect 36544 8628 36596 8634
rect 36544 8570 36596 8576
rect 36176 8492 36228 8498
rect 36176 8434 36228 8440
rect 36268 8492 36320 8498
rect 36268 8434 36320 8440
rect 36082 8392 36138 8401
rect 36082 8327 36138 8336
rect 36096 8294 36124 8327
rect 36084 8288 36136 8294
rect 36084 8230 36136 8236
rect 36096 8022 36124 8230
rect 36084 8016 36136 8022
rect 36084 7958 36136 7964
rect 35992 6656 36044 6662
rect 35992 6598 36044 6604
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 36084 6112 36136 6118
rect 36084 6054 36136 6060
rect 35992 5840 36044 5846
rect 35992 5782 36044 5788
rect 35440 5636 35492 5642
rect 35440 5578 35492 5584
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 34888 5228 34940 5234
rect 34888 5170 34940 5176
rect 35164 5228 35216 5234
rect 35164 5170 35216 5176
rect 36004 5098 36032 5782
rect 36096 5778 36124 6054
rect 36188 5930 36216 8434
rect 36280 8022 36308 8434
rect 36268 8016 36320 8022
rect 36268 7958 36320 7964
rect 36648 6882 36676 8774
rect 36726 8664 36782 8673
rect 36726 8599 36782 8608
rect 36740 8566 36768 8599
rect 36728 8560 36780 8566
rect 36728 8502 36780 8508
rect 36464 6854 36676 6882
rect 36188 5902 36308 5930
rect 36176 5840 36228 5846
rect 36176 5782 36228 5788
rect 36084 5772 36136 5778
rect 36084 5714 36136 5720
rect 35992 5092 36044 5098
rect 35992 5034 36044 5040
rect 35532 5024 35584 5030
rect 35532 4966 35584 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34428 4752 34480 4758
rect 34428 4694 34480 4700
rect 34060 4684 34112 4690
rect 34060 4626 34112 4632
rect 33784 4616 33836 4622
rect 33704 4576 33784 4604
rect 33784 4558 33836 4564
rect 33600 4548 33652 4554
rect 33600 4490 33652 4496
rect 33612 4214 33640 4490
rect 31864 4134 31984 4162
rect 33600 4208 33652 4214
rect 33600 4150 33652 4156
rect 31864 3942 31892 4134
rect 34072 4078 34100 4626
rect 35544 4622 35572 4966
rect 35532 4616 35584 4622
rect 35532 4558 35584 4564
rect 36096 4554 36124 5714
rect 36188 5234 36216 5782
rect 36280 5370 36308 5902
rect 36268 5364 36320 5370
rect 36268 5306 36320 5312
rect 36176 5228 36228 5234
rect 36176 5170 36228 5176
rect 36360 5228 36412 5234
rect 36464 5216 36492 6854
rect 36636 6792 36688 6798
rect 36636 6734 36688 6740
rect 36648 6458 36676 6734
rect 36832 6644 36860 8894
rect 37016 8242 37044 9046
rect 37200 8566 37228 14418
rect 37292 12238 37320 14418
rect 37464 12912 37516 12918
rect 37462 12880 37464 12889
rect 37516 12880 37518 12889
rect 37462 12815 37518 12824
rect 37372 12368 37424 12374
rect 37372 12310 37424 12316
rect 37280 12232 37332 12238
rect 37280 12174 37332 12180
rect 37280 11688 37332 11694
rect 37280 11630 37332 11636
rect 37292 10674 37320 11630
rect 37280 10668 37332 10674
rect 37280 10610 37332 10616
rect 37280 9920 37332 9926
rect 37280 9862 37332 9868
rect 37292 9518 37320 9862
rect 37280 9512 37332 9518
rect 37280 9454 37332 9460
rect 37280 9104 37332 9110
rect 37280 9046 37332 9052
rect 37292 8566 37320 9046
rect 37188 8560 37240 8566
rect 37188 8502 37240 8508
rect 37280 8560 37332 8566
rect 37280 8502 37332 8508
rect 37200 8430 37228 8502
rect 37188 8424 37240 8430
rect 37188 8366 37240 8372
rect 37280 8424 37332 8430
rect 37280 8366 37332 8372
rect 37292 8242 37320 8366
rect 37384 8294 37412 12310
rect 37568 12306 37596 14418
rect 37740 14272 37792 14278
rect 37740 14214 37792 14220
rect 37752 12918 37780 14214
rect 37844 13530 37872 15422
rect 37936 14618 37964 15438
rect 37924 14612 37976 14618
rect 37924 14554 37976 14560
rect 37832 13524 37884 13530
rect 37832 13466 37884 13472
rect 37832 13320 37884 13326
rect 37832 13262 37884 13268
rect 37844 12986 37872 13262
rect 38028 13258 38056 19314
rect 38304 19310 38332 19450
rect 38292 19304 38344 19310
rect 38292 19246 38344 19252
rect 38200 19168 38252 19174
rect 38200 19110 38252 19116
rect 38384 19168 38436 19174
rect 38384 19110 38436 19116
rect 38212 18970 38240 19110
rect 38108 18964 38160 18970
rect 38108 18906 38160 18912
rect 38200 18964 38252 18970
rect 38200 18906 38252 18912
rect 38120 18850 38148 18906
rect 38292 18896 38344 18902
rect 38120 18844 38292 18850
rect 38120 18838 38344 18844
rect 38120 18822 38332 18838
rect 38108 18352 38160 18358
rect 38108 18294 38160 18300
rect 38016 13252 38068 13258
rect 38016 13194 38068 13200
rect 37832 12980 37884 12986
rect 37832 12922 37884 12928
rect 37924 12980 37976 12986
rect 37924 12922 37976 12928
rect 37740 12912 37792 12918
rect 37740 12854 37792 12860
rect 37648 12844 37700 12850
rect 37648 12786 37700 12792
rect 37556 12300 37608 12306
rect 37556 12242 37608 12248
rect 37464 11892 37516 11898
rect 37464 11834 37516 11840
rect 37476 11014 37504 11834
rect 37568 11830 37596 12242
rect 37556 11824 37608 11830
rect 37556 11766 37608 11772
rect 37660 11336 37688 12786
rect 37936 12434 37964 12922
rect 38120 12918 38148 18294
rect 38292 18148 38344 18154
rect 38292 18090 38344 18096
rect 38198 17640 38254 17649
rect 38198 17575 38200 17584
rect 38252 17575 38254 17584
rect 38200 17546 38252 17552
rect 38200 16788 38252 16794
rect 38200 16730 38252 16736
rect 38212 16250 38240 16730
rect 38200 16244 38252 16250
rect 38200 16186 38252 16192
rect 38200 13320 38252 13326
rect 38200 13262 38252 13268
rect 38108 12912 38160 12918
rect 38108 12854 38160 12860
rect 38212 12714 38240 13262
rect 38304 13190 38332 18090
rect 38396 18086 38424 19110
rect 38384 18080 38436 18086
rect 38382 18048 38384 18057
rect 38436 18048 38438 18057
rect 38382 17983 38438 17992
rect 38488 17814 38516 19450
rect 38476 17808 38528 17814
rect 38476 17750 38528 17756
rect 38384 17196 38436 17202
rect 38384 17138 38436 17144
rect 38396 16794 38424 17138
rect 38384 16788 38436 16794
rect 38384 16730 38436 16736
rect 38488 16726 38516 17750
rect 38580 17746 38608 20946
rect 38672 20942 38700 21286
rect 38660 20936 38712 20942
rect 38660 20878 38712 20884
rect 38936 20936 38988 20942
rect 38936 20878 38988 20884
rect 38948 19922 38976 20878
rect 38936 19916 38988 19922
rect 38936 19858 38988 19864
rect 38844 19712 38896 19718
rect 38844 19654 38896 19660
rect 38752 19304 38804 19310
rect 38752 19246 38804 19252
rect 38764 18970 38792 19246
rect 38752 18964 38804 18970
rect 38752 18906 38804 18912
rect 38856 18766 38884 19654
rect 38936 19372 38988 19378
rect 38936 19314 38988 19320
rect 38844 18760 38896 18766
rect 38844 18702 38896 18708
rect 38752 18080 38804 18086
rect 38752 18022 38804 18028
rect 38568 17740 38620 17746
rect 38568 17682 38620 17688
rect 38580 17202 38608 17682
rect 38764 17270 38792 18022
rect 38844 17876 38896 17882
rect 38844 17818 38896 17824
rect 38752 17264 38804 17270
rect 38752 17206 38804 17212
rect 38568 17196 38620 17202
rect 38568 17138 38620 17144
rect 38476 16720 38528 16726
rect 38476 16662 38528 16668
rect 38752 15700 38804 15706
rect 38752 15642 38804 15648
rect 38568 15564 38620 15570
rect 38568 15506 38620 15512
rect 38384 13524 38436 13530
rect 38384 13466 38436 13472
rect 38396 13326 38424 13466
rect 38384 13320 38436 13326
rect 38384 13262 38436 13268
rect 38292 13184 38344 13190
rect 38292 13126 38344 13132
rect 38304 12986 38332 13126
rect 38292 12980 38344 12986
rect 38292 12922 38344 12928
rect 38290 12880 38346 12889
rect 38290 12815 38292 12824
rect 38344 12815 38346 12824
rect 38292 12786 38344 12792
rect 38200 12708 38252 12714
rect 38200 12650 38252 12656
rect 38212 12434 38240 12650
rect 38396 12434 38424 13262
rect 38580 12850 38608 15506
rect 38568 12844 38620 12850
rect 38568 12786 38620 12792
rect 37936 12406 38056 12434
rect 37832 12232 37884 12238
rect 37832 12174 37884 12180
rect 37844 11762 37872 12174
rect 37832 11756 37884 11762
rect 37832 11698 37884 11704
rect 37568 11308 37688 11336
rect 37464 11008 37516 11014
rect 37464 10950 37516 10956
rect 37568 9625 37596 11308
rect 37844 11286 37872 11698
rect 37832 11280 37884 11286
rect 37832 11222 37884 11228
rect 37648 11212 37700 11218
rect 37648 11154 37700 11160
rect 37660 10606 37688 11154
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 37648 10600 37700 10606
rect 37648 10542 37700 10548
rect 37554 9616 37610 9625
rect 37660 9586 37688 10542
rect 37554 9551 37610 9560
rect 37648 9580 37700 9586
rect 37648 9522 37700 9528
rect 37464 9444 37516 9450
rect 37464 9386 37516 9392
rect 37476 9042 37504 9386
rect 37464 9036 37516 9042
rect 37464 8978 37516 8984
rect 37476 8362 37504 8978
rect 37648 8900 37700 8906
rect 37648 8842 37700 8848
rect 37556 8628 37608 8634
rect 37556 8570 37608 8576
rect 37568 8498 37596 8570
rect 37660 8498 37688 8842
rect 37556 8492 37608 8498
rect 37556 8434 37608 8440
rect 37648 8492 37700 8498
rect 37648 8434 37700 8440
rect 37464 8356 37516 8362
rect 37464 8298 37516 8304
rect 37016 8214 37320 8242
rect 37372 8288 37424 8294
rect 37372 8230 37424 8236
rect 36912 6656 36964 6662
rect 36832 6616 36912 6644
rect 36912 6598 36964 6604
rect 36636 6452 36688 6458
rect 36636 6394 36688 6400
rect 37016 6338 37044 8214
rect 37660 7954 37688 8434
rect 37280 7948 37332 7954
rect 37280 7890 37332 7896
rect 37648 7948 37700 7954
rect 37648 7890 37700 7896
rect 37292 7546 37320 7890
rect 37280 7540 37332 7546
rect 37280 7482 37332 7488
rect 37372 7472 37424 7478
rect 37372 7414 37424 7420
rect 37384 6934 37412 7414
rect 37372 6928 37424 6934
rect 37844 6905 37872 10610
rect 37924 9512 37976 9518
rect 37924 9454 37976 9460
rect 37936 9178 37964 9454
rect 37924 9172 37976 9178
rect 37924 9114 37976 9120
rect 38028 9042 38056 12406
rect 38120 12406 38240 12434
rect 38304 12406 38424 12434
rect 38120 12238 38148 12406
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 38108 12096 38160 12102
rect 38108 12038 38160 12044
rect 38120 11558 38148 12038
rect 38108 11552 38160 11558
rect 38108 11494 38160 11500
rect 38200 11552 38252 11558
rect 38200 11494 38252 11500
rect 38016 9036 38068 9042
rect 38016 8978 38068 8984
rect 38120 8566 38148 11494
rect 38212 11218 38240 11494
rect 38200 11212 38252 11218
rect 38200 11154 38252 11160
rect 38200 9648 38252 9654
rect 38200 9590 38252 9596
rect 38212 8786 38240 9590
rect 38304 8974 38332 12406
rect 38476 12232 38528 12238
rect 38476 12174 38528 12180
rect 38384 12096 38436 12102
rect 38384 12038 38436 12044
rect 38396 11762 38424 12038
rect 38488 11830 38516 12174
rect 38476 11824 38528 11830
rect 38476 11766 38528 11772
rect 38384 11756 38436 11762
rect 38384 11698 38436 11704
rect 38580 11558 38608 12786
rect 38568 11552 38620 11558
rect 38568 11494 38620 11500
rect 38580 10742 38608 11494
rect 38660 11076 38712 11082
rect 38660 11018 38712 11024
rect 38672 10742 38700 11018
rect 38568 10736 38620 10742
rect 38568 10678 38620 10684
rect 38660 10736 38712 10742
rect 38660 10678 38712 10684
rect 38672 9674 38700 10678
rect 38764 10674 38792 15642
rect 38856 13938 38884 17818
rect 38948 17134 38976 19314
rect 39040 19310 39068 28494
rect 39212 27396 39264 27402
rect 39212 27338 39264 27344
rect 39224 27062 39252 27338
rect 39212 27056 39264 27062
rect 39212 26998 39264 27004
rect 39224 25226 39252 26998
rect 39212 25220 39264 25226
rect 39212 25162 39264 25168
rect 39120 24064 39172 24070
rect 39120 24006 39172 24012
rect 39132 23730 39160 24006
rect 39224 23866 39252 25162
rect 39212 23860 39264 23866
rect 39212 23802 39264 23808
rect 39120 23724 39172 23730
rect 39120 23666 39172 23672
rect 39120 23112 39172 23118
rect 39120 23054 39172 23060
rect 39132 22778 39160 23054
rect 39120 22772 39172 22778
rect 39120 22714 39172 22720
rect 39212 22704 39264 22710
rect 39212 22646 39264 22652
rect 39224 22522 39252 22646
rect 39132 22494 39252 22522
rect 39132 19394 39160 22494
rect 39316 22488 39344 39200
rect 39396 37188 39448 37194
rect 39396 37130 39448 37136
rect 39408 29306 39436 37130
rect 39960 36922 39988 39200
rect 40500 37256 40552 37262
rect 40500 37198 40552 37204
rect 39948 36916 40000 36922
rect 39948 36858 40000 36864
rect 40408 36848 40460 36854
rect 40408 36790 40460 36796
rect 39488 36576 39540 36582
rect 39488 36518 39540 36524
rect 39500 36106 39528 36518
rect 40420 36106 40448 36790
rect 40512 36786 40540 37198
rect 40604 36922 40632 39200
rect 40868 37256 40920 37262
rect 40868 37198 40920 37204
rect 40592 36916 40644 36922
rect 40592 36858 40644 36864
rect 40880 36786 40908 37198
rect 41248 36922 41276 39200
rect 41892 36922 41920 39200
rect 42536 36922 42564 39200
rect 43180 36922 43208 39200
rect 43824 37398 43852 39200
rect 43812 37392 43864 37398
rect 43812 37334 43864 37340
rect 43904 37188 43956 37194
rect 43904 37130 43956 37136
rect 44364 37188 44416 37194
rect 44364 37130 44416 37136
rect 41236 36916 41288 36922
rect 41236 36858 41288 36864
rect 41880 36916 41932 36922
rect 41880 36858 41932 36864
rect 42524 36916 42576 36922
rect 42524 36858 42576 36864
rect 43168 36916 43220 36922
rect 43168 36858 43220 36864
rect 40500 36780 40552 36786
rect 40500 36722 40552 36728
rect 40868 36780 40920 36786
rect 40868 36722 40920 36728
rect 42524 36780 42576 36786
rect 42524 36722 42576 36728
rect 43076 36780 43128 36786
rect 43076 36722 43128 36728
rect 42248 36712 42300 36718
rect 42248 36654 42300 36660
rect 42260 36242 42288 36654
rect 42536 36378 42564 36722
rect 43088 36378 43116 36722
rect 43536 36712 43588 36718
rect 43536 36654 43588 36660
rect 43548 36378 43576 36654
rect 42524 36372 42576 36378
rect 42524 36314 42576 36320
rect 43076 36372 43128 36378
rect 43076 36314 43128 36320
rect 43536 36372 43588 36378
rect 43536 36314 43588 36320
rect 43720 36372 43772 36378
rect 43720 36314 43772 36320
rect 42248 36236 42300 36242
rect 42248 36178 42300 36184
rect 39488 36100 39540 36106
rect 39488 36042 39540 36048
rect 40408 36100 40460 36106
rect 40408 36042 40460 36048
rect 41972 36100 42024 36106
rect 41972 36042 42024 36048
rect 40420 34610 40448 36042
rect 40684 36032 40736 36038
rect 40684 35974 40736 35980
rect 40696 35698 40724 35974
rect 41984 35834 42012 36042
rect 41972 35828 42024 35834
rect 41972 35770 42024 35776
rect 41328 35760 41380 35766
rect 41328 35702 41380 35708
rect 40684 35692 40736 35698
rect 40684 35634 40736 35640
rect 40868 35692 40920 35698
rect 40868 35634 40920 35640
rect 40408 34604 40460 34610
rect 40408 34546 40460 34552
rect 39488 34400 39540 34406
rect 39488 34342 39540 34348
rect 40040 34400 40092 34406
rect 40040 34342 40092 34348
rect 39500 34202 39528 34342
rect 39488 34196 39540 34202
rect 39488 34138 39540 34144
rect 39948 33992 40000 33998
rect 39948 33934 40000 33940
rect 39960 33658 39988 33934
rect 40052 33930 40080 34342
rect 40040 33924 40092 33930
rect 40040 33866 40092 33872
rect 39948 33652 40000 33658
rect 39948 33594 40000 33600
rect 39488 33584 39540 33590
rect 40052 33538 40080 33866
rect 40696 33862 40724 35634
rect 40880 33998 40908 35634
rect 41236 34604 41288 34610
rect 41236 34546 41288 34552
rect 41144 34196 41196 34202
rect 41144 34138 41196 34144
rect 40960 34060 41012 34066
rect 40960 34002 41012 34008
rect 40868 33992 40920 33998
rect 40868 33934 40920 33940
rect 40684 33856 40736 33862
rect 40684 33798 40736 33804
rect 40696 33674 40724 33798
rect 39488 33526 39540 33532
rect 39500 32910 39528 33526
rect 39868 33510 40080 33538
rect 40604 33646 40724 33674
rect 40880 33658 40908 33934
rect 40868 33652 40920 33658
rect 39868 33318 39896 33510
rect 40604 33318 40632 33646
rect 40868 33594 40920 33600
rect 40684 33584 40736 33590
rect 40684 33526 40736 33532
rect 39672 33312 39724 33318
rect 39672 33254 39724 33260
rect 39856 33312 39908 33318
rect 39856 33254 39908 33260
rect 40592 33312 40644 33318
rect 40592 33254 40644 33260
rect 39488 32904 39540 32910
rect 39488 32846 39540 32852
rect 39684 32774 39712 33254
rect 39868 32978 39896 33254
rect 40696 33114 40724 33526
rect 40684 33108 40736 33114
rect 40684 33050 40736 33056
rect 39856 32972 39908 32978
rect 39856 32914 39908 32920
rect 39672 32768 39724 32774
rect 39672 32710 39724 32716
rect 39948 32768 40000 32774
rect 39948 32710 40000 32716
rect 39684 32366 39712 32710
rect 39672 32360 39724 32366
rect 39672 32302 39724 32308
rect 39960 30394 39988 32710
rect 40684 31884 40736 31890
rect 40684 31826 40736 31832
rect 40500 31680 40552 31686
rect 40500 31622 40552 31628
rect 40512 31414 40540 31622
rect 40696 31482 40724 31826
rect 40880 31482 40908 33594
rect 40972 33522 41000 34002
rect 41052 33992 41104 33998
rect 41052 33934 41104 33940
rect 41064 33658 41092 33934
rect 41052 33652 41104 33658
rect 41052 33594 41104 33600
rect 40960 33516 41012 33522
rect 40960 33458 41012 33464
rect 40684 31476 40736 31482
rect 40604 31436 40684 31464
rect 40500 31408 40552 31414
rect 40500 31350 40552 31356
rect 40604 31142 40632 31436
rect 40684 31418 40736 31424
rect 40868 31476 40920 31482
rect 40868 31418 40920 31424
rect 40684 31272 40736 31278
rect 40684 31214 40736 31220
rect 40592 31136 40644 31142
rect 40592 31078 40644 31084
rect 40696 30938 40724 31214
rect 40972 31210 41000 33458
rect 41156 33318 41184 34138
rect 41144 33312 41196 33318
rect 41144 33254 41196 33260
rect 41248 32910 41276 34546
rect 41340 34490 41368 35702
rect 42260 35630 42288 36178
rect 43732 35766 43760 36314
rect 43720 35760 43772 35766
rect 43720 35702 43772 35708
rect 42248 35624 42300 35630
rect 42248 35566 42300 35572
rect 42260 34610 42288 35566
rect 43732 35222 43760 35702
rect 43720 35216 43772 35222
rect 43720 35158 43772 35164
rect 43352 35080 43404 35086
rect 43352 35022 43404 35028
rect 43536 35080 43588 35086
rect 43536 35022 43588 35028
rect 42800 34944 42852 34950
rect 42800 34886 42852 34892
rect 42812 34678 42840 34886
rect 42800 34672 42852 34678
rect 42800 34614 42852 34620
rect 42248 34604 42300 34610
rect 42248 34546 42300 34552
rect 41340 34462 41460 34490
rect 41328 33992 41380 33998
rect 41328 33934 41380 33940
rect 41340 33522 41368 33934
rect 41328 33516 41380 33522
rect 41328 33458 41380 33464
rect 41236 32904 41288 32910
rect 41236 32846 41288 32852
rect 40960 31204 41012 31210
rect 40960 31146 41012 31152
rect 40776 31136 40828 31142
rect 40776 31078 40828 31084
rect 40684 30932 40736 30938
rect 40684 30874 40736 30880
rect 40592 30728 40644 30734
rect 40592 30670 40644 30676
rect 40224 30660 40276 30666
rect 40224 30602 40276 30608
rect 39948 30388 40000 30394
rect 39948 30330 40000 30336
rect 40236 30326 40264 30602
rect 40224 30320 40276 30326
rect 40224 30262 40276 30268
rect 40236 29510 40264 30262
rect 40604 30190 40632 30670
rect 40788 30326 40816 31078
rect 41248 30666 41276 32846
rect 41432 31822 41460 34462
rect 42156 33924 42208 33930
rect 42156 33866 42208 33872
rect 42168 33522 42196 33866
rect 42156 33516 42208 33522
rect 42156 33458 42208 33464
rect 41604 33380 41656 33386
rect 41604 33322 41656 33328
rect 41616 32774 41644 33322
rect 42168 33318 42196 33458
rect 42156 33312 42208 33318
rect 42156 33254 42208 33260
rect 42260 32978 42288 34546
rect 43364 34202 43392 35022
rect 43352 34196 43404 34202
rect 43352 34138 43404 34144
rect 43548 33998 43576 35022
rect 42432 33992 42484 33998
rect 42432 33934 42484 33940
rect 43536 33992 43588 33998
rect 43536 33934 43588 33940
rect 42444 33522 42472 33934
rect 43812 33652 43864 33658
rect 43812 33594 43864 33600
rect 42432 33516 42484 33522
rect 42432 33458 42484 33464
rect 43824 33114 43852 33594
rect 43812 33108 43864 33114
rect 43812 33050 43864 33056
rect 42248 32972 42300 32978
rect 42248 32914 42300 32920
rect 42708 32972 42760 32978
rect 42708 32914 42760 32920
rect 41604 32768 41656 32774
rect 41604 32710 41656 32716
rect 41420 31816 41472 31822
rect 41420 31758 41472 31764
rect 41696 31816 41748 31822
rect 41696 31758 41748 31764
rect 41708 31346 41736 31758
rect 41696 31340 41748 31346
rect 41696 31282 41748 31288
rect 42524 31340 42576 31346
rect 42524 31282 42576 31288
rect 42536 30938 42564 31282
rect 42524 30932 42576 30938
rect 42524 30874 42576 30880
rect 42720 30802 42748 32914
rect 43824 32434 43852 33050
rect 43812 32428 43864 32434
rect 43812 32370 43864 32376
rect 43536 32292 43588 32298
rect 43536 32234 43588 32240
rect 43548 31754 43576 32234
rect 43824 31822 43852 32370
rect 43812 31816 43864 31822
rect 43812 31758 43864 31764
rect 43548 31726 43668 31754
rect 42892 31408 42944 31414
rect 42892 31350 42944 31356
rect 42800 31136 42852 31142
rect 42800 31078 42852 31084
rect 42708 30796 42760 30802
rect 42708 30738 42760 30744
rect 41236 30660 41288 30666
rect 41236 30602 41288 30608
rect 40776 30320 40828 30326
rect 40776 30262 40828 30268
rect 42812 30258 42840 31078
rect 42904 30258 42932 31350
rect 43076 30660 43128 30666
rect 43076 30602 43128 30608
rect 43088 30394 43116 30602
rect 43640 30598 43668 31726
rect 43628 30592 43680 30598
rect 43628 30534 43680 30540
rect 43076 30388 43128 30394
rect 43076 30330 43128 30336
rect 43640 30258 43668 30534
rect 42800 30252 42852 30258
rect 42800 30194 42852 30200
rect 42892 30252 42944 30258
rect 42892 30194 42944 30200
rect 43628 30252 43680 30258
rect 43628 30194 43680 30200
rect 40592 30184 40644 30190
rect 40592 30126 40644 30132
rect 42432 30184 42484 30190
rect 42432 30126 42484 30132
rect 43444 30184 43496 30190
rect 43444 30126 43496 30132
rect 40960 30048 41012 30054
rect 40960 29990 41012 29996
rect 40972 29714 41000 29990
rect 40960 29708 41012 29714
rect 40960 29650 41012 29656
rect 40224 29504 40276 29510
rect 40224 29446 40276 29452
rect 39396 29300 39448 29306
rect 39396 29242 39448 29248
rect 40132 28960 40184 28966
rect 40132 28902 40184 28908
rect 40144 28626 40172 28902
rect 40132 28620 40184 28626
rect 40132 28562 40184 28568
rect 40236 28422 40264 29446
rect 41144 29232 41196 29238
rect 41144 29174 41196 29180
rect 40868 29164 40920 29170
rect 40868 29106 40920 29112
rect 40880 28626 40908 29106
rect 41156 29102 41184 29174
rect 41144 29096 41196 29102
rect 41144 29038 41196 29044
rect 40868 28620 40920 28626
rect 40868 28562 40920 28568
rect 40224 28416 40276 28422
rect 40224 28358 40276 28364
rect 40880 28082 40908 28562
rect 40868 28076 40920 28082
rect 40868 28018 40920 28024
rect 40408 26920 40460 26926
rect 40408 26862 40460 26868
rect 40420 26586 40448 26862
rect 41156 26586 41184 29038
rect 41420 28416 41472 28422
rect 41248 28364 41420 28370
rect 41248 28358 41472 28364
rect 41248 28342 41460 28358
rect 41248 28014 41276 28342
rect 41236 28008 41288 28014
rect 41236 27950 41288 27956
rect 41248 27402 41276 27950
rect 41236 27396 41288 27402
rect 41236 27338 41288 27344
rect 41248 26926 41276 27338
rect 41236 26920 41288 26926
rect 41236 26862 41288 26868
rect 40408 26580 40460 26586
rect 40408 26522 40460 26528
rect 41144 26580 41196 26586
rect 41144 26522 41196 26528
rect 41248 26382 41276 26862
rect 41236 26376 41288 26382
rect 41236 26318 41288 26324
rect 40868 26240 40920 26246
rect 40868 26182 40920 26188
rect 40880 26042 40908 26182
rect 40868 26036 40920 26042
rect 40868 25978 40920 25984
rect 40880 25362 40908 25978
rect 41236 25832 41288 25838
rect 41236 25774 41288 25780
rect 40868 25356 40920 25362
rect 40868 25298 40920 25304
rect 41248 25158 41276 25774
rect 42444 25498 42472 30126
rect 42616 29572 42668 29578
rect 42616 29514 42668 29520
rect 42628 29306 42656 29514
rect 42616 29300 42668 29306
rect 42616 29242 42668 29248
rect 42984 29300 43036 29306
rect 42984 29242 43036 29248
rect 42708 29164 42760 29170
rect 42708 29106 42760 29112
rect 42720 27674 42748 29106
rect 42800 29028 42852 29034
rect 42800 28970 42852 28976
rect 42812 28694 42840 28970
rect 42800 28688 42852 28694
rect 42800 28630 42852 28636
rect 42812 28218 42840 28630
rect 42892 28416 42944 28422
rect 42892 28358 42944 28364
rect 42800 28212 42852 28218
rect 42800 28154 42852 28160
rect 42904 28150 42932 28358
rect 42892 28144 42944 28150
rect 42892 28086 42944 28092
rect 42800 28076 42852 28082
rect 42800 28018 42852 28024
rect 42708 27668 42760 27674
rect 42628 27628 42708 27656
rect 42432 25492 42484 25498
rect 42432 25434 42484 25440
rect 42524 25424 42576 25430
rect 42524 25366 42576 25372
rect 41420 25288 41472 25294
rect 41420 25230 41472 25236
rect 42156 25288 42208 25294
rect 42156 25230 42208 25236
rect 39764 25152 39816 25158
rect 39764 25094 39816 25100
rect 41236 25152 41288 25158
rect 41236 25094 41288 25100
rect 39776 24818 39804 25094
rect 39764 24812 39816 24818
rect 39764 24754 39816 24760
rect 39672 24404 39724 24410
rect 39672 24346 39724 24352
rect 39488 23792 39540 23798
rect 39488 23734 39540 23740
rect 39316 22460 39436 22488
rect 39210 22400 39266 22409
rect 39210 22335 39266 22344
rect 39224 21010 39252 22335
rect 39408 22114 39436 22460
rect 39316 22086 39436 22114
rect 39212 21004 39264 21010
rect 39212 20946 39264 20952
rect 39224 20058 39252 20946
rect 39316 20369 39344 22086
rect 39500 21622 39528 23734
rect 39684 23662 39712 24346
rect 39672 23656 39724 23662
rect 39672 23598 39724 23604
rect 39580 23044 39632 23050
rect 39580 22986 39632 22992
rect 39592 22642 39620 22986
rect 39580 22636 39632 22642
rect 39580 22578 39632 22584
rect 39684 21622 39712 23598
rect 39776 23186 39804 24754
rect 40040 24132 40092 24138
rect 40040 24074 40092 24080
rect 40052 23866 40080 24074
rect 40408 24064 40460 24070
rect 40406 24032 40408 24041
rect 40460 24032 40462 24041
rect 40406 23967 40462 23976
rect 40040 23860 40092 23866
rect 40040 23802 40092 23808
rect 40316 23724 40368 23730
rect 40316 23666 40368 23672
rect 40328 23322 40356 23666
rect 40316 23316 40368 23322
rect 40316 23258 40368 23264
rect 39948 23248 40000 23254
rect 39948 23190 40000 23196
rect 39764 23180 39816 23186
rect 39764 23122 39816 23128
rect 39960 22778 39988 23190
rect 40224 23044 40276 23050
rect 40224 22986 40276 22992
rect 40236 22778 40264 22986
rect 40500 22976 40552 22982
rect 40500 22918 40552 22924
rect 39948 22772 40000 22778
rect 39948 22714 40000 22720
rect 40224 22772 40276 22778
rect 40224 22714 40276 22720
rect 40512 22438 40540 22918
rect 41248 22778 41276 25094
rect 41236 22772 41288 22778
rect 41432 22760 41460 25230
rect 41696 25220 41748 25226
rect 41696 25162 41748 25168
rect 41708 24886 41736 25162
rect 41696 24880 41748 24886
rect 41696 24822 41748 24828
rect 41708 23526 41736 24822
rect 42168 24614 42196 25230
rect 42156 24608 42208 24614
rect 42156 24550 42208 24556
rect 42064 24336 42116 24342
rect 42064 24278 42116 24284
rect 42076 23798 42104 24278
rect 42064 23792 42116 23798
rect 42064 23734 42116 23740
rect 41696 23520 41748 23526
rect 41696 23462 41748 23468
rect 42076 23066 42104 23734
rect 41892 23038 42104 23066
rect 41512 22772 41564 22778
rect 41432 22732 41512 22760
rect 41236 22714 41288 22720
rect 41512 22714 41564 22720
rect 40224 22432 40276 22438
rect 40222 22400 40224 22409
rect 40500 22432 40552 22438
rect 40276 22400 40278 22409
rect 40500 22374 40552 22380
rect 40222 22335 40278 22344
rect 39856 21888 39908 21894
rect 39856 21830 39908 21836
rect 39488 21616 39540 21622
rect 39488 21558 39540 21564
rect 39672 21616 39724 21622
rect 39672 21558 39724 21564
rect 39500 21078 39528 21558
rect 39488 21072 39540 21078
rect 39488 21014 39540 21020
rect 39684 21010 39712 21558
rect 39764 21480 39816 21486
rect 39764 21422 39816 21428
rect 39776 21146 39804 21422
rect 39868 21146 39896 21830
rect 39764 21140 39816 21146
rect 39764 21082 39816 21088
rect 39856 21140 39908 21146
rect 39856 21082 39908 21088
rect 39672 21004 39724 21010
rect 39672 20946 39724 20952
rect 39396 20936 39448 20942
rect 39396 20878 39448 20884
rect 39408 20602 39436 20878
rect 40132 20868 40184 20874
rect 40132 20810 40184 20816
rect 40144 20602 40172 20810
rect 39396 20596 39448 20602
rect 39396 20538 39448 20544
rect 40132 20596 40184 20602
rect 40132 20538 40184 20544
rect 39764 20460 39816 20466
rect 39764 20402 39816 20408
rect 39856 20460 39908 20466
rect 39856 20402 39908 20408
rect 40040 20460 40092 20466
rect 40040 20402 40092 20408
rect 39302 20360 39358 20369
rect 39302 20295 39358 20304
rect 39488 20256 39540 20262
rect 39488 20198 39540 20204
rect 39212 20052 39264 20058
rect 39212 19994 39264 20000
rect 39132 19366 39344 19394
rect 39028 19304 39080 19310
rect 39028 19246 39080 19252
rect 39120 19236 39172 19242
rect 39120 19178 39172 19184
rect 39132 18850 39160 19178
rect 39040 18822 39160 18850
rect 39040 18766 39068 18822
rect 39028 18760 39080 18766
rect 39028 18702 39080 18708
rect 39212 18692 39264 18698
rect 39212 18634 39264 18640
rect 39028 17672 39080 17678
rect 39028 17614 39080 17620
rect 39040 17542 39068 17614
rect 39028 17536 39080 17542
rect 39028 17478 39080 17484
rect 38936 17128 38988 17134
rect 38936 17070 38988 17076
rect 38948 16590 38976 17070
rect 39040 16590 39068 17478
rect 38936 16584 38988 16590
rect 38936 16526 38988 16532
rect 39028 16584 39080 16590
rect 39028 16526 39080 16532
rect 39224 16522 39252 18634
rect 39316 18154 39344 19366
rect 39396 19304 39448 19310
rect 39396 19246 39448 19252
rect 39408 18630 39436 19246
rect 39396 18624 39448 18630
rect 39396 18566 39448 18572
rect 39408 18426 39436 18566
rect 39396 18420 39448 18426
rect 39396 18362 39448 18368
rect 39304 18148 39356 18154
rect 39304 18090 39356 18096
rect 39408 17814 39436 18362
rect 39396 17808 39448 17814
rect 39396 17750 39448 17756
rect 39500 17105 39528 20198
rect 39580 19916 39632 19922
rect 39580 19858 39632 19864
rect 39592 19378 39620 19858
rect 39580 19372 39632 19378
rect 39776 19360 39804 20402
rect 39868 20262 39896 20402
rect 39856 20256 39908 20262
rect 39856 20198 39908 20204
rect 39948 20256 40000 20262
rect 39948 20198 40000 20204
rect 39960 20058 39988 20198
rect 39948 20052 40000 20058
rect 39948 19994 40000 20000
rect 39856 19372 39908 19378
rect 39776 19332 39856 19360
rect 39580 19314 39632 19320
rect 39856 19314 39908 19320
rect 39856 19168 39908 19174
rect 39856 19110 39908 19116
rect 39868 19009 39896 19110
rect 39854 19000 39910 19009
rect 39854 18935 39910 18944
rect 39580 18760 39632 18766
rect 39580 18702 39632 18708
rect 39486 17096 39542 17105
rect 39486 17031 39542 17040
rect 39488 16584 39540 16590
rect 39488 16526 39540 16532
rect 39212 16516 39264 16522
rect 39212 16458 39264 16464
rect 39304 15496 39356 15502
rect 39304 15438 39356 15444
rect 39120 15088 39172 15094
rect 39120 15030 39172 15036
rect 38844 13932 38896 13938
rect 38844 13874 38896 13880
rect 39132 13326 39160 15030
rect 39316 14822 39344 15438
rect 39394 15192 39450 15201
rect 39394 15127 39450 15136
rect 39408 15094 39436 15127
rect 39396 15088 39448 15094
rect 39396 15030 39448 15036
rect 39500 15026 39528 16526
rect 39488 15020 39540 15026
rect 39488 14962 39540 14968
rect 39304 14816 39356 14822
rect 39304 14758 39356 14764
rect 39316 14006 39344 14758
rect 39500 14414 39528 14962
rect 39488 14408 39540 14414
rect 39488 14350 39540 14356
rect 39304 14000 39356 14006
rect 39304 13942 39356 13948
rect 39396 13728 39448 13734
rect 39396 13670 39448 13676
rect 39408 13530 39436 13670
rect 39396 13524 39448 13530
rect 39396 13466 39448 13472
rect 39120 13320 39172 13326
rect 39120 13262 39172 13268
rect 39132 12170 39160 13262
rect 39120 12164 39172 12170
rect 39120 12106 39172 12112
rect 39500 11762 39528 14350
rect 39592 14006 39620 18702
rect 39672 17604 39724 17610
rect 39672 17546 39724 17552
rect 39684 15910 39712 17546
rect 39960 16998 39988 19994
rect 40052 19514 40080 20402
rect 40040 19508 40092 19514
rect 40040 19450 40092 19456
rect 40314 19408 40370 19417
rect 40224 19372 40276 19378
rect 40314 19343 40316 19352
rect 40224 19314 40276 19320
rect 40368 19343 40370 19352
rect 40316 19314 40368 19320
rect 40040 19304 40092 19310
rect 40040 19246 40092 19252
rect 40236 19258 40264 19314
rect 40052 17785 40080 19246
rect 40236 19242 40356 19258
rect 40236 19236 40368 19242
rect 40236 19230 40316 19236
rect 40316 19178 40368 19184
rect 40132 19168 40184 19174
rect 40132 19110 40184 19116
rect 40144 18970 40172 19110
rect 40132 18964 40184 18970
rect 40132 18906 40184 18912
rect 40224 18216 40276 18222
rect 40224 18158 40276 18164
rect 40038 17776 40094 17785
rect 40038 17711 40094 17720
rect 40052 17678 40080 17711
rect 40236 17678 40264 18158
rect 40328 17678 40356 19178
rect 40406 19136 40462 19145
rect 40406 19071 40462 19080
rect 40040 17672 40092 17678
rect 40040 17614 40092 17620
rect 40224 17672 40276 17678
rect 40224 17614 40276 17620
rect 40316 17672 40368 17678
rect 40316 17614 40368 17620
rect 40236 17134 40264 17614
rect 40224 17128 40276 17134
rect 40224 17070 40276 17076
rect 39948 16992 40000 16998
rect 39948 16934 40000 16940
rect 39672 15904 39724 15910
rect 39672 15846 39724 15852
rect 40040 15428 40092 15434
rect 40040 15370 40092 15376
rect 40132 15428 40184 15434
rect 40132 15370 40184 15376
rect 39672 15020 39724 15026
rect 39672 14962 39724 14968
rect 39764 15020 39816 15026
rect 39764 14962 39816 14968
rect 39684 14550 39712 14962
rect 39672 14544 39724 14550
rect 39672 14486 39724 14492
rect 39776 14482 39804 14962
rect 39764 14476 39816 14482
rect 39764 14418 39816 14424
rect 39856 14476 39908 14482
rect 39856 14418 39908 14424
rect 39868 14074 39896 14418
rect 39856 14068 39908 14074
rect 39856 14010 39908 14016
rect 39580 14000 39632 14006
rect 39632 13960 39712 13988
rect 39580 13942 39632 13948
rect 39684 12434 39712 13960
rect 40052 13546 40080 15370
rect 40144 15162 40172 15370
rect 40132 15156 40184 15162
rect 40132 15098 40184 15104
rect 40420 13818 40448 19071
rect 40512 18970 40540 22374
rect 41892 22273 41920 23038
rect 42064 22772 42116 22778
rect 42064 22714 42116 22720
rect 41878 22264 41934 22273
rect 40592 22228 40644 22234
rect 41878 22199 41934 22208
rect 40592 22170 40644 22176
rect 40604 21418 40632 22170
rect 41604 21956 41656 21962
rect 41604 21898 41656 21904
rect 41788 21956 41840 21962
rect 41788 21898 41840 21904
rect 40592 21412 40644 21418
rect 40592 21354 40644 21360
rect 40604 19417 40632 21354
rect 41144 20868 41196 20874
rect 41144 20810 41196 20816
rect 41156 20602 41184 20810
rect 41512 20800 41564 20806
rect 41512 20742 41564 20748
rect 41144 20596 41196 20602
rect 41144 20538 41196 20544
rect 41524 20398 41552 20742
rect 41616 20466 41644 21898
rect 41800 21146 41828 21898
rect 41788 21140 41840 21146
rect 41788 21082 41840 21088
rect 41604 20460 41656 20466
rect 41604 20402 41656 20408
rect 41052 20392 41104 20398
rect 41052 20334 41104 20340
rect 41512 20392 41564 20398
rect 41512 20334 41564 20340
rect 40684 19916 40736 19922
rect 40684 19858 40736 19864
rect 40590 19408 40646 19417
rect 40696 19378 40724 19858
rect 40868 19780 40920 19786
rect 40868 19722 40920 19728
rect 40774 19408 40830 19417
rect 40590 19343 40646 19352
rect 40684 19372 40736 19378
rect 40604 19258 40632 19343
rect 40774 19343 40776 19352
rect 40684 19314 40736 19320
rect 40828 19343 40830 19352
rect 40880 19360 40908 19722
rect 41064 19417 41092 20334
rect 41800 19553 41828 21082
rect 41786 19544 41842 19553
rect 41786 19479 41842 19488
rect 41050 19408 41106 19417
rect 40960 19372 41012 19378
rect 40880 19332 40960 19360
rect 40776 19314 40828 19320
rect 41050 19343 41106 19352
rect 40960 19314 41012 19320
rect 40604 19230 40908 19258
rect 40500 18964 40552 18970
rect 40500 18906 40552 18912
rect 40684 18896 40736 18902
rect 40684 18838 40736 18844
rect 40696 18290 40724 18838
rect 40880 18698 40908 19230
rect 40868 18692 40920 18698
rect 40868 18634 40920 18640
rect 40684 18284 40736 18290
rect 40684 18226 40736 18232
rect 40880 17882 40908 18634
rect 40868 17876 40920 17882
rect 40868 17818 40920 17824
rect 40868 17740 40920 17746
rect 40868 17682 40920 17688
rect 40592 17604 40644 17610
rect 40592 17546 40644 17552
rect 40604 15706 40632 17546
rect 40880 16658 40908 17682
rect 40972 17678 41000 19314
rect 41050 19272 41106 19281
rect 41050 19207 41106 19216
rect 41064 18970 41092 19207
rect 41512 19168 41564 19174
rect 41512 19110 41564 19116
rect 41052 18964 41104 18970
rect 41052 18906 41104 18912
rect 41064 18766 41092 18906
rect 41052 18760 41104 18766
rect 41052 18702 41104 18708
rect 41524 18358 41552 19110
rect 41696 18624 41748 18630
rect 41696 18566 41748 18572
rect 41512 18352 41564 18358
rect 41512 18294 41564 18300
rect 41328 17876 41380 17882
rect 41328 17818 41380 17824
rect 41340 17746 41368 17818
rect 41328 17740 41380 17746
rect 41328 17682 41380 17688
rect 40960 17672 41012 17678
rect 40960 17614 41012 17620
rect 41420 17604 41472 17610
rect 41420 17546 41472 17552
rect 41328 17536 41380 17542
rect 41328 17478 41380 17484
rect 41236 17264 41288 17270
rect 41236 17206 41288 17212
rect 41052 17196 41104 17202
rect 41052 17138 41104 17144
rect 41064 16794 41092 17138
rect 41052 16788 41104 16794
rect 41052 16730 41104 16736
rect 40868 16652 40920 16658
rect 40868 16594 40920 16600
rect 40592 15700 40644 15706
rect 40592 15642 40644 15648
rect 40880 15570 40908 16594
rect 41248 15688 41276 17206
rect 41340 17202 41368 17478
rect 41432 17202 41460 17546
rect 41328 17196 41380 17202
rect 41328 17138 41380 17144
rect 41420 17196 41472 17202
rect 41420 17138 41472 17144
rect 41418 17096 41474 17105
rect 41418 17031 41420 17040
rect 41472 17031 41474 17040
rect 41420 17002 41472 17008
rect 41328 16992 41380 16998
rect 41328 16934 41380 16940
rect 41340 16658 41368 16934
rect 41328 16652 41380 16658
rect 41328 16594 41380 16600
rect 41524 16250 41552 18294
rect 41708 17202 41736 18566
rect 41696 17196 41748 17202
rect 41696 17138 41748 17144
rect 41708 17066 41736 17138
rect 41696 17060 41748 17066
rect 41696 17002 41748 17008
rect 41512 16244 41564 16250
rect 41512 16186 41564 16192
rect 41420 15700 41472 15706
rect 41248 15660 41420 15688
rect 41420 15642 41472 15648
rect 40868 15564 40920 15570
rect 40868 15506 40920 15512
rect 41432 15434 41460 15642
rect 41420 15428 41472 15434
rect 41420 15370 41472 15376
rect 41432 15201 41460 15370
rect 41604 15360 41656 15366
rect 41604 15302 41656 15308
rect 41418 15192 41474 15201
rect 41418 15127 41474 15136
rect 41050 15056 41106 15065
rect 41616 15026 41644 15302
rect 41050 14991 41052 15000
rect 41104 14991 41106 15000
rect 41604 15020 41656 15026
rect 41052 14962 41104 14968
rect 41604 14962 41656 14968
rect 41788 15020 41840 15026
rect 41788 14962 41840 14968
rect 41420 14884 41472 14890
rect 41420 14826 41472 14832
rect 40590 13968 40646 13977
rect 40590 13903 40592 13912
rect 40644 13903 40646 13912
rect 40592 13874 40644 13880
rect 40420 13790 40540 13818
rect 40408 13728 40460 13734
rect 40408 13670 40460 13676
rect 39960 13518 40080 13546
rect 40420 13530 40448 13670
rect 40512 13530 40540 13790
rect 40408 13524 40460 13530
rect 39764 13456 39816 13462
rect 39764 13398 39816 13404
rect 39592 12406 39712 12434
rect 39488 11756 39540 11762
rect 39488 11698 39540 11704
rect 39028 11008 39080 11014
rect 39028 10950 39080 10956
rect 38844 10804 38896 10810
rect 38844 10746 38896 10752
rect 38752 10668 38804 10674
rect 38752 10610 38804 10616
rect 38856 10062 38884 10746
rect 39040 10742 39068 10950
rect 39592 10810 39620 12406
rect 39672 11620 39724 11626
rect 39672 11562 39724 11568
rect 39684 11286 39712 11562
rect 39672 11280 39724 11286
rect 39672 11222 39724 11228
rect 39670 10976 39726 10985
rect 39670 10911 39726 10920
rect 39580 10804 39632 10810
rect 39580 10746 39632 10752
rect 39028 10736 39080 10742
rect 39028 10678 39080 10684
rect 39684 10266 39712 10911
rect 39672 10260 39724 10266
rect 39672 10202 39724 10208
rect 39684 10062 39712 10202
rect 39776 10198 39804 13398
rect 39856 13320 39908 13326
rect 39856 13262 39908 13268
rect 39868 12782 39896 13262
rect 39960 13138 39988 13518
rect 40408 13466 40460 13472
rect 40500 13524 40552 13530
rect 40500 13466 40552 13472
rect 40040 13456 40092 13462
rect 40040 13398 40092 13404
rect 40052 13326 40080 13398
rect 40512 13326 40540 13466
rect 40776 13456 40828 13462
rect 40774 13424 40776 13433
rect 40828 13424 40830 13433
rect 40774 13359 40830 13368
rect 40040 13320 40092 13326
rect 40040 13262 40092 13268
rect 40500 13320 40552 13326
rect 40500 13262 40552 13268
rect 40776 13320 40828 13326
rect 40776 13262 40828 13268
rect 40132 13252 40184 13258
rect 40132 13194 40184 13200
rect 39960 13110 40080 13138
rect 39856 12776 39908 12782
rect 39856 12718 39908 12724
rect 39764 10192 39816 10198
rect 39764 10134 39816 10140
rect 39856 10124 39908 10130
rect 39856 10066 39908 10072
rect 38844 10056 38896 10062
rect 38844 9998 38896 10004
rect 39212 10056 39264 10062
rect 39672 10056 39724 10062
rect 39264 10004 39344 10010
rect 39212 9998 39344 10004
rect 39672 9998 39724 10004
rect 39224 9982 39344 9998
rect 38672 9654 38976 9674
rect 38672 9648 38988 9654
rect 38672 9646 38936 9648
rect 38936 9590 38988 9596
rect 38384 9376 38436 9382
rect 38384 9318 38436 9324
rect 38396 9178 38424 9318
rect 38384 9172 38436 9178
rect 38384 9114 38436 9120
rect 38568 9104 38620 9110
rect 38568 9046 38620 9052
rect 38292 8968 38344 8974
rect 38292 8910 38344 8916
rect 38384 8968 38436 8974
rect 38384 8910 38436 8916
rect 38476 8968 38528 8974
rect 38476 8910 38528 8916
rect 38396 8838 38424 8910
rect 38384 8832 38436 8838
rect 38212 8780 38384 8786
rect 38212 8774 38436 8780
rect 38212 8758 38424 8774
rect 38488 8634 38516 8910
rect 38476 8628 38528 8634
rect 38476 8570 38528 8576
rect 38108 8560 38160 8566
rect 38108 8502 38160 8508
rect 38016 8356 38068 8362
rect 38016 8298 38068 8304
rect 37372 6870 37424 6876
rect 37830 6896 37886 6905
rect 37188 6860 37240 6866
rect 37830 6831 37886 6840
rect 37188 6802 37240 6808
rect 36636 6316 36688 6322
rect 36636 6258 36688 6264
rect 36832 6310 37044 6338
rect 36648 5710 36676 6258
rect 36832 5914 36860 6310
rect 36912 6248 36964 6254
rect 36912 6190 36964 6196
rect 36820 5908 36872 5914
rect 36820 5850 36872 5856
rect 36832 5710 36860 5850
rect 36924 5710 36952 6190
rect 36636 5704 36688 5710
rect 36636 5646 36688 5652
rect 36820 5704 36872 5710
rect 36820 5646 36872 5652
rect 36912 5704 36964 5710
rect 36912 5646 36964 5652
rect 36924 5370 36952 5646
rect 37200 5574 37228 6802
rect 37464 6792 37516 6798
rect 37464 6734 37516 6740
rect 37476 5846 37504 6734
rect 37556 6180 37608 6186
rect 37556 6122 37608 6128
rect 37464 5840 37516 5846
rect 37464 5782 37516 5788
rect 37476 5710 37504 5782
rect 37464 5704 37516 5710
rect 37464 5646 37516 5652
rect 37372 5636 37424 5642
rect 37372 5578 37424 5584
rect 37188 5568 37240 5574
rect 37188 5510 37240 5516
rect 36544 5364 36596 5370
rect 36544 5306 36596 5312
rect 36912 5364 36964 5370
rect 36912 5306 36964 5312
rect 36556 5234 36584 5306
rect 36412 5188 36492 5216
rect 36544 5228 36596 5234
rect 36360 5170 36412 5176
rect 36544 5170 36596 5176
rect 36372 4622 36400 5170
rect 37096 5160 37148 5166
rect 37200 5114 37228 5510
rect 37384 5234 37412 5578
rect 37464 5568 37516 5574
rect 37464 5510 37516 5516
rect 37476 5234 37504 5510
rect 37372 5228 37424 5234
rect 37372 5170 37424 5176
rect 37464 5228 37516 5234
rect 37464 5170 37516 5176
rect 37148 5108 37228 5114
rect 37096 5102 37228 5108
rect 37108 5086 37228 5102
rect 36452 5024 36504 5030
rect 36452 4966 36504 4972
rect 36360 4616 36412 4622
rect 36360 4558 36412 4564
rect 35992 4548 36044 4554
rect 35992 4490 36044 4496
rect 36084 4548 36136 4554
rect 36084 4490 36136 4496
rect 35256 4480 35308 4486
rect 35256 4422 35308 4428
rect 35268 4078 35296 4422
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 36004 4282 36032 4490
rect 35992 4276 36044 4282
rect 35992 4218 36044 4224
rect 36096 4146 36124 4490
rect 36360 4480 36412 4486
rect 36360 4422 36412 4428
rect 36268 4208 36320 4214
rect 36268 4150 36320 4156
rect 36084 4140 36136 4146
rect 36004 4100 36084 4128
rect 34060 4072 34112 4078
rect 34060 4014 34112 4020
rect 35256 4072 35308 4078
rect 35256 4014 35308 4020
rect 31852 3936 31904 3942
rect 31852 3878 31904 3884
rect 31944 3936 31996 3942
rect 31944 3878 31996 3884
rect 31760 3664 31812 3670
rect 31760 3606 31812 3612
rect 30196 3596 30248 3602
rect 30196 3538 30248 3544
rect 31864 3534 31892 3878
rect 31956 3738 31984 3878
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 31944 3732 31996 3738
rect 31944 3674 31996 3680
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 31864 3194 31892 3470
rect 31944 3392 31996 3398
rect 31944 3334 31996 3340
rect 31852 3188 31904 3194
rect 31852 3130 31904 3136
rect 31956 3058 31984 3334
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 36004 3194 36032 4100
rect 36084 4082 36136 4088
rect 36176 3936 36228 3942
rect 36176 3878 36228 3884
rect 35992 3188 36044 3194
rect 35992 3130 36044 3136
rect 31944 3052 31996 3058
rect 31944 2994 31996 3000
rect 36188 2990 36216 3878
rect 36280 3126 36308 4150
rect 36372 4146 36400 4422
rect 36464 4146 36492 4966
rect 36360 4140 36412 4146
rect 36360 4082 36412 4088
rect 36452 4140 36504 4146
rect 36452 4082 36504 4088
rect 37108 4078 37136 5086
rect 37568 5030 37596 6122
rect 37188 5024 37240 5030
rect 37188 4966 37240 4972
rect 37556 5024 37608 5030
rect 37556 4966 37608 4972
rect 37200 4690 37228 4966
rect 37188 4684 37240 4690
rect 37188 4626 37240 4632
rect 37096 4072 37148 4078
rect 37096 4014 37148 4020
rect 36268 3120 36320 3126
rect 36268 3062 36320 3068
rect 37108 2990 37136 4014
rect 37568 4010 37596 4966
rect 37648 4548 37700 4554
rect 37648 4490 37700 4496
rect 37660 4214 37688 4490
rect 37844 4282 37872 6831
rect 37832 4276 37884 4282
rect 37832 4218 37884 4224
rect 37648 4208 37700 4214
rect 37648 4150 37700 4156
rect 37556 4004 37608 4010
rect 37556 3946 37608 3952
rect 36176 2984 36228 2990
rect 36176 2926 36228 2932
rect 37096 2984 37148 2990
rect 37096 2926 37148 2932
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 32968 2446 32996 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 38028 2446 38056 8298
rect 38120 6866 38148 8502
rect 38580 8480 38608 9046
rect 38844 8832 38896 8838
rect 38844 8774 38896 8780
rect 38488 8452 38608 8480
rect 38292 8288 38344 8294
rect 38292 8230 38344 8236
rect 38304 6934 38332 8230
rect 38488 7954 38516 8452
rect 38476 7948 38528 7954
rect 38476 7890 38528 7896
rect 38292 6928 38344 6934
rect 38292 6870 38344 6876
rect 38108 6860 38160 6866
rect 38160 6820 38240 6848
rect 38108 6802 38160 6808
rect 38108 6656 38160 6662
rect 38108 6598 38160 6604
rect 38120 6322 38148 6598
rect 38108 6316 38160 6322
rect 38108 6258 38160 6264
rect 38212 6254 38240 6820
rect 38304 6798 38332 6870
rect 38292 6792 38344 6798
rect 38292 6734 38344 6740
rect 38384 6724 38436 6730
rect 38384 6666 38436 6672
rect 38200 6248 38252 6254
rect 38200 6190 38252 6196
rect 38108 6112 38160 6118
rect 38108 6054 38160 6060
rect 38120 5778 38148 6054
rect 38108 5772 38160 5778
rect 38108 5714 38160 5720
rect 38396 5302 38424 6666
rect 38488 6186 38516 7890
rect 38856 7886 38884 8774
rect 38844 7880 38896 7886
rect 38844 7822 38896 7828
rect 38660 7744 38712 7750
rect 38660 7686 38712 7692
rect 38752 7744 38804 7750
rect 38752 7686 38804 7692
rect 38672 7546 38700 7686
rect 38660 7540 38712 7546
rect 38660 7482 38712 7488
rect 38764 7342 38792 7686
rect 38752 7336 38804 7342
rect 38752 7278 38804 7284
rect 38752 7200 38804 7206
rect 38752 7142 38804 7148
rect 38764 6798 38792 7142
rect 38752 6792 38804 6798
rect 38752 6734 38804 6740
rect 38764 6390 38792 6734
rect 38752 6384 38804 6390
rect 38752 6326 38804 6332
rect 38476 6180 38528 6186
rect 38476 6122 38528 6128
rect 38384 5296 38436 5302
rect 38384 5238 38436 5244
rect 38396 4758 38424 5238
rect 38384 4752 38436 4758
rect 38384 4694 38436 4700
rect 38200 4208 38252 4214
rect 38200 4150 38252 4156
rect 38212 3670 38240 4150
rect 38856 3942 38884 7822
rect 38844 3936 38896 3942
rect 38844 3878 38896 3884
rect 38200 3664 38252 3670
rect 38200 3606 38252 3612
rect 38212 2446 38240 3606
rect 38948 3466 38976 9590
rect 39316 9382 39344 9982
rect 39304 9376 39356 9382
rect 39304 9318 39356 9324
rect 39488 9376 39540 9382
rect 39488 9318 39540 9324
rect 39212 8356 39264 8362
rect 39212 8298 39264 8304
rect 39224 7886 39252 8298
rect 39316 7886 39344 9318
rect 39500 8974 39528 9318
rect 39488 8968 39540 8974
rect 39488 8910 39540 8916
rect 39868 7954 39896 10066
rect 40052 9654 40080 13110
rect 40144 12918 40172 13194
rect 40408 13184 40460 13190
rect 40408 13126 40460 13132
rect 40132 12912 40184 12918
rect 40132 12854 40184 12860
rect 40144 11626 40172 12854
rect 40224 12232 40276 12238
rect 40224 12174 40276 12180
rect 40132 11620 40184 11626
rect 40132 11562 40184 11568
rect 40236 10606 40264 12174
rect 40224 10600 40276 10606
rect 40224 10542 40276 10548
rect 40236 10130 40264 10542
rect 40224 10124 40276 10130
rect 40224 10066 40276 10072
rect 40224 9988 40276 9994
rect 40224 9930 40276 9936
rect 40236 9722 40264 9930
rect 40224 9716 40276 9722
rect 40224 9658 40276 9664
rect 40040 9648 40092 9654
rect 40040 9590 40092 9596
rect 40316 9376 40368 9382
rect 40316 9318 40368 9324
rect 40328 9110 40356 9318
rect 40316 9104 40368 9110
rect 40316 9046 40368 9052
rect 40328 8430 40356 9046
rect 40316 8424 40368 8430
rect 40316 8366 40368 8372
rect 40132 8288 40184 8294
rect 40132 8230 40184 8236
rect 40144 7954 40172 8230
rect 39856 7948 39908 7954
rect 39856 7890 39908 7896
rect 40132 7948 40184 7954
rect 40132 7890 40184 7896
rect 39212 7880 39264 7886
rect 39212 7822 39264 7828
rect 39304 7880 39356 7886
rect 39304 7822 39356 7828
rect 39316 6866 39344 7822
rect 39868 7410 39896 7890
rect 39856 7404 39908 7410
rect 39856 7346 39908 7352
rect 39304 6860 39356 6866
rect 39304 6802 39356 6808
rect 39764 6248 39816 6254
rect 39764 6190 39816 6196
rect 39776 5914 39804 6190
rect 39764 5908 39816 5914
rect 39764 5850 39816 5856
rect 39856 4616 39908 4622
rect 39856 4558 39908 4564
rect 39580 4208 39632 4214
rect 39580 4150 39632 4156
rect 39592 3942 39620 4150
rect 39580 3936 39632 3942
rect 39580 3878 39632 3884
rect 38936 3460 38988 3466
rect 38936 3402 38988 3408
rect 39868 3126 39896 4558
rect 40132 4548 40184 4554
rect 40132 4490 40184 4496
rect 40144 4282 40172 4490
rect 40132 4276 40184 4282
rect 40132 4218 40184 4224
rect 39856 3120 39908 3126
rect 39856 3062 39908 3068
rect 38660 3052 38712 3058
rect 38660 2994 38712 3000
rect 40040 3052 40092 3058
rect 40040 2994 40092 3000
rect 38672 2650 38700 2994
rect 39488 2916 39540 2922
rect 39488 2858 39540 2864
rect 39396 2848 39448 2854
rect 39316 2808 39396 2836
rect 38660 2644 38712 2650
rect 38660 2586 38712 2592
rect 32956 2440 33008 2446
rect 32956 2382 33008 2388
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 38200 2440 38252 2446
rect 38200 2382 38252 2388
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 32876 800 32904 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 39316 800 39344 2808
rect 39396 2790 39448 2796
rect 39500 2514 39528 2858
rect 40052 2650 40080 2994
rect 40420 2774 40448 13126
rect 40592 12844 40644 12850
rect 40592 12786 40644 12792
rect 40604 11898 40632 12786
rect 40684 12640 40736 12646
rect 40684 12582 40736 12588
rect 40696 12306 40724 12582
rect 40684 12300 40736 12306
rect 40684 12242 40736 12248
rect 40592 11892 40644 11898
rect 40592 11834 40644 11840
rect 40684 9580 40736 9586
rect 40684 9522 40736 9528
rect 40696 8838 40724 9522
rect 40684 8832 40736 8838
rect 40684 8774 40736 8780
rect 40788 8401 40816 13262
rect 41432 12850 41460 14826
rect 41800 14414 41828 14962
rect 41512 14408 41564 14414
rect 41512 14350 41564 14356
rect 41788 14408 41840 14414
rect 41788 14350 41840 14356
rect 41524 13394 41552 14350
rect 41696 14340 41748 14346
rect 41696 14282 41748 14288
rect 41708 13682 41736 14282
rect 41892 14278 41920 22199
rect 41972 21956 42024 21962
rect 41972 21898 42024 21904
rect 41984 20942 42012 21898
rect 41972 20936 42024 20942
rect 41972 20878 42024 20884
rect 42076 15178 42104 22714
rect 42168 21962 42196 24550
rect 42248 24200 42300 24206
rect 42248 24142 42300 24148
rect 42260 23594 42288 24142
rect 42340 24064 42392 24070
rect 42340 24006 42392 24012
rect 42248 23588 42300 23594
rect 42248 23530 42300 23536
rect 42260 23118 42288 23530
rect 42352 23322 42380 24006
rect 42340 23316 42392 23322
rect 42340 23258 42392 23264
rect 42248 23112 42300 23118
rect 42248 23054 42300 23060
rect 42156 21956 42208 21962
rect 42156 21898 42208 21904
rect 42156 21616 42208 21622
rect 42156 21558 42208 21564
rect 42168 20874 42196 21558
rect 42156 20868 42208 20874
rect 42156 20810 42208 20816
rect 42260 18630 42288 23054
rect 42352 22642 42380 23258
rect 42536 23186 42564 25366
rect 42628 25294 42656 27628
rect 42708 27610 42760 27616
rect 42812 26994 42840 28018
rect 42996 28014 43024 29242
rect 43456 29238 43484 30126
rect 43444 29232 43496 29238
rect 43444 29174 43496 29180
rect 43076 29096 43128 29102
rect 43076 29038 43128 29044
rect 42984 28008 43036 28014
rect 42904 27968 42984 27996
rect 42904 27606 42932 27968
rect 42984 27950 43036 27956
rect 42984 27872 43036 27878
rect 42984 27814 43036 27820
rect 42892 27600 42944 27606
rect 42892 27542 42944 27548
rect 42996 27470 43024 27814
rect 42984 27464 43036 27470
rect 42984 27406 43036 27412
rect 42800 26988 42852 26994
rect 42800 26930 42852 26936
rect 42708 26784 42760 26790
rect 42708 26726 42760 26732
rect 42616 25288 42668 25294
rect 42616 25230 42668 25236
rect 42628 24993 42656 25230
rect 42614 24984 42670 24993
rect 42614 24919 42670 24928
rect 42616 24812 42668 24818
rect 42616 24754 42668 24760
rect 42720 24800 42748 26726
rect 42800 26580 42852 26586
rect 42800 26522 42852 26528
rect 42812 25906 42840 26522
rect 43088 26042 43116 29038
rect 43640 28994 43668 30194
rect 43812 30048 43864 30054
rect 43812 29990 43864 29996
rect 43824 29646 43852 29990
rect 43812 29640 43864 29646
rect 43812 29582 43864 29588
rect 43456 28966 43668 28994
rect 43456 28762 43484 28966
rect 43444 28756 43496 28762
rect 43444 28698 43496 28704
rect 43168 28416 43220 28422
rect 43168 28358 43220 28364
rect 43076 26036 43128 26042
rect 43076 25978 43128 25984
rect 42800 25900 42852 25906
rect 42800 25842 42852 25848
rect 42812 25430 42840 25842
rect 42800 25424 42852 25430
rect 42852 25372 42932 25378
rect 42800 25366 42932 25372
rect 42812 25350 42932 25366
rect 42904 24818 42932 25350
rect 43088 24954 43116 25978
rect 43180 25974 43208 28358
rect 43352 27464 43404 27470
rect 43352 27406 43404 27412
rect 43260 27328 43312 27334
rect 43260 27270 43312 27276
rect 43272 26926 43300 27270
rect 43364 26926 43392 27406
rect 43260 26920 43312 26926
rect 43260 26862 43312 26868
rect 43352 26920 43404 26926
rect 43352 26862 43404 26868
rect 43456 26874 43484 28698
rect 43536 28552 43588 28558
rect 43536 28494 43588 28500
rect 43548 28082 43576 28494
rect 43536 28076 43588 28082
rect 43536 28018 43588 28024
rect 43720 28076 43772 28082
rect 43720 28018 43772 28024
rect 43548 27674 43576 28018
rect 43628 27872 43680 27878
rect 43628 27814 43680 27820
rect 43536 27668 43588 27674
rect 43536 27610 43588 27616
rect 43640 27470 43668 27814
rect 43732 27470 43760 28018
rect 43628 27464 43680 27470
rect 43628 27406 43680 27412
rect 43720 27464 43772 27470
rect 43720 27406 43772 27412
rect 43640 27010 43668 27406
rect 43732 27130 43760 27406
rect 43720 27124 43772 27130
rect 43720 27066 43772 27072
rect 43548 26994 43668 27010
rect 43536 26988 43668 26994
rect 43588 26982 43668 26988
rect 43536 26930 43588 26936
rect 43456 26846 43576 26874
rect 43640 26858 43668 26982
rect 43168 25968 43220 25974
rect 43168 25910 43220 25916
rect 43180 25362 43208 25910
rect 43168 25356 43220 25362
rect 43168 25298 43220 25304
rect 43076 24948 43128 24954
rect 43076 24890 43128 24896
rect 43180 24818 43208 25298
rect 43352 25220 43404 25226
rect 43352 25162 43404 25168
rect 42800 24812 42852 24818
rect 42720 24772 42800 24800
rect 42628 24342 42656 24754
rect 42616 24336 42668 24342
rect 42616 24278 42668 24284
rect 42720 24206 42748 24772
rect 42800 24754 42852 24760
rect 42892 24812 42944 24818
rect 42892 24754 42944 24760
rect 43168 24812 43220 24818
rect 43168 24754 43220 24760
rect 43364 24682 43392 25162
rect 43352 24676 43404 24682
rect 43352 24618 43404 24624
rect 43076 24404 43128 24410
rect 43076 24346 43128 24352
rect 42708 24200 42760 24206
rect 42708 24142 42760 24148
rect 43088 24120 43116 24346
rect 43260 24268 43312 24274
rect 43260 24210 43312 24216
rect 43272 24120 43300 24210
rect 43088 24092 43300 24120
rect 42892 24064 42944 24070
rect 42892 24006 42944 24012
rect 42708 23792 42760 23798
rect 42708 23734 42760 23740
rect 42720 23254 42748 23734
rect 42708 23248 42760 23254
rect 42708 23190 42760 23196
rect 42524 23180 42576 23186
rect 42524 23122 42576 23128
rect 42524 23044 42576 23050
rect 42524 22986 42576 22992
rect 42340 22636 42392 22642
rect 42340 22578 42392 22584
rect 42536 22098 42564 22986
rect 42616 22976 42668 22982
rect 42616 22918 42668 22924
rect 42628 22642 42656 22918
rect 42720 22642 42748 23190
rect 42904 23050 42932 24006
rect 43088 23186 43116 24092
rect 43076 23180 43128 23186
rect 43076 23122 43128 23128
rect 42984 23112 43036 23118
rect 42984 23054 43036 23060
rect 42892 23044 42944 23050
rect 42892 22986 42944 22992
rect 42904 22953 42932 22986
rect 42890 22944 42946 22953
rect 42890 22879 42946 22888
rect 42616 22636 42668 22642
rect 42616 22578 42668 22584
rect 42708 22636 42760 22642
rect 42708 22578 42760 22584
rect 42524 22092 42576 22098
rect 42524 22034 42576 22040
rect 42616 22024 42668 22030
rect 42616 21966 42668 21972
rect 42628 21418 42656 21966
rect 42800 21956 42852 21962
rect 42800 21898 42852 21904
rect 42616 21412 42668 21418
rect 42616 21354 42668 21360
rect 42812 20874 42840 21898
rect 42524 20868 42576 20874
rect 42524 20810 42576 20816
rect 42800 20868 42852 20874
rect 42800 20810 42852 20816
rect 42536 20330 42564 20810
rect 42708 20800 42760 20806
rect 42708 20742 42760 20748
rect 42524 20324 42576 20330
rect 42524 20266 42576 20272
rect 42720 19854 42748 20742
rect 42708 19848 42760 19854
rect 42708 19790 42760 19796
rect 42616 19508 42668 19514
rect 42616 19450 42668 19456
rect 42340 19440 42392 19446
rect 42340 19382 42392 19388
rect 42248 18624 42300 18630
rect 42248 18566 42300 18572
rect 42248 18216 42300 18222
rect 42248 18158 42300 18164
rect 42260 17882 42288 18158
rect 42248 17876 42300 17882
rect 42248 17818 42300 17824
rect 42352 17082 42380 19382
rect 42432 17740 42484 17746
rect 42432 17682 42484 17688
rect 42524 17740 42576 17746
rect 42524 17682 42576 17688
rect 42444 17134 42472 17682
rect 42260 17054 42380 17082
rect 42432 17128 42484 17134
rect 42432 17070 42484 17076
rect 42156 15428 42208 15434
rect 42156 15370 42208 15376
rect 41984 15150 42104 15178
rect 42168 15162 42196 15370
rect 42156 15156 42208 15162
rect 41880 14272 41932 14278
rect 41880 14214 41932 14220
rect 41616 13654 41736 13682
rect 41512 13388 41564 13394
rect 41512 13330 41564 13336
rect 41420 12844 41472 12850
rect 41420 12786 41472 12792
rect 41616 12434 41644 13654
rect 41696 13524 41748 13530
rect 41696 13466 41748 13472
rect 41708 13326 41736 13466
rect 41696 13320 41748 13326
rect 41696 13262 41748 13268
rect 41616 12406 41736 12434
rect 41708 11558 41736 12406
rect 41696 11552 41748 11558
rect 41696 11494 41748 11500
rect 41708 10742 41736 11494
rect 41788 11348 41840 11354
rect 41788 11290 41840 11296
rect 41800 11218 41828 11290
rect 41788 11212 41840 11218
rect 41788 11154 41840 11160
rect 41696 10736 41748 10742
rect 41696 10678 41748 10684
rect 41800 10674 41828 11154
rect 41420 10668 41472 10674
rect 41420 10610 41472 10616
rect 41788 10668 41840 10674
rect 41788 10610 41840 10616
rect 41236 9920 41288 9926
rect 41236 9862 41288 9868
rect 40868 8832 40920 8838
rect 40868 8774 40920 8780
rect 40880 8430 40908 8774
rect 40868 8424 40920 8430
rect 40774 8392 40830 8401
rect 40868 8366 40920 8372
rect 40774 8327 40830 8336
rect 40788 7546 40816 8327
rect 41248 7886 41276 9862
rect 41432 8566 41460 10610
rect 41696 10600 41748 10606
rect 41696 10542 41748 10548
rect 41708 9926 41736 10542
rect 41696 9920 41748 9926
rect 41696 9862 41748 9868
rect 41708 9518 41736 9862
rect 41696 9512 41748 9518
rect 41696 9454 41748 9460
rect 41696 8900 41748 8906
rect 41696 8842 41748 8848
rect 41708 8566 41736 8842
rect 41788 8832 41840 8838
rect 41788 8774 41840 8780
rect 41420 8560 41472 8566
rect 41420 8502 41472 8508
rect 41696 8560 41748 8566
rect 41696 8502 41748 8508
rect 41236 7880 41288 7886
rect 41236 7822 41288 7828
rect 40776 7540 40828 7546
rect 40776 7482 40828 7488
rect 40776 7404 40828 7410
rect 40776 7346 40828 7352
rect 40498 7032 40554 7041
rect 40498 6967 40554 6976
rect 40512 6798 40540 6967
rect 40500 6792 40552 6798
rect 40500 6734 40552 6740
rect 40788 6730 40816 7346
rect 41144 6928 41196 6934
rect 41144 6870 41196 6876
rect 40960 6792 41012 6798
rect 40960 6734 41012 6740
rect 41050 6760 41106 6769
rect 40684 6724 40736 6730
rect 40684 6666 40736 6672
rect 40776 6724 40828 6730
rect 40776 6666 40828 6672
rect 40696 5710 40724 6666
rect 40972 6458 41000 6734
rect 41156 6730 41184 6870
rect 41050 6695 41106 6704
rect 41144 6724 41196 6730
rect 40960 6452 41012 6458
rect 40960 6394 41012 6400
rect 41064 6254 41092 6695
rect 41144 6666 41196 6672
rect 41144 6384 41196 6390
rect 41248 6372 41276 7822
rect 41432 7206 41460 8502
rect 41512 8492 41564 8498
rect 41512 8434 41564 8440
rect 41524 7410 41552 8434
rect 41512 7404 41564 7410
rect 41512 7346 41564 7352
rect 41696 7404 41748 7410
rect 41696 7346 41748 7352
rect 41420 7200 41472 7206
rect 41420 7142 41472 7148
rect 41326 7032 41382 7041
rect 41326 6967 41382 6976
rect 41196 6344 41276 6372
rect 41144 6326 41196 6332
rect 41052 6248 41104 6254
rect 41052 6190 41104 6196
rect 41144 6248 41196 6254
rect 41144 6190 41196 6196
rect 40684 5704 40736 5710
rect 40684 5646 40736 5652
rect 41156 5574 41184 6190
rect 41248 5642 41276 6344
rect 41236 5636 41288 5642
rect 41236 5578 41288 5584
rect 41144 5568 41196 5574
rect 41144 5510 41196 5516
rect 40776 4684 40828 4690
rect 40776 4626 40828 4632
rect 40788 3942 40816 4626
rect 41248 4622 41276 5578
rect 41340 4758 41368 6967
rect 41432 5846 41460 7142
rect 41512 6860 41564 6866
rect 41512 6802 41564 6808
rect 41524 6769 41552 6802
rect 41510 6760 41566 6769
rect 41510 6695 41566 6704
rect 41512 6656 41564 6662
rect 41512 6598 41564 6604
rect 41604 6656 41656 6662
rect 41604 6598 41656 6604
rect 41524 6118 41552 6598
rect 41616 6390 41644 6598
rect 41708 6458 41736 7346
rect 41800 7342 41828 8774
rect 41892 8022 41920 14214
rect 41984 13734 42012 15150
rect 42156 15098 42208 15104
rect 42064 15020 42116 15026
rect 42064 14962 42116 14968
rect 42076 14618 42104 14962
rect 42156 14816 42208 14822
rect 42156 14758 42208 14764
rect 42064 14612 42116 14618
rect 42064 14554 42116 14560
rect 42168 14414 42196 14758
rect 42156 14408 42208 14414
rect 42156 14350 42208 14356
rect 42260 14362 42288 17054
rect 42340 16992 42392 16998
rect 42536 16980 42564 17682
rect 42628 17678 42656 19450
rect 42904 19446 42932 22879
rect 42996 21962 43024 23054
rect 43168 22568 43220 22574
rect 43166 22536 43168 22545
rect 43220 22536 43222 22545
rect 43166 22471 43222 22480
rect 43076 22092 43128 22098
rect 43076 22034 43128 22040
rect 43088 21962 43116 22034
rect 43364 21962 43392 24618
rect 43444 24608 43496 24614
rect 43444 24550 43496 24556
rect 43456 22982 43484 24550
rect 43548 24041 43576 26846
rect 43628 26852 43680 26858
rect 43628 26794 43680 26800
rect 43640 26382 43668 26794
rect 43732 26790 43760 27066
rect 43720 26784 43772 26790
rect 43720 26726 43772 26732
rect 43628 26376 43680 26382
rect 43628 26318 43680 26324
rect 43720 25152 43772 25158
rect 43720 25094 43772 25100
rect 43732 24614 43760 25094
rect 43916 24834 43944 37130
rect 44376 36378 44404 37130
rect 44468 36922 44496 39200
rect 45112 37466 45140 39200
rect 45100 37460 45152 37466
rect 45100 37402 45152 37408
rect 45756 36922 45784 39200
rect 46400 37466 46428 39200
rect 46388 37460 46440 37466
rect 46388 37402 46440 37408
rect 46112 37188 46164 37194
rect 46112 37130 46164 37136
rect 46124 36922 46152 37130
rect 47044 36922 47072 39200
rect 47688 36922 47716 39200
rect 48332 36922 48360 39200
rect 48976 36922 49004 39200
rect 49620 36922 49648 39200
rect 50264 36922 50292 39200
rect 50908 36922 50936 39200
rect 51552 36922 51580 39200
rect 52196 36922 52224 39200
rect 52840 36922 52868 39200
rect 53484 36922 53512 39200
rect 54128 36922 54156 39200
rect 54772 36922 54800 39200
rect 55416 36922 55444 39200
rect 56060 36922 56088 39200
rect 56704 36922 56732 39200
rect 57348 36922 57376 39200
rect 57992 36922 58020 39200
rect 58636 36922 58664 39200
rect 59280 36922 59308 39200
rect 59924 36922 59952 39200
rect 60568 36922 60596 39200
rect 61212 36922 61240 39200
rect 61856 36922 61884 39200
rect 62500 36922 62528 39200
rect 63144 36922 63172 39200
rect 63788 36922 63816 39200
rect 64432 36922 64460 39200
rect 65076 36922 65104 39200
rect 65720 37890 65748 39200
rect 66364 37890 66392 39200
rect 65536 37862 65748 37890
rect 66272 37862 66392 37890
rect 65536 36922 65564 37862
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 66272 37210 66300 37862
rect 66180 37182 66300 37210
rect 44456 36916 44508 36922
rect 44456 36858 44508 36864
rect 45744 36916 45796 36922
rect 45744 36858 45796 36864
rect 46112 36916 46164 36922
rect 46112 36858 46164 36864
rect 47032 36916 47084 36922
rect 47032 36858 47084 36864
rect 47676 36916 47728 36922
rect 47676 36858 47728 36864
rect 48320 36916 48372 36922
rect 48320 36858 48372 36864
rect 48964 36916 49016 36922
rect 48964 36858 49016 36864
rect 49608 36916 49660 36922
rect 49608 36858 49660 36864
rect 50252 36916 50304 36922
rect 50252 36858 50304 36864
rect 50896 36916 50948 36922
rect 50896 36858 50948 36864
rect 51540 36916 51592 36922
rect 51540 36858 51592 36864
rect 52184 36916 52236 36922
rect 52184 36858 52236 36864
rect 52828 36916 52880 36922
rect 52828 36858 52880 36864
rect 53472 36916 53524 36922
rect 53472 36858 53524 36864
rect 54116 36916 54168 36922
rect 54116 36858 54168 36864
rect 54760 36916 54812 36922
rect 54760 36858 54812 36864
rect 55404 36916 55456 36922
rect 55404 36858 55456 36864
rect 56048 36916 56100 36922
rect 56048 36858 56100 36864
rect 56692 36916 56744 36922
rect 56692 36858 56744 36864
rect 57336 36916 57388 36922
rect 57336 36858 57388 36864
rect 57980 36916 58032 36922
rect 57980 36858 58032 36864
rect 58624 36916 58676 36922
rect 58624 36858 58676 36864
rect 59268 36916 59320 36922
rect 59268 36858 59320 36864
rect 59912 36916 59964 36922
rect 59912 36858 59964 36864
rect 60556 36916 60608 36922
rect 60556 36858 60608 36864
rect 61200 36916 61252 36922
rect 61200 36858 61252 36864
rect 61844 36916 61896 36922
rect 61844 36858 61896 36864
rect 62488 36916 62540 36922
rect 62488 36858 62540 36864
rect 63132 36916 63184 36922
rect 63132 36858 63184 36864
rect 63776 36916 63828 36922
rect 63776 36858 63828 36864
rect 64420 36916 64472 36922
rect 64420 36858 64472 36864
rect 65064 36916 65116 36922
rect 65064 36858 65116 36864
rect 65524 36916 65576 36922
rect 66180 36904 66208 37182
rect 66314 37020 66622 37029
rect 66314 37018 66320 37020
rect 66376 37018 66400 37020
rect 66456 37018 66480 37020
rect 66536 37018 66560 37020
rect 66616 37018 66622 37020
rect 66376 36966 66378 37018
rect 66558 36966 66560 37018
rect 66314 36964 66320 36966
rect 66376 36964 66400 36966
rect 66456 36964 66480 36966
rect 66536 36964 66560 36966
rect 66616 36964 66622 36966
rect 66314 36955 66622 36964
rect 67008 36922 67036 39200
rect 67652 36922 67680 39200
rect 68296 36922 68324 39200
rect 68940 36922 68968 39200
rect 69584 36922 69612 39200
rect 70228 36922 70256 39200
rect 70872 36922 70900 39200
rect 71516 36922 71544 39200
rect 72160 36922 72188 39200
rect 72804 36922 72832 39200
rect 73448 36922 73476 39200
rect 66260 36916 66312 36922
rect 66180 36876 66260 36904
rect 65524 36858 65576 36864
rect 66260 36858 66312 36864
rect 66996 36916 67048 36922
rect 66996 36858 67048 36864
rect 67640 36916 67692 36922
rect 67640 36858 67692 36864
rect 68284 36916 68336 36922
rect 68284 36858 68336 36864
rect 68928 36916 68980 36922
rect 68928 36858 68980 36864
rect 69572 36916 69624 36922
rect 69572 36858 69624 36864
rect 70216 36916 70268 36922
rect 70216 36858 70268 36864
rect 70860 36916 70912 36922
rect 70860 36858 70912 36864
rect 71504 36916 71556 36922
rect 71504 36858 71556 36864
rect 72148 36916 72200 36922
rect 72148 36858 72200 36864
rect 72792 36916 72844 36922
rect 72792 36858 72844 36864
rect 73436 36916 73488 36922
rect 73436 36858 73488 36864
rect 44916 36848 44968 36854
rect 44916 36790 44968 36796
rect 44548 36576 44600 36582
rect 44548 36518 44600 36524
rect 44364 36372 44416 36378
rect 44364 36314 44416 36320
rect 44088 36168 44140 36174
rect 44088 36110 44140 36116
rect 44364 36168 44416 36174
rect 44364 36110 44416 36116
rect 44100 35154 44128 36110
rect 44272 36032 44324 36038
rect 44272 35974 44324 35980
rect 44284 35834 44312 35974
rect 44272 35828 44324 35834
rect 44272 35770 44324 35776
rect 44088 35148 44140 35154
rect 44088 35090 44140 35096
rect 44100 34950 44128 35090
rect 44272 35080 44324 35086
rect 44272 35022 44324 35028
rect 44088 34944 44140 34950
rect 44088 34886 44140 34892
rect 44284 34610 44312 35022
rect 44272 34604 44324 34610
rect 44272 34546 44324 34552
rect 44284 34406 44312 34546
rect 44272 34400 44324 34406
rect 44272 34342 44324 34348
rect 44284 33862 44312 34342
rect 44272 33856 44324 33862
rect 44272 33798 44324 33804
rect 44180 33652 44232 33658
rect 44180 33594 44232 33600
rect 44192 32434 44220 33594
rect 44284 33522 44312 33798
rect 44272 33516 44324 33522
rect 44272 33458 44324 33464
rect 44284 33114 44312 33458
rect 44272 33108 44324 33114
rect 44272 33050 44324 33056
rect 44376 32858 44404 36110
rect 44560 35698 44588 36518
rect 44548 35692 44600 35698
rect 44548 35634 44600 35640
rect 44732 35692 44784 35698
rect 44732 35634 44784 35640
rect 44560 35034 44588 35634
rect 44744 35290 44772 35634
rect 44732 35284 44784 35290
rect 44732 35226 44784 35232
rect 44560 35018 44680 35034
rect 44560 35012 44692 35018
rect 44560 35006 44640 35012
rect 44640 34954 44692 34960
rect 44652 34678 44680 34954
rect 44640 34672 44692 34678
rect 44640 34614 44692 34620
rect 44652 33318 44680 34614
rect 44744 33522 44772 35226
rect 44732 33516 44784 33522
rect 44732 33458 44784 33464
rect 44744 33386 44772 33458
rect 44732 33380 44784 33386
rect 44732 33322 44784 33328
rect 44640 33312 44692 33318
rect 44640 33254 44692 33260
rect 44284 32830 44404 32858
rect 44548 32904 44600 32910
rect 44652 32892 44680 33254
rect 44732 32904 44784 32910
rect 44652 32864 44732 32892
rect 44548 32846 44600 32852
rect 44732 32846 44784 32852
rect 44180 32428 44232 32434
rect 44180 32370 44232 32376
rect 44192 31958 44220 32370
rect 44180 31952 44232 31958
rect 44180 31894 44232 31900
rect 44284 31346 44312 32830
rect 44364 32768 44416 32774
rect 44364 32710 44416 32716
rect 44456 32768 44508 32774
rect 44456 32710 44508 32716
rect 44376 31822 44404 32710
rect 44468 32434 44496 32710
rect 44456 32428 44508 32434
rect 44560 32416 44588 32846
rect 44640 32428 44692 32434
rect 44560 32388 44640 32416
rect 44456 32370 44508 32376
rect 44640 32370 44692 32376
rect 44468 32026 44496 32370
rect 44456 32020 44508 32026
rect 44456 31962 44508 31968
rect 44548 31952 44600 31958
rect 44548 31894 44600 31900
rect 44364 31816 44416 31822
rect 44364 31758 44416 31764
rect 44560 31414 44588 31894
rect 44652 31890 44680 32370
rect 44640 31884 44692 31890
rect 44640 31826 44692 31832
rect 44548 31408 44600 31414
rect 44548 31350 44600 31356
rect 44272 31340 44324 31346
rect 44272 31282 44324 31288
rect 44364 29572 44416 29578
rect 44364 29514 44416 29520
rect 44376 29306 44404 29514
rect 44364 29300 44416 29306
rect 44364 29242 44416 29248
rect 44272 29164 44324 29170
rect 44272 29106 44324 29112
rect 43996 29096 44048 29102
rect 43996 29038 44048 29044
rect 44008 28994 44036 29038
rect 44284 28994 44312 29106
rect 44376 29102 44404 29242
rect 44560 29186 44588 31350
rect 44928 30326 44956 36790
rect 45008 36780 45060 36786
rect 45008 36722 45060 36728
rect 45928 36780 45980 36786
rect 45928 36722 45980 36728
rect 47768 36780 47820 36786
rect 47768 36722 47820 36728
rect 48780 36780 48832 36786
rect 48780 36722 48832 36728
rect 52920 36780 52972 36786
rect 52920 36722 52972 36728
rect 53288 36780 53340 36786
rect 53288 36722 53340 36728
rect 58072 36780 58124 36786
rect 58072 36722 58124 36728
rect 60648 36780 60700 36786
rect 60648 36722 60700 36728
rect 61016 36780 61068 36786
rect 61016 36722 61068 36728
rect 63132 36780 63184 36786
rect 63132 36722 63184 36728
rect 68284 36780 68336 36786
rect 68284 36722 68336 36728
rect 72240 36780 72292 36786
rect 72240 36722 72292 36728
rect 45020 36378 45048 36722
rect 45940 36394 45968 36722
rect 45008 36372 45060 36378
rect 45008 36314 45060 36320
rect 45848 36366 45968 36394
rect 47780 36378 47808 36722
rect 48792 36378 48820 36722
rect 52932 36378 52960 36722
rect 53300 36378 53328 36722
rect 58084 36378 58112 36722
rect 60660 36378 60688 36722
rect 61028 36378 61056 36722
rect 63144 36378 63172 36722
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 68296 36378 68324 36722
rect 72252 36378 72280 36722
rect 47768 36372 47820 36378
rect 45744 36236 45796 36242
rect 45744 36178 45796 36184
rect 45756 35766 45784 36178
rect 45744 35760 45796 35766
rect 45744 35702 45796 35708
rect 45756 34950 45784 35702
rect 45744 34944 45796 34950
rect 45744 34886 45796 34892
rect 45848 34746 45876 36366
rect 47768 36314 47820 36320
rect 48780 36372 48832 36378
rect 48780 36314 48832 36320
rect 52920 36372 52972 36378
rect 52920 36314 52972 36320
rect 53288 36372 53340 36378
rect 53288 36314 53340 36320
rect 58072 36372 58124 36378
rect 58072 36314 58124 36320
rect 60648 36372 60700 36378
rect 60648 36314 60700 36320
rect 61016 36372 61068 36378
rect 61016 36314 61068 36320
rect 63132 36372 63184 36378
rect 63132 36314 63184 36320
rect 68284 36372 68336 36378
rect 68284 36314 68336 36320
rect 72240 36372 72292 36378
rect 72240 36314 72292 36320
rect 46112 36168 46164 36174
rect 46112 36110 46164 36116
rect 46480 36168 46532 36174
rect 46480 36110 46532 36116
rect 45928 36032 45980 36038
rect 45928 35974 45980 35980
rect 45940 35766 45968 35974
rect 45928 35760 45980 35766
rect 45928 35702 45980 35708
rect 45928 35624 45980 35630
rect 45980 35572 46060 35578
rect 45928 35566 46060 35572
rect 45940 35550 46060 35566
rect 45836 34740 45888 34746
rect 45836 34682 45888 34688
rect 45100 34128 45152 34134
rect 45100 34070 45152 34076
rect 45112 33862 45140 34070
rect 45100 33856 45152 33862
rect 45100 33798 45152 33804
rect 45112 33590 45140 33798
rect 45928 33652 45980 33658
rect 45928 33594 45980 33600
rect 45100 33584 45152 33590
rect 45100 33526 45152 33532
rect 45192 33380 45244 33386
rect 45192 33322 45244 33328
rect 45204 33114 45232 33322
rect 45192 33108 45244 33114
rect 45192 33050 45244 33056
rect 45376 33040 45428 33046
rect 45376 32982 45428 32988
rect 45192 32972 45244 32978
rect 45192 32914 45244 32920
rect 45204 32570 45232 32914
rect 45388 32910 45416 32982
rect 45940 32978 45968 33594
rect 46032 33454 46060 35550
rect 46124 35290 46152 36110
rect 46492 35834 46520 36110
rect 66314 35932 66622 35941
rect 66314 35930 66320 35932
rect 66376 35930 66400 35932
rect 66456 35930 66480 35932
rect 66536 35930 66560 35932
rect 66616 35930 66622 35932
rect 66376 35878 66378 35930
rect 66558 35878 66560 35930
rect 66314 35876 66320 35878
rect 66376 35876 66400 35878
rect 66456 35876 66480 35878
rect 66536 35876 66560 35878
rect 66616 35876 66622 35878
rect 66314 35867 66622 35876
rect 46480 35828 46532 35834
rect 46480 35770 46532 35776
rect 46112 35284 46164 35290
rect 46112 35226 46164 35232
rect 46492 35154 46520 35770
rect 48780 35488 48832 35494
rect 48780 35430 48832 35436
rect 46480 35148 46532 35154
rect 46480 35090 46532 35096
rect 46848 35080 46900 35086
rect 46848 35022 46900 35028
rect 46112 34604 46164 34610
rect 46112 34546 46164 34552
rect 46124 33658 46152 34546
rect 46112 33652 46164 33658
rect 46112 33594 46164 33600
rect 46204 33652 46256 33658
rect 46204 33594 46256 33600
rect 46020 33448 46072 33454
rect 46020 33390 46072 33396
rect 46032 33318 46060 33390
rect 46020 33312 46072 33318
rect 46020 33254 46072 33260
rect 45928 32972 45980 32978
rect 45928 32914 45980 32920
rect 45376 32904 45428 32910
rect 45376 32846 45428 32852
rect 45192 32564 45244 32570
rect 45192 32506 45244 32512
rect 45940 32502 45968 32914
rect 46020 32904 46072 32910
rect 46020 32846 46072 32852
rect 46032 32502 46060 32846
rect 46216 32842 46244 33594
rect 46860 33522 46888 35022
rect 48792 33590 48820 35430
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 66314 34844 66622 34853
rect 66314 34842 66320 34844
rect 66376 34842 66400 34844
rect 66456 34842 66480 34844
rect 66536 34842 66560 34844
rect 66616 34842 66622 34844
rect 66376 34790 66378 34842
rect 66558 34790 66560 34842
rect 66314 34788 66320 34790
rect 66376 34788 66400 34790
rect 66456 34788 66480 34790
rect 66536 34788 66560 34790
rect 66616 34788 66622 34790
rect 66314 34779 66622 34788
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 66314 33756 66622 33765
rect 66314 33754 66320 33756
rect 66376 33754 66400 33756
rect 66456 33754 66480 33756
rect 66536 33754 66560 33756
rect 66616 33754 66622 33756
rect 66376 33702 66378 33754
rect 66558 33702 66560 33754
rect 66314 33700 66320 33702
rect 66376 33700 66400 33702
rect 66456 33700 66480 33702
rect 66536 33700 66560 33702
rect 66616 33700 66622 33702
rect 66314 33691 66622 33700
rect 47676 33584 47728 33590
rect 47676 33526 47728 33532
rect 48780 33584 48832 33590
rect 48780 33526 48832 33532
rect 46388 33516 46440 33522
rect 46388 33458 46440 33464
rect 46848 33516 46900 33522
rect 46848 33458 46900 33464
rect 46204 32836 46256 32842
rect 46204 32778 46256 32784
rect 46112 32768 46164 32774
rect 46112 32710 46164 32716
rect 45560 32496 45612 32502
rect 45560 32438 45612 32444
rect 45928 32496 45980 32502
rect 45928 32438 45980 32444
rect 46020 32496 46072 32502
rect 46020 32438 46072 32444
rect 45572 32230 45600 32438
rect 45560 32224 45612 32230
rect 45560 32166 45612 32172
rect 45376 31816 45428 31822
rect 45376 31758 45428 31764
rect 45100 31680 45152 31686
rect 45100 31622 45152 31628
rect 45112 31142 45140 31622
rect 45100 31136 45152 31142
rect 45100 31078 45152 31084
rect 45284 31136 45336 31142
rect 45284 31078 45336 31084
rect 45296 30666 45324 31078
rect 45284 30660 45336 30666
rect 45284 30602 45336 30608
rect 44916 30320 44968 30326
rect 44916 30262 44968 30268
rect 44824 30252 44876 30258
rect 44824 30194 44876 30200
rect 44836 30054 44864 30194
rect 44824 30048 44876 30054
rect 44822 30016 44824 30025
rect 44876 30016 44878 30025
rect 44822 29951 44878 29960
rect 44560 29158 44680 29186
rect 44364 29096 44416 29102
rect 44364 29038 44416 29044
rect 44008 28966 44312 28994
rect 44548 29028 44600 29034
rect 44548 28970 44600 28976
rect 44008 28490 44036 28966
rect 43996 28484 44048 28490
rect 43996 28426 44048 28432
rect 44180 28076 44232 28082
rect 44180 28018 44232 28024
rect 44192 27538 44220 28018
rect 44180 27532 44232 27538
rect 44180 27474 44232 27480
rect 44192 27010 44220 27474
rect 44192 26982 44312 27010
rect 44284 26926 44312 26982
rect 44272 26920 44324 26926
rect 44272 26862 44324 26868
rect 44180 26852 44232 26858
rect 44180 26794 44232 26800
rect 44088 26512 44140 26518
rect 44088 26454 44140 26460
rect 43824 24806 43944 24834
rect 44100 24818 44128 26454
rect 44192 25770 44220 26794
rect 44456 26308 44508 26314
rect 44456 26250 44508 26256
rect 44180 25764 44232 25770
rect 44180 25706 44232 25712
rect 44364 25696 44416 25702
rect 44364 25638 44416 25644
rect 44270 24984 44326 24993
rect 44376 24954 44404 25638
rect 44270 24919 44326 24928
rect 44364 24948 44416 24954
rect 44088 24812 44140 24818
rect 43720 24608 43772 24614
rect 43720 24550 43772 24556
rect 43534 24032 43590 24041
rect 43534 23967 43590 23976
rect 43732 23730 43760 24550
rect 43824 23866 43852 24806
rect 44088 24754 44140 24760
rect 43904 24744 43956 24750
rect 43904 24686 43956 24692
rect 43916 24410 43944 24686
rect 44100 24614 44128 24754
rect 44088 24608 44140 24614
rect 44088 24550 44140 24556
rect 43904 24404 43956 24410
rect 43904 24346 43956 24352
rect 44100 24120 44128 24550
rect 44180 24132 44232 24138
rect 44100 24092 44180 24120
rect 44180 24074 44232 24080
rect 43812 23860 43864 23866
rect 43812 23802 43864 23808
rect 43720 23724 43772 23730
rect 43720 23666 43772 23672
rect 44180 23724 44232 23730
rect 44180 23666 44232 23672
rect 43628 23656 43680 23662
rect 43628 23598 43680 23604
rect 43640 23118 43668 23598
rect 43628 23112 43680 23118
rect 43732 23100 43760 23666
rect 44192 23610 44220 23666
rect 44100 23582 44220 23610
rect 44100 23186 44128 23582
rect 44180 23520 44232 23526
rect 44180 23462 44232 23468
rect 44088 23180 44140 23186
rect 44088 23122 44140 23128
rect 43812 23112 43864 23118
rect 43732 23072 43812 23100
rect 43628 23054 43680 23060
rect 43812 23054 43864 23060
rect 43904 23112 43956 23118
rect 43904 23054 43956 23060
rect 43444 22976 43496 22982
rect 43444 22918 43496 22924
rect 43536 22568 43588 22574
rect 43536 22510 43588 22516
rect 43548 21962 43576 22510
rect 43916 22098 43944 23054
rect 44192 22778 44220 23462
rect 44284 23186 44312 24919
rect 44364 24890 44416 24896
rect 44376 24206 44404 24890
rect 44468 24818 44496 26250
rect 44560 25906 44588 28970
rect 44548 25900 44600 25906
rect 44548 25842 44600 25848
rect 44456 24812 44508 24818
rect 44456 24754 44508 24760
rect 44364 24200 44416 24206
rect 44364 24142 44416 24148
rect 44364 24064 44416 24070
rect 44364 24006 44416 24012
rect 44376 23730 44404 24006
rect 44468 23730 44496 24754
rect 44652 23798 44680 29158
rect 45100 29164 45152 29170
rect 45100 29106 45152 29112
rect 45112 28558 45140 29106
rect 45100 28552 45152 28558
rect 45100 28494 45152 28500
rect 45112 28082 45140 28494
rect 45284 28416 45336 28422
rect 45284 28358 45336 28364
rect 44732 28076 44784 28082
rect 44732 28018 44784 28024
rect 45100 28076 45152 28082
rect 45100 28018 45152 28024
rect 44744 27946 44772 28018
rect 44732 27940 44784 27946
rect 44732 27882 44784 27888
rect 44744 26382 44772 27882
rect 45296 26994 45324 28358
rect 45284 26988 45336 26994
rect 45284 26930 45336 26936
rect 44824 26920 44876 26926
rect 44824 26862 44876 26868
rect 44732 26376 44784 26382
rect 44732 26318 44784 26324
rect 44744 25770 44772 26318
rect 44836 26246 44864 26862
rect 45008 26376 45060 26382
rect 45008 26318 45060 26324
rect 44824 26240 44876 26246
rect 44824 26182 44876 26188
rect 44836 25906 44864 26182
rect 45020 25974 45048 26318
rect 45296 26246 45324 26930
rect 45284 26240 45336 26246
rect 45284 26182 45336 26188
rect 45008 25968 45060 25974
rect 45008 25910 45060 25916
rect 45296 25906 45324 26182
rect 44824 25900 44876 25906
rect 44824 25842 44876 25848
rect 45284 25900 45336 25906
rect 45284 25842 45336 25848
rect 44732 25764 44784 25770
rect 44732 25706 44784 25712
rect 44836 24818 44864 25842
rect 45296 24818 45324 25842
rect 44824 24812 44876 24818
rect 44824 24754 44876 24760
rect 45284 24812 45336 24818
rect 45284 24754 45336 24760
rect 45296 24342 45324 24754
rect 45284 24336 45336 24342
rect 45284 24278 45336 24284
rect 45296 23798 45324 24278
rect 44640 23792 44692 23798
rect 44640 23734 44692 23740
rect 45284 23792 45336 23798
rect 45284 23734 45336 23740
rect 44364 23724 44416 23730
rect 44364 23666 44416 23672
rect 44456 23724 44508 23730
rect 44456 23666 44508 23672
rect 44272 23180 44324 23186
rect 44272 23122 44324 23128
rect 44284 23089 44312 23122
rect 44270 23080 44326 23089
rect 44270 23015 44326 23024
rect 44376 22794 44404 23666
rect 44456 23520 44508 23526
rect 44456 23462 44508 23468
rect 44180 22772 44232 22778
rect 44180 22714 44232 22720
rect 44284 22766 44404 22794
rect 44284 22574 44312 22766
rect 44364 22704 44416 22710
rect 44364 22646 44416 22652
rect 44272 22568 44324 22574
rect 44272 22510 44324 22516
rect 44284 22234 44312 22510
rect 44272 22228 44324 22234
rect 44272 22170 44324 22176
rect 43996 22160 44048 22166
rect 43994 22128 43996 22137
rect 44048 22128 44050 22137
rect 43904 22092 43956 22098
rect 43994 22063 44050 22072
rect 43904 22034 43956 22040
rect 42984 21956 43036 21962
rect 42984 21898 43036 21904
rect 43076 21956 43128 21962
rect 43076 21898 43128 21904
rect 43352 21956 43404 21962
rect 43352 21898 43404 21904
rect 43536 21956 43588 21962
rect 43536 21898 43588 21904
rect 43904 21956 43956 21962
rect 43904 21898 43956 21904
rect 42996 20942 43024 21898
rect 42984 20936 43036 20942
rect 42984 20878 43036 20884
rect 42996 19922 43024 20878
rect 43364 20874 43392 21898
rect 43352 20868 43404 20874
rect 43352 20810 43404 20816
rect 43916 20602 43944 21898
rect 43904 20596 43956 20602
rect 43904 20538 43956 20544
rect 42984 19916 43036 19922
rect 42984 19858 43036 19864
rect 43444 19508 43496 19514
rect 43444 19450 43496 19456
rect 43628 19508 43680 19514
rect 43628 19450 43680 19456
rect 42892 19440 42944 19446
rect 42892 19382 42944 19388
rect 43260 19304 43312 19310
rect 43260 19246 43312 19252
rect 43272 18698 43300 19246
rect 43260 18692 43312 18698
rect 43260 18634 43312 18640
rect 43168 18624 43220 18630
rect 43168 18566 43220 18572
rect 42984 18420 43036 18426
rect 42984 18362 43036 18368
rect 42708 18284 42760 18290
rect 42708 18226 42760 18232
rect 42616 17672 42668 17678
rect 42616 17614 42668 17620
rect 42720 17270 42748 18226
rect 42800 18216 42852 18222
rect 42800 18158 42852 18164
rect 42708 17264 42760 17270
rect 42708 17206 42760 17212
rect 42392 16952 42564 16980
rect 42340 16934 42392 16940
rect 42340 14612 42392 14618
rect 42340 14554 42392 14560
rect 42352 14482 42380 14554
rect 42340 14476 42392 14482
rect 42340 14418 42392 14424
rect 42260 14334 42380 14362
rect 42248 14272 42300 14278
rect 42248 14214 42300 14220
rect 42260 13802 42288 14214
rect 42248 13796 42300 13802
rect 42248 13738 42300 13744
rect 41972 13728 42024 13734
rect 41972 13670 42024 13676
rect 42352 13530 42380 14334
rect 42340 13524 42392 13530
rect 42340 13466 42392 13472
rect 42248 12844 42300 12850
rect 42248 12786 42300 12792
rect 42156 12776 42208 12782
rect 42156 12718 42208 12724
rect 42168 12442 42196 12718
rect 42156 12436 42208 12442
rect 42156 12378 42208 12384
rect 42168 12306 42196 12378
rect 42156 12300 42208 12306
rect 42156 12242 42208 12248
rect 42260 11354 42288 12786
rect 42248 11348 42300 11354
rect 42248 11290 42300 11296
rect 42064 11144 42116 11150
rect 42064 11086 42116 11092
rect 41972 11008 42024 11014
rect 41972 10950 42024 10956
rect 41984 9994 42012 10950
rect 42076 10810 42104 11086
rect 42248 11008 42300 11014
rect 42248 10950 42300 10956
rect 42064 10804 42116 10810
rect 42064 10746 42116 10752
rect 42064 10668 42116 10674
rect 42064 10610 42116 10616
rect 41972 9988 42024 9994
rect 41972 9930 42024 9936
rect 41972 9376 42024 9382
rect 41972 9318 42024 9324
rect 41984 8974 42012 9318
rect 42076 8974 42104 10610
rect 42260 10606 42288 10950
rect 42248 10600 42300 10606
rect 42248 10542 42300 10548
rect 41972 8968 42024 8974
rect 41972 8910 42024 8916
rect 42064 8968 42116 8974
rect 42064 8910 42116 8916
rect 41984 8090 42012 8910
rect 42076 8294 42104 8910
rect 42064 8288 42116 8294
rect 42064 8230 42116 8236
rect 41972 8084 42024 8090
rect 41972 8026 42024 8032
rect 41880 8016 41932 8022
rect 41880 7958 41932 7964
rect 41880 7880 41932 7886
rect 41880 7822 41932 7828
rect 41788 7336 41840 7342
rect 41788 7278 41840 7284
rect 41696 6452 41748 6458
rect 41696 6394 41748 6400
rect 41604 6384 41656 6390
rect 41604 6326 41656 6332
rect 41512 6112 41564 6118
rect 41512 6054 41564 6060
rect 41420 5840 41472 5846
rect 41420 5782 41472 5788
rect 41708 5710 41736 6394
rect 41696 5704 41748 5710
rect 41696 5646 41748 5652
rect 41800 5574 41828 7278
rect 41892 5710 41920 7822
rect 41984 7478 42012 8026
rect 41972 7472 42024 7478
rect 41972 7414 42024 7420
rect 42260 6186 42288 10542
rect 42340 9580 42392 9586
rect 42340 9522 42392 9528
rect 42352 8838 42380 9522
rect 42340 8832 42392 8838
rect 42340 8774 42392 8780
rect 42338 8528 42394 8537
rect 42338 8463 42340 8472
rect 42392 8463 42394 8472
rect 42340 8434 42392 8440
rect 42340 7812 42392 7818
rect 42340 7754 42392 7760
rect 42352 7410 42380 7754
rect 42340 7404 42392 7410
rect 42340 7346 42392 7352
rect 42444 6866 42472 16952
rect 42812 16658 42840 18158
rect 42892 18080 42944 18086
rect 42892 18022 42944 18028
rect 42904 17746 42932 18022
rect 42892 17740 42944 17746
rect 42892 17682 42944 17688
rect 42996 17202 43024 18362
rect 43076 18216 43128 18222
rect 43076 18158 43128 18164
rect 43088 17338 43116 18158
rect 43180 17678 43208 18566
rect 43168 17672 43220 17678
rect 43166 17640 43168 17649
rect 43220 17640 43222 17649
rect 43166 17575 43222 17584
rect 43168 17536 43220 17542
rect 43168 17478 43220 17484
rect 43076 17332 43128 17338
rect 43076 17274 43128 17280
rect 42984 17196 43036 17202
rect 42984 17138 43036 17144
rect 43180 16794 43208 17478
rect 43168 16788 43220 16794
rect 43168 16730 43220 16736
rect 42800 16652 42852 16658
rect 42800 16594 42852 16600
rect 42616 16448 42668 16454
rect 42616 16390 42668 16396
rect 42524 16244 42576 16250
rect 42524 16186 42576 16192
rect 42536 13462 42564 16186
rect 42628 15706 42656 16390
rect 42616 15700 42668 15706
rect 42616 15642 42668 15648
rect 42628 15434 42656 15642
rect 42616 15428 42668 15434
rect 42616 15370 42668 15376
rect 42984 15020 43036 15026
rect 42984 14962 43036 14968
rect 42996 14793 43024 14962
rect 42982 14784 43038 14793
rect 42982 14719 43038 14728
rect 43076 14612 43128 14618
rect 43076 14554 43128 14560
rect 42800 14408 42852 14414
rect 42800 14350 42852 14356
rect 42708 13524 42760 13530
rect 42708 13466 42760 13472
rect 42524 13456 42576 13462
rect 42524 13398 42576 13404
rect 42524 12164 42576 12170
rect 42524 12106 42576 12112
rect 42536 11830 42564 12106
rect 42524 11824 42576 11830
rect 42524 11766 42576 11772
rect 42720 9602 42748 13466
rect 42812 12374 42840 14350
rect 42892 13320 42944 13326
rect 42892 13262 42944 13268
rect 42904 12442 42932 13262
rect 42984 13184 43036 13190
rect 42984 13126 43036 13132
rect 42996 12918 43024 13126
rect 42984 12912 43036 12918
rect 42984 12854 43036 12860
rect 42892 12436 42944 12442
rect 42892 12378 42944 12384
rect 42800 12368 42852 12374
rect 42800 12310 42852 12316
rect 42536 9574 42748 9602
rect 42800 9580 42852 9586
rect 42536 7546 42564 9574
rect 42800 9522 42852 9528
rect 42708 9512 42760 9518
rect 42708 9454 42760 9460
rect 42616 9172 42668 9178
rect 42616 9114 42668 9120
rect 42628 9042 42656 9114
rect 42616 9036 42668 9042
rect 42616 8978 42668 8984
rect 42720 8498 42748 9454
rect 42812 8634 42840 9522
rect 42890 9344 42946 9353
rect 42890 9279 42946 9288
rect 42904 9178 42932 9279
rect 42892 9172 42944 9178
rect 42892 9114 42944 9120
rect 42800 8628 42852 8634
rect 42800 8570 42852 8576
rect 42890 8528 42946 8537
rect 42616 8492 42668 8498
rect 42616 8434 42668 8440
rect 42708 8492 42760 8498
rect 42890 8463 42892 8472
rect 42708 8434 42760 8440
rect 42944 8463 42946 8472
rect 42984 8492 43036 8498
rect 42892 8434 42944 8440
rect 42984 8434 43036 8440
rect 42628 8090 42656 8434
rect 42708 8288 42760 8294
rect 42708 8230 42760 8236
rect 42616 8084 42668 8090
rect 42616 8026 42668 8032
rect 42616 7812 42668 7818
rect 42616 7754 42668 7760
rect 42524 7540 42576 7546
rect 42524 7482 42576 7488
rect 42432 6860 42484 6866
rect 42432 6802 42484 6808
rect 42444 6458 42472 6802
rect 42432 6452 42484 6458
rect 42432 6394 42484 6400
rect 42248 6180 42300 6186
rect 42248 6122 42300 6128
rect 42536 6118 42564 7482
rect 42628 7410 42656 7754
rect 42720 7750 42748 8230
rect 42708 7744 42760 7750
rect 42708 7686 42760 7692
rect 42616 7404 42668 7410
rect 42616 7346 42668 7352
rect 42524 6112 42576 6118
rect 42524 6054 42576 6060
rect 41880 5704 41932 5710
rect 41880 5646 41932 5652
rect 41420 5568 41472 5574
rect 41420 5510 41472 5516
rect 41788 5568 41840 5574
rect 41788 5510 41840 5516
rect 41328 4752 41380 4758
rect 41328 4694 41380 4700
rect 41236 4616 41288 4622
rect 41236 4558 41288 4564
rect 41144 4140 41196 4146
rect 41432 4128 41460 5510
rect 41800 5234 41828 5510
rect 41892 5302 41920 5646
rect 42628 5370 42656 7346
rect 42800 6792 42852 6798
rect 42800 6734 42852 6740
rect 42812 6254 42840 6734
rect 42800 6248 42852 6254
rect 42800 6190 42852 6196
rect 42616 5364 42668 5370
rect 42616 5306 42668 5312
rect 41880 5296 41932 5302
rect 41880 5238 41932 5244
rect 41788 5228 41840 5234
rect 41788 5170 41840 5176
rect 41800 4214 41828 5170
rect 41972 4752 42024 4758
rect 41972 4694 42024 4700
rect 41984 4214 42012 4694
rect 42628 4214 42656 5306
rect 42812 4622 42840 6190
rect 42892 5296 42944 5302
rect 42892 5238 42944 5244
rect 42800 4616 42852 4622
rect 42800 4558 42852 4564
rect 41788 4208 41840 4214
rect 41788 4150 41840 4156
rect 41972 4208 42024 4214
rect 41972 4150 42024 4156
rect 42616 4208 42668 4214
rect 42616 4150 42668 4156
rect 41196 4100 41460 4128
rect 41144 4082 41196 4088
rect 40880 4010 41552 4026
rect 40868 4004 41552 4010
rect 40920 3998 41552 4004
rect 40868 3946 40920 3952
rect 41524 3942 41552 3998
rect 40776 3936 40828 3942
rect 40776 3878 40828 3884
rect 41420 3936 41472 3942
rect 41420 3878 41472 3884
rect 41512 3936 41564 3942
rect 41512 3878 41564 3884
rect 41432 3466 41460 3878
rect 42812 3602 42840 4558
rect 42904 4146 42932 5238
rect 42996 5216 43024 8434
rect 43088 8090 43116 14554
rect 43272 10044 43300 18634
rect 43352 18624 43404 18630
rect 43352 18566 43404 18572
rect 43364 18358 43392 18566
rect 43352 18352 43404 18358
rect 43352 18294 43404 18300
rect 43456 17882 43484 19450
rect 43536 18760 43588 18766
rect 43536 18702 43588 18708
rect 43444 17876 43496 17882
rect 43444 17818 43496 17824
rect 43352 17672 43404 17678
rect 43456 17660 43484 17818
rect 43404 17632 43484 17660
rect 43352 17614 43404 17620
rect 43444 17536 43496 17542
rect 43444 17478 43496 17484
rect 43456 17202 43484 17478
rect 43548 17241 43576 18702
rect 43534 17232 43590 17241
rect 43444 17196 43496 17202
rect 43534 17167 43590 17176
rect 43444 17138 43496 17144
rect 43640 16998 43668 19450
rect 43720 19372 43772 19378
rect 44008 19334 44036 22063
rect 44272 21888 44324 21894
rect 44272 21830 44324 21836
rect 44088 20868 44140 20874
rect 44088 20810 44140 20816
rect 44100 20534 44128 20810
rect 44284 20806 44312 21830
rect 44272 20800 44324 20806
rect 44272 20742 44324 20748
rect 44376 20534 44404 22646
rect 44468 22409 44496 23462
rect 44652 23100 44680 23734
rect 45388 23254 45416 31758
rect 45940 31754 45968 32438
rect 46124 32230 46152 32710
rect 46216 32298 46244 32778
rect 46400 32570 46428 33458
rect 46860 33046 46888 33458
rect 47688 33318 47716 33526
rect 47768 33448 47820 33454
rect 47768 33390 47820 33396
rect 48044 33448 48096 33454
rect 48044 33390 48096 33396
rect 47492 33312 47544 33318
rect 47492 33254 47544 33260
rect 47676 33312 47728 33318
rect 47676 33254 47728 33260
rect 46848 33040 46900 33046
rect 46848 32982 46900 32988
rect 47504 32910 47532 33254
rect 47688 32910 47716 33254
rect 47780 32978 47808 33390
rect 48056 33114 48084 33390
rect 48044 33108 48096 33114
rect 48044 33050 48096 33056
rect 48792 32978 48820 33526
rect 49608 33312 49660 33318
rect 49608 33254 49660 33260
rect 49620 32978 49648 33254
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 47768 32972 47820 32978
rect 47768 32914 47820 32920
rect 48780 32972 48832 32978
rect 48780 32914 48832 32920
rect 49608 32972 49660 32978
rect 49608 32914 49660 32920
rect 47216 32904 47268 32910
rect 47216 32846 47268 32852
rect 47308 32904 47360 32910
rect 47308 32846 47360 32852
rect 47492 32904 47544 32910
rect 47492 32846 47544 32852
rect 47584 32904 47636 32910
rect 47584 32846 47636 32852
rect 47676 32904 47728 32910
rect 47676 32846 47728 32852
rect 46572 32768 46624 32774
rect 46572 32710 46624 32716
rect 46388 32564 46440 32570
rect 46388 32506 46440 32512
rect 46584 32366 46612 32710
rect 47228 32502 47256 32846
rect 47216 32496 47268 32502
rect 47216 32438 47268 32444
rect 46572 32360 46624 32366
rect 46572 32302 46624 32308
rect 46204 32292 46256 32298
rect 46204 32234 46256 32240
rect 46112 32224 46164 32230
rect 46112 32166 46164 32172
rect 46388 32224 46440 32230
rect 46388 32166 46440 32172
rect 46400 32026 46428 32166
rect 46388 32020 46440 32026
rect 46388 31962 46440 31968
rect 45940 31748 46164 31754
rect 45940 31726 46112 31748
rect 46112 31690 46164 31696
rect 46296 31748 46348 31754
rect 46296 31690 46348 31696
rect 46124 31278 46152 31690
rect 46308 31346 46336 31690
rect 46400 31346 46428 31962
rect 46584 31754 46612 32302
rect 47320 32230 47348 32846
rect 47596 32570 47624 32846
rect 48792 32842 48820 32914
rect 48780 32836 48832 32842
rect 48780 32778 48832 32784
rect 47584 32564 47636 32570
rect 47584 32506 47636 32512
rect 47768 32428 47820 32434
rect 47768 32370 47820 32376
rect 47308 32224 47360 32230
rect 47308 32166 47360 32172
rect 47124 32020 47176 32026
rect 47124 31962 47176 31968
rect 46572 31748 46624 31754
rect 46572 31690 46624 31696
rect 47136 31346 47164 31962
rect 46296 31340 46348 31346
rect 46296 31282 46348 31288
rect 46388 31340 46440 31346
rect 46388 31282 46440 31288
rect 46572 31340 46624 31346
rect 46572 31282 46624 31288
rect 47124 31340 47176 31346
rect 47124 31282 47176 31288
rect 46112 31272 46164 31278
rect 46112 31214 46164 31220
rect 46584 30870 46612 31282
rect 47320 31278 47348 32166
rect 47780 32026 47808 32370
rect 48044 32360 48096 32366
rect 48044 32302 48096 32308
rect 48056 32230 48084 32302
rect 48044 32224 48096 32230
rect 48044 32166 48096 32172
rect 47768 32020 47820 32026
rect 47768 31962 47820 31968
rect 46756 31272 46808 31278
rect 46756 31214 46808 31220
rect 47308 31272 47360 31278
rect 47308 31214 47360 31220
rect 46768 30938 46796 31214
rect 47216 31136 47268 31142
rect 47216 31078 47268 31084
rect 46756 30932 46808 30938
rect 46756 30874 46808 30880
rect 46572 30864 46624 30870
rect 46572 30806 46624 30812
rect 47228 30802 47256 31078
rect 47216 30796 47268 30802
rect 47216 30738 47268 30744
rect 46940 30660 46992 30666
rect 46940 30602 46992 30608
rect 46952 30054 46980 30602
rect 48792 30598 48820 32778
rect 49792 32768 49844 32774
rect 49792 32710 49844 32716
rect 49804 32434 49832 32710
rect 66314 32668 66622 32677
rect 66314 32666 66320 32668
rect 66376 32666 66400 32668
rect 66456 32666 66480 32668
rect 66536 32666 66560 32668
rect 66616 32666 66622 32668
rect 66376 32614 66378 32666
rect 66558 32614 66560 32666
rect 66314 32612 66320 32614
rect 66376 32612 66400 32614
rect 66456 32612 66480 32614
rect 66536 32612 66560 32614
rect 66616 32612 66622 32614
rect 66314 32603 66622 32612
rect 49792 32428 49844 32434
rect 49792 32370 49844 32376
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 66314 31580 66622 31589
rect 66314 31578 66320 31580
rect 66376 31578 66400 31580
rect 66456 31578 66480 31580
rect 66536 31578 66560 31580
rect 66616 31578 66622 31580
rect 66376 31526 66378 31578
rect 66558 31526 66560 31578
rect 66314 31524 66320 31526
rect 66376 31524 66400 31526
rect 66456 31524 66480 31526
rect 66536 31524 66560 31526
rect 66616 31524 66622 31526
rect 66314 31515 66622 31524
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 48228 30592 48280 30598
rect 48228 30534 48280 30540
rect 48780 30592 48832 30598
rect 48780 30534 48832 30540
rect 48240 30054 48268 30534
rect 66314 30492 66622 30501
rect 66314 30490 66320 30492
rect 66376 30490 66400 30492
rect 66456 30490 66480 30492
rect 66536 30490 66560 30492
rect 66616 30490 66622 30492
rect 66376 30438 66378 30490
rect 66558 30438 66560 30490
rect 66314 30436 66320 30438
rect 66376 30436 66400 30438
rect 66456 30436 66480 30438
rect 66536 30436 66560 30438
rect 66616 30436 66622 30438
rect 66314 30427 66622 30436
rect 46940 30048 46992 30054
rect 46940 29990 46992 29996
rect 48228 30048 48280 30054
rect 48228 29990 48280 29996
rect 47676 29232 47728 29238
rect 47676 29174 47728 29180
rect 46204 29164 46256 29170
rect 46204 29106 46256 29112
rect 47492 29164 47544 29170
rect 47492 29106 47544 29112
rect 45836 29096 45888 29102
rect 45836 29038 45888 29044
rect 46020 29096 46072 29102
rect 46020 29038 46072 29044
rect 45468 28620 45520 28626
rect 45468 28562 45520 28568
rect 45480 28422 45508 28562
rect 45468 28416 45520 28422
rect 45468 28358 45520 28364
rect 45468 28144 45520 28150
rect 45468 28086 45520 28092
rect 45480 26382 45508 28086
rect 45848 27878 45876 29038
rect 46032 28558 46060 29038
rect 46020 28552 46072 28558
rect 46020 28494 46072 28500
rect 46216 28490 46244 29106
rect 46480 28960 46532 28966
rect 46480 28902 46532 28908
rect 46492 28558 46520 28902
rect 46572 28688 46624 28694
rect 46572 28630 46624 28636
rect 46480 28552 46532 28558
rect 46480 28494 46532 28500
rect 46204 28484 46256 28490
rect 46204 28426 46256 28432
rect 45928 28212 45980 28218
rect 45928 28154 45980 28160
rect 45836 27872 45888 27878
rect 45836 27814 45888 27820
rect 45848 27470 45876 27814
rect 45836 27464 45888 27470
rect 45836 27406 45888 27412
rect 45848 26450 45876 27406
rect 45940 27334 45968 28154
rect 46584 28082 46612 28630
rect 47504 28626 47532 29106
rect 47492 28620 47544 28626
rect 47492 28562 47544 28568
rect 46664 28484 46716 28490
rect 46664 28426 46716 28432
rect 46676 28150 46704 28426
rect 47504 28218 47532 28562
rect 47492 28212 47544 28218
rect 47492 28154 47544 28160
rect 46664 28144 46716 28150
rect 46664 28086 46716 28092
rect 46572 28076 46624 28082
rect 46572 28018 46624 28024
rect 46112 28008 46164 28014
rect 46112 27950 46164 27956
rect 46124 27878 46152 27950
rect 46020 27872 46072 27878
rect 46020 27814 46072 27820
rect 46112 27872 46164 27878
rect 46112 27814 46164 27820
rect 45928 27328 45980 27334
rect 45928 27270 45980 27276
rect 45940 26858 45968 27270
rect 46032 27130 46060 27814
rect 46020 27124 46072 27130
rect 46020 27066 46072 27072
rect 45928 26852 45980 26858
rect 45928 26794 45980 26800
rect 46032 26518 46060 27066
rect 46020 26512 46072 26518
rect 46020 26454 46072 26460
rect 45836 26444 45888 26450
rect 45836 26386 45888 26392
rect 45468 26376 45520 26382
rect 45468 26318 45520 26324
rect 45480 25974 45508 26318
rect 46124 26314 46152 27814
rect 46480 26376 46532 26382
rect 46480 26318 46532 26324
rect 46112 26308 46164 26314
rect 46112 26250 46164 26256
rect 46492 26042 46520 26318
rect 46480 26036 46532 26042
rect 46480 25978 46532 25984
rect 45468 25968 45520 25974
rect 45468 25910 45520 25916
rect 46584 25294 46612 28018
rect 47688 27878 47716 29174
rect 48240 28422 48268 29990
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 66314 29404 66622 29413
rect 66314 29402 66320 29404
rect 66376 29402 66400 29404
rect 66456 29402 66480 29404
rect 66536 29402 66560 29404
rect 66616 29402 66622 29404
rect 66376 29350 66378 29402
rect 66558 29350 66560 29402
rect 66314 29348 66320 29350
rect 66376 29348 66400 29350
rect 66456 29348 66480 29350
rect 66536 29348 66560 29350
rect 66616 29348 66622 29350
rect 66314 29339 66622 29348
rect 48504 29164 48556 29170
rect 48504 29106 48556 29112
rect 48320 28960 48372 28966
rect 48320 28902 48372 28908
rect 48228 28416 48280 28422
rect 48228 28358 48280 28364
rect 48332 28082 48360 28902
rect 48516 28218 48544 29106
rect 49240 28960 49292 28966
rect 49240 28902 49292 28908
rect 49252 28626 49280 28902
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 49240 28620 49292 28626
rect 49240 28562 49292 28568
rect 49516 28552 49568 28558
rect 49516 28494 49568 28500
rect 48504 28212 48556 28218
rect 48504 28154 48556 28160
rect 48320 28076 48372 28082
rect 48320 28018 48372 28024
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 46756 26308 46808 26314
rect 46756 26250 46808 26256
rect 46768 26042 46796 26250
rect 46756 26036 46808 26042
rect 46756 25978 46808 25984
rect 46768 25770 46796 25978
rect 47688 25838 47716 27814
rect 49332 27328 49384 27334
rect 49332 27270 49384 27276
rect 48412 27124 48464 27130
rect 48412 27066 48464 27072
rect 48424 26314 48452 27066
rect 48504 26920 48556 26926
rect 48504 26862 48556 26868
rect 49148 26920 49200 26926
rect 49148 26862 49200 26868
rect 48516 26450 48544 26862
rect 49160 26586 49188 26862
rect 49148 26580 49200 26586
rect 49148 26522 49200 26528
rect 48504 26444 48556 26450
rect 48504 26386 48556 26392
rect 49344 26382 49372 27270
rect 49528 26518 49556 28494
rect 55956 28416 56008 28422
rect 55956 28358 56008 28364
rect 51264 27328 51316 27334
rect 51264 27270 51316 27276
rect 51276 26926 51304 27270
rect 53932 27056 53984 27062
rect 53932 26998 53984 27004
rect 51172 26920 51224 26926
rect 51172 26862 51224 26868
rect 51264 26920 51316 26926
rect 51264 26862 51316 26868
rect 52368 26920 52420 26926
rect 52368 26862 52420 26868
rect 49976 26784 50028 26790
rect 49976 26726 50028 26732
rect 51080 26784 51132 26790
rect 51080 26726 51132 26732
rect 49516 26512 49568 26518
rect 49516 26454 49568 26460
rect 49988 26450 50016 26726
rect 51092 26518 51120 26726
rect 51080 26512 51132 26518
rect 51080 26454 51132 26460
rect 49976 26444 50028 26450
rect 49976 26386 50028 26392
rect 49332 26376 49384 26382
rect 49332 26318 49384 26324
rect 48412 26308 48464 26314
rect 48412 26250 48464 26256
rect 48504 26308 48556 26314
rect 48504 26250 48556 26256
rect 49884 26308 49936 26314
rect 49884 26250 49936 26256
rect 47676 25832 47728 25838
rect 47676 25774 47728 25780
rect 47952 25832 48004 25838
rect 47952 25774 48004 25780
rect 46756 25764 46808 25770
rect 46756 25706 46808 25712
rect 46572 25288 46624 25294
rect 46572 25230 46624 25236
rect 46388 24948 46440 24954
rect 46388 24890 46440 24896
rect 45468 24744 45520 24750
rect 45468 24686 45520 24692
rect 45480 24274 45508 24686
rect 45468 24268 45520 24274
rect 45468 24210 45520 24216
rect 45744 24132 45796 24138
rect 45744 24074 45796 24080
rect 45756 23866 45784 24074
rect 45834 24032 45890 24041
rect 45834 23967 45890 23976
rect 45744 23860 45796 23866
rect 45744 23802 45796 23808
rect 45848 23662 45876 23967
rect 46400 23730 46428 24890
rect 46388 23724 46440 23730
rect 46388 23666 46440 23672
rect 45836 23656 45888 23662
rect 45836 23598 45888 23604
rect 45376 23248 45428 23254
rect 45376 23190 45428 23196
rect 44732 23180 44784 23186
rect 44732 23122 44784 23128
rect 45192 23180 45244 23186
rect 45192 23122 45244 23128
rect 44560 23072 44680 23100
rect 44454 22400 44510 22409
rect 44454 22335 44510 22344
rect 44088 20528 44140 20534
rect 44364 20528 44416 20534
rect 44088 20470 44140 20476
rect 44284 20476 44364 20482
rect 44284 20470 44416 20476
rect 44100 19786 44128 20470
rect 44284 20454 44404 20470
rect 44180 20324 44232 20330
rect 44180 20266 44232 20272
rect 44088 19780 44140 19786
rect 44088 19722 44140 19728
rect 44192 19378 44220 20266
rect 44284 19718 44312 20454
rect 44364 20256 44416 20262
rect 44364 20198 44416 20204
rect 44376 20097 44404 20198
rect 44362 20088 44418 20097
rect 44362 20023 44418 20032
rect 44272 19712 44324 19718
rect 44272 19654 44324 19660
rect 44284 19514 44312 19654
rect 44272 19508 44324 19514
rect 44272 19450 44324 19456
rect 43720 19314 43772 19320
rect 43732 18766 43760 19314
rect 43916 19306 44036 19334
rect 44180 19372 44232 19378
rect 44180 19314 44232 19320
rect 43812 19168 43864 19174
rect 43812 19110 43864 19116
rect 43720 18760 43772 18766
rect 43720 18702 43772 18708
rect 43720 17536 43772 17542
rect 43720 17478 43772 17484
rect 43732 17202 43760 17478
rect 43720 17196 43772 17202
rect 43720 17138 43772 17144
rect 43628 16992 43680 16998
rect 43628 16934 43680 16940
rect 43352 15904 43404 15910
rect 43352 15846 43404 15852
rect 43364 15162 43392 15846
rect 43536 15496 43588 15502
rect 43536 15438 43588 15444
rect 43548 15366 43576 15438
rect 43444 15360 43496 15366
rect 43444 15302 43496 15308
rect 43536 15360 43588 15366
rect 43536 15302 43588 15308
rect 43720 15360 43772 15366
rect 43720 15302 43772 15308
rect 43456 15162 43484 15302
rect 43352 15156 43404 15162
rect 43352 15098 43404 15104
rect 43444 15156 43496 15162
rect 43444 15098 43496 15104
rect 43352 14544 43404 14550
rect 43352 14486 43404 14492
rect 43364 14396 43392 14486
rect 43548 14414 43576 15302
rect 43732 14958 43760 15302
rect 43720 14952 43772 14958
rect 43720 14894 43772 14900
rect 43628 14816 43680 14822
rect 43824 14793 43852 19110
rect 43628 14758 43680 14764
rect 43810 14784 43866 14793
rect 43640 14482 43668 14758
rect 43810 14719 43866 14728
rect 43916 14618 43944 19306
rect 44364 18352 44416 18358
rect 44364 18294 44416 18300
rect 44376 16590 44404 18294
rect 44364 16584 44416 16590
rect 44364 16526 44416 16532
rect 44272 16448 44324 16454
rect 44272 16390 44324 16396
rect 43996 15020 44048 15026
rect 43996 14962 44048 14968
rect 44008 14618 44036 14962
rect 44088 14816 44140 14822
rect 44088 14758 44140 14764
rect 43904 14612 43956 14618
rect 43904 14554 43956 14560
rect 43996 14612 44048 14618
rect 43996 14554 44048 14560
rect 43628 14476 43680 14482
rect 43628 14418 43680 14424
rect 43536 14408 43588 14414
rect 43364 14368 43536 14396
rect 43536 14350 43588 14356
rect 43640 12238 43668 14418
rect 44100 14006 44128 14758
rect 44088 14000 44140 14006
rect 44088 13942 44140 13948
rect 44180 13524 44232 13530
rect 44180 13466 44232 13472
rect 44192 12374 44220 13466
rect 44284 12918 44312 16390
rect 44468 16250 44496 22335
rect 44560 22094 44588 23072
rect 44744 23050 44772 23122
rect 45204 23050 45232 23122
rect 46400 23118 46428 23666
rect 45376 23112 45428 23118
rect 45374 23080 45376 23089
rect 46020 23112 46072 23118
rect 45428 23080 45430 23089
rect 44732 23044 44784 23050
rect 44732 22986 44784 22992
rect 45192 23044 45244 23050
rect 46020 23054 46072 23060
rect 46388 23112 46440 23118
rect 46388 23054 46440 23060
rect 47308 23112 47360 23118
rect 47308 23054 47360 23060
rect 45374 23015 45430 23024
rect 45192 22986 45244 22992
rect 44640 22976 44692 22982
rect 44640 22918 44692 22924
rect 45008 22976 45060 22982
rect 45100 22976 45152 22982
rect 45008 22918 45060 22924
rect 45098 22944 45100 22953
rect 45152 22944 45154 22953
rect 44652 22710 44680 22918
rect 44640 22704 44692 22710
rect 44640 22646 44692 22652
rect 45020 22642 45048 22918
rect 45098 22879 45154 22888
rect 45192 22772 45244 22778
rect 45192 22714 45244 22720
rect 45008 22636 45060 22642
rect 45008 22578 45060 22584
rect 44916 22432 44968 22438
rect 44916 22374 44968 22380
rect 44560 22066 44680 22094
rect 44548 20868 44600 20874
rect 44548 20810 44600 20816
rect 44560 19990 44588 20810
rect 44548 19984 44600 19990
rect 44548 19926 44600 19932
rect 44548 19780 44600 19786
rect 44548 19722 44600 19728
rect 44560 19378 44588 19722
rect 44548 19372 44600 19378
rect 44548 19314 44600 19320
rect 44652 19310 44680 22066
rect 44928 21486 44956 22374
rect 45204 22166 45232 22714
rect 45744 22636 45796 22642
rect 45744 22578 45796 22584
rect 45284 22228 45336 22234
rect 45284 22170 45336 22176
rect 45192 22160 45244 22166
rect 45192 22102 45244 22108
rect 45100 21956 45152 21962
rect 45100 21898 45152 21904
rect 45112 21554 45140 21898
rect 45100 21548 45152 21554
rect 45100 21490 45152 21496
rect 44916 21480 44968 21486
rect 44916 21422 44968 21428
rect 44732 20868 44784 20874
rect 44732 20810 44784 20816
rect 44744 19689 44772 20810
rect 44730 19680 44786 19689
rect 44730 19615 44786 19624
rect 44640 19304 44692 19310
rect 44640 19246 44692 19252
rect 44652 18698 44680 19246
rect 44640 18692 44692 18698
rect 44640 18634 44692 18640
rect 44548 18080 44600 18086
rect 44548 18022 44600 18028
rect 44560 17785 44588 18022
rect 44546 17776 44602 17785
rect 44546 17711 44548 17720
rect 44600 17711 44602 17720
rect 44548 17682 44600 17688
rect 44456 16244 44508 16250
rect 44456 16186 44508 16192
rect 44468 16153 44496 16186
rect 44454 16144 44510 16153
rect 44454 16079 44510 16088
rect 44364 14884 44416 14890
rect 44364 14826 44416 14832
rect 44376 14346 44404 14826
rect 44640 14476 44692 14482
rect 44640 14418 44692 14424
rect 44364 14340 44416 14346
rect 44364 14282 44416 14288
rect 44272 12912 44324 12918
rect 44272 12854 44324 12860
rect 44272 12708 44324 12714
rect 44272 12650 44324 12656
rect 44180 12368 44232 12374
rect 44180 12310 44232 12316
rect 43628 12232 43680 12238
rect 43628 12174 43680 12180
rect 43352 11144 43404 11150
rect 43352 11086 43404 11092
rect 43364 10674 43392 11086
rect 43640 10792 43668 12174
rect 44192 11354 44220 12310
rect 44284 12102 44312 12650
rect 44272 12096 44324 12102
rect 44272 12038 44324 12044
rect 44180 11348 44232 11354
rect 44180 11290 44232 11296
rect 44180 11144 44232 11150
rect 44180 11086 44232 11092
rect 44192 10810 44220 11086
rect 44272 11008 44324 11014
rect 44272 10950 44324 10956
rect 44180 10804 44232 10810
rect 43640 10764 43760 10792
rect 43732 10674 43760 10764
rect 44180 10746 44232 10752
rect 44284 10742 44312 10950
rect 44272 10736 44324 10742
rect 44272 10678 44324 10684
rect 43352 10668 43404 10674
rect 43352 10610 43404 10616
rect 43628 10668 43680 10674
rect 43628 10610 43680 10616
rect 43720 10668 43772 10674
rect 43720 10610 43772 10616
rect 43364 10266 43392 10610
rect 43352 10260 43404 10266
rect 43352 10202 43404 10208
rect 43536 10260 43588 10266
rect 43536 10202 43588 10208
rect 43352 10056 43404 10062
rect 43272 10016 43352 10044
rect 43352 9998 43404 10004
rect 43548 9586 43576 10202
rect 43260 9580 43312 9586
rect 43260 9522 43312 9528
rect 43536 9580 43588 9586
rect 43536 9522 43588 9528
rect 43272 9178 43300 9522
rect 43260 9172 43312 9178
rect 43260 9114 43312 9120
rect 43640 8945 43668 10610
rect 43996 10600 44048 10606
rect 43996 10542 44048 10548
rect 44008 10130 44036 10542
rect 44272 10464 44324 10470
rect 44272 10406 44324 10412
rect 43996 10124 44048 10130
rect 43996 10066 44048 10072
rect 43904 10056 43956 10062
rect 43904 9998 43956 10004
rect 43720 9376 43772 9382
rect 43720 9318 43772 9324
rect 43626 8936 43682 8945
rect 43626 8871 43682 8880
rect 43168 8628 43220 8634
rect 43168 8570 43220 8576
rect 43536 8628 43588 8634
rect 43536 8570 43588 8576
rect 43076 8084 43128 8090
rect 43076 8026 43128 8032
rect 43076 7200 43128 7206
rect 43076 7142 43128 7148
rect 43088 6390 43116 7142
rect 43076 6384 43128 6390
rect 43076 6326 43128 6332
rect 43076 5228 43128 5234
rect 42996 5188 43076 5216
rect 43076 5170 43128 5176
rect 43076 4548 43128 4554
rect 43076 4490 43128 4496
rect 42984 4480 43036 4486
rect 42984 4422 43036 4428
rect 42892 4140 42944 4146
rect 42892 4082 42944 4088
rect 42904 3670 42932 4082
rect 42996 3670 43024 4422
rect 43088 4282 43116 4490
rect 43076 4276 43128 4282
rect 43076 4218 43128 4224
rect 42892 3664 42944 3670
rect 42892 3606 42944 3612
rect 42984 3664 43036 3670
rect 42984 3606 43036 3612
rect 42800 3596 42852 3602
rect 42800 3538 42852 3544
rect 42996 3482 43024 3606
rect 42720 3466 43024 3482
rect 41420 3460 41472 3466
rect 41420 3402 41472 3408
rect 42708 3460 43024 3466
rect 42760 3454 43024 3460
rect 42708 3402 42760 3408
rect 41420 2848 41472 2854
rect 41420 2790 41472 2796
rect 40420 2746 40724 2774
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 40696 2514 40724 2746
rect 39488 2508 39540 2514
rect 39488 2450 39540 2456
rect 40684 2508 40736 2514
rect 40684 2450 40736 2456
rect 41432 2446 41460 2790
rect 43180 2774 43208 8570
rect 43352 8492 43404 8498
rect 43352 8434 43404 8440
rect 43364 8090 43392 8434
rect 43352 8084 43404 8090
rect 43352 8026 43404 8032
rect 43548 7970 43576 8570
rect 43732 8566 43760 9318
rect 43812 8832 43864 8838
rect 43812 8774 43864 8780
rect 43720 8560 43772 8566
rect 43720 8502 43772 8508
rect 43824 8498 43852 8774
rect 43812 8492 43864 8498
rect 43812 8434 43864 8440
rect 43720 8424 43772 8430
rect 43720 8366 43772 8372
rect 43732 8265 43760 8366
rect 43718 8256 43774 8265
rect 43718 8191 43774 8200
rect 43364 7942 43576 7970
rect 43364 7274 43392 7942
rect 43720 7404 43772 7410
rect 43720 7346 43772 7352
rect 43352 7268 43404 7274
rect 43352 7210 43404 7216
rect 43364 6866 43392 7210
rect 43732 7041 43760 7346
rect 43718 7032 43774 7041
rect 43718 6967 43774 6976
rect 43352 6860 43404 6866
rect 43352 6802 43404 6808
rect 43260 6724 43312 6730
rect 43260 6666 43312 6672
rect 43272 6458 43300 6666
rect 43260 6452 43312 6458
rect 43260 6394 43312 6400
rect 43364 6322 43392 6802
rect 43352 6316 43404 6322
rect 43352 6258 43404 6264
rect 43720 6112 43772 6118
rect 43720 6054 43772 6060
rect 43444 5024 43496 5030
rect 43444 4966 43496 4972
rect 43456 4146 43484 4966
rect 43628 4820 43680 4826
rect 43628 4762 43680 4768
rect 43444 4140 43496 4146
rect 43444 4082 43496 4088
rect 43260 3664 43312 3670
rect 43260 3606 43312 3612
rect 43088 2746 43208 2774
rect 43088 2446 43116 2746
rect 43168 2576 43220 2582
rect 43168 2518 43220 2524
rect 41420 2440 41472 2446
rect 41420 2382 41472 2388
rect 43076 2440 43128 2446
rect 43076 2382 43128 2388
rect 42524 2304 42576 2310
rect 42524 2246 42576 2252
rect 42536 800 42564 2246
rect 43180 800 43208 2518
rect 43272 2446 43300 3606
rect 43640 3466 43668 4762
rect 43732 4010 43760 6054
rect 43916 5234 43944 9998
rect 44284 9994 44312 10406
rect 44272 9988 44324 9994
rect 44272 9930 44324 9936
rect 44376 9674 44404 14282
rect 44652 13462 44680 14418
rect 44548 13456 44600 13462
rect 44548 13398 44600 13404
rect 44640 13456 44692 13462
rect 44640 13398 44692 13404
rect 44456 13320 44508 13326
rect 44456 13262 44508 13268
rect 44468 12782 44496 13262
rect 44560 12850 44588 13398
rect 44640 13184 44692 13190
rect 44640 13126 44692 13132
rect 44548 12844 44600 12850
rect 44548 12786 44600 12792
rect 44456 12776 44508 12782
rect 44456 12718 44508 12724
rect 44560 12442 44588 12786
rect 44548 12436 44600 12442
rect 44548 12378 44600 12384
rect 44284 9646 44404 9674
rect 44180 9036 44232 9042
rect 44180 8978 44232 8984
rect 44088 8968 44140 8974
rect 44086 8936 44088 8945
rect 44140 8936 44142 8945
rect 44086 8871 44142 8880
rect 44192 8498 44220 8978
rect 44180 8492 44232 8498
rect 44180 8434 44232 8440
rect 44192 8022 44220 8434
rect 44180 8016 44232 8022
rect 44180 7958 44232 7964
rect 44284 7002 44312 9646
rect 44364 8968 44416 8974
rect 44364 8910 44416 8916
rect 44456 8968 44508 8974
rect 44456 8910 44508 8916
rect 44272 6996 44324 7002
rect 44272 6938 44324 6944
rect 44284 6848 44312 6938
rect 44192 6820 44312 6848
rect 44192 6458 44220 6820
rect 44272 6724 44324 6730
rect 44272 6666 44324 6672
rect 44180 6452 44232 6458
rect 44180 6394 44232 6400
rect 44192 5370 44220 6394
rect 44180 5364 44232 5370
rect 44180 5306 44232 5312
rect 43904 5228 43956 5234
rect 43904 5170 43956 5176
rect 43720 4004 43772 4010
rect 43720 3946 43772 3952
rect 43916 3466 43944 5170
rect 44284 4690 44312 6666
rect 44376 5914 44404 8910
rect 44468 7546 44496 8910
rect 44652 8786 44680 13126
rect 44744 9081 44772 19615
rect 44824 19168 44876 19174
rect 44824 19110 44876 19116
rect 44836 11150 44864 19110
rect 44928 16250 44956 21422
rect 45204 20942 45232 22102
rect 45296 21554 45324 22170
rect 45756 21962 45784 22578
rect 45560 21956 45612 21962
rect 45560 21898 45612 21904
rect 45744 21956 45796 21962
rect 45744 21898 45796 21904
rect 45376 21616 45428 21622
rect 45376 21558 45428 21564
rect 45284 21548 45336 21554
rect 45284 21490 45336 21496
rect 45388 21010 45416 21558
rect 45572 21078 45600 21898
rect 45560 21072 45612 21078
rect 45560 21014 45612 21020
rect 45376 21004 45428 21010
rect 45376 20946 45428 20952
rect 45572 20942 45600 21014
rect 45192 20936 45244 20942
rect 45192 20878 45244 20884
rect 45560 20936 45612 20942
rect 45560 20878 45612 20884
rect 45192 20800 45244 20806
rect 45192 20742 45244 20748
rect 45204 20398 45232 20742
rect 46032 20534 46060 23054
rect 46400 22030 46428 23054
rect 46664 23044 46716 23050
rect 46664 22986 46716 22992
rect 46388 22024 46440 22030
rect 46388 21966 46440 21972
rect 46676 21622 46704 22986
rect 47216 22568 47268 22574
rect 47216 22510 47268 22516
rect 47228 22234 47256 22510
rect 47216 22228 47268 22234
rect 47216 22170 47268 22176
rect 46756 22160 46808 22166
rect 46754 22128 46756 22137
rect 46808 22128 46810 22137
rect 46754 22063 46810 22072
rect 47032 22024 47084 22030
rect 47032 21966 47084 21972
rect 46940 21888 46992 21894
rect 46940 21830 46992 21836
rect 46664 21616 46716 21622
rect 46664 21558 46716 21564
rect 46112 21412 46164 21418
rect 46112 21354 46164 21360
rect 46124 21146 46152 21354
rect 46204 21344 46256 21350
rect 46204 21286 46256 21292
rect 46112 21140 46164 21146
rect 46112 21082 46164 21088
rect 46020 20528 46072 20534
rect 46020 20470 46072 20476
rect 45192 20392 45244 20398
rect 45192 20334 45244 20340
rect 45204 19514 45232 20334
rect 46032 19990 46060 20470
rect 46020 19984 46072 19990
rect 46020 19926 46072 19932
rect 45192 19508 45244 19514
rect 45192 19450 45244 19456
rect 46216 19145 46244 21286
rect 46676 20466 46704 21558
rect 46952 21554 46980 21830
rect 46940 21548 46992 21554
rect 46940 21490 46992 21496
rect 46756 20936 46808 20942
rect 46756 20878 46808 20884
rect 46664 20460 46716 20466
rect 46664 20402 46716 20408
rect 46676 19854 46704 20402
rect 46664 19848 46716 19854
rect 46664 19790 46716 19796
rect 46202 19136 46258 19145
rect 46202 19071 46258 19080
rect 45192 18760 45244 18766
rect 45192 18702 45244 18708
rect 45008 17128 45060 17134
rect 45008 17070 45060 17076
rect 45020 16658 45048 17070
rect 45008 16652 45060 16658
rect 45008 16594 45060 16600
rect 44916 16244 44968 16250
rect 44916 16186 44968 16192
rect 45008 14816 45060 14822
rect 45008 14758 45060 14764
rect 44916 14544 44968 14550
rect 44916 14486 44968 14492
rect 44928 13326 44956 14486
rect 45020 14346 45048 14758
rect 45100 14476 45152 14482
rect 45100 14418 45152 14424
rect 45008 14340 45060 14346
rect 45008 14282 45060 14288
rect 45020 13530 45048 14282
rect 45112 13734 45140 14418
rect 45204 14385 45232 18702
rect 45560 18216 45612 18222
rect 45560 18158 45612 18164
rect 45572 17882 45600 18158
rect 45560 17876 45612 17882
rect 45560 17818 45612 17824
rect 46296 17808 46348 17814
rect 46296 17750 46348 17756
rect 46020 17672 46072 17678
rect 45926 17640 45982 17649
rect 46020 17614 46072 17620
rect 46112 17672 46164 17678
rect 46112 17614 46164 17620
rect 45926 17575 45928 17584
rect 45980 17575 45982 17584
rect 45928 17546 45980 17552
rect 45652 17332 45704 17338
rect 45652 17274 45704 17280
rect 45468 17196 45520 17202
rect 45468 17138 45520 17144
rect 45560 17196 45612 17202
rect 45560 17138 45612 17144
rect 45480 16726 45508 17138
rect 45572 16794 45600 17138
rect 45560 16788 45612 16794
rect 45560 16730 45612 16736
rect 45468 16720 45520 16726
rect 45664 16674 45692 17274
rect 45940 17270 45968 17546
rect 45928 17264 45980 17270
rect 45928 17206 45980 17212
rect 45744 17196 45796 17202
rect 45744 17138 45796 17144
rect 45468 16662 45520 16668
rect 45572 16646 45692 16674
rect 45756 16658 45784 17138
rect 45836 17060 45888 17066
rect 45836 17002 45888 17008
rect 45744 16652 45796 16658
rect 45468 16108 45520 16114
rect 45468 16050 45520 16056
rect 45480 15366 45508 16050
rect 45468 15360 45520 15366
rect 45468 15302 45520 15308
rect 45376 14952 45428 14958
rect 45480 14929 45508 15302
rect 45572 15026 45600 16646
rect 45744 16594 45796 16600
rect 45652 16244 45704 16250
rect 45652 16186 45704 16192
rect 45560 15020 45612 15026
rect 45560 14962 45612 14968
rect 45376 14894 45428 14900
rect 45466 14920 45522 14929
rect 45190 14376 45246 14385
rect 45190 14311 45192 14320
rect 45244 14311 45246 14320
rect 45192 14282 45244 14288
rect 45284 14272 45336 14278
rect 45284 14214 45336 14220
rect 45100 13728 45152 13734
rect 45100 13670 45152 13676
rect 45008 13524 45060 13530
rect 45008 13466 45060 13472
rect 44916 13320 44968 13326
rect 44916 13262 44968 13268
rect 44928 12714 44956 13262
rect 45112 12986 45140 13670
rect 45296 13326 45324 14214
rect 45388 13734 45416 14894
rect 45466 14855 45522 14864
rect 45376 13728 45428 13734
rect 45376 13670 45428 13676
rect 45284 13320 45336 13326
rect 45284 13262 45336 13268
rect 45100 12980 45152 12986
rect 45100 12922 45152 12928
rect 45112 12850 45140 12922
rect 45100 12844 45152 12850
rect 45100 12786 45152 12792
rect 44916 12708 44968 12714
rect 44916 12650 44968 12656
rect 45296 12434 45324 13262
rect 45388 13258 45416 13670
rect 45664 13433 45692 16186
rect 45756 16114 45784 16594
rect 45744 16108 45796 16114
rect 45744 16050 45796 16056
rect 45744 15564 45796 15570
rect 45744 15506 45796 15512
rect 45756 14482 45784 15506
rect 45848 15473 45876 17002
rect 45940 16046 45968 17206
rect 46032 17134 46060 17614
rect 46124 17338 46152 17614
rect 46204 17536 46256 17542
rect 46204 17478 46256 17484
rect 46112 17332 46164 17338
rect 46112 17274 46164 17280
rect 46216 17202 46244 17478
rect 46204 17196 46256 17202
rect 46204 17138 46256 17144
rect 46020 17128 46072 17134
rect 46020 17070 46072 17076
rect 46032 16794 46060 17070
rect 46020 16788 46072 16794
rect 46020 16730 46072 16736
rect 46112 16584 46164 16590
rect 46112 16526 46164 16532
rect 46020 16244 46072 16250
rect 46020 16186 46072 16192
rect 45928 16040 45980 16046
rect 45928 15982 45980 15988
rect 46032 15858 46060 16186
rect 46124 15910 46152 16526
rect 46216 16114 46244 17138
rect 46308 16998 46336 17750
rect 46296 16992 46348 16998
rect 46296 16934 46348 16940
rect 46308 16794 46336 16934
rect 46296 16788 46348 16794
rect 46296 16730 46348 16736
rect 46480 16584 46532 16590
rect 46480 16526 46532 16532
rect 46492 16250 46520 16526
rect 46480 16244 46532 16250
rect 46480 16186 46532 16192
rect 46204 16108 46256 16114
rect 46204 16050 46256 16056
rect 46768 15910 46796 20878
rect 46848 19984 46900 19990
rect 46848 19926 46900 19932
rect 46860 19446 46888 19926
rect 46952 19854 46980 21490
rect 47044 20602 47072 21966
rect 47124 21072 47176 21078
rect 47124 21014 47176 21020
rect 47136 20874 47164 21014
rect 47124 20868 47176 20874
rect 47124 20810 47176 20816
rect 47032 20596 47084 20602
rect 47032 20538 47084 20544
rect 46940 19848 46992 19854
rect 46940 19790 46992 19796
rect 47044 19718 47072 20538
rect 47032 19712 47084 19718
rect 47032 19654 47084 19660
rect 47136 19514 47164 20810
rect 47214 20632 47270 20641
rect 47214 20567 47270 20576
rect 47228 20534 47256 20567
rect 47216 20528 47268 20534
rect 47216 20470 47268 20476
rect 47320 20466 47348 23054
rect 47398 22672 47454 22681
rect 47398 22607 47454 22616
rect 47412 22234 47440 22607
rect 47400 22228 47452 22234
rect 47400 22170 47452 22176
rect 47412 22098 47440 22170
rect 47400 22092 47452 22098
rect 47400 22034 47452 22040
rect 47400 21344 47452 21350
rect 47400 21286 47452 21292
rect 47308 20460 47360 20466
rect 47308 20402 47360 20408
rect 47412 20398 47440 21286
rect 47400 20392 47452 20398
rect 47400 20334 47452 20340
rect 47412 20058 47440 20334
rect 47400 20052 47452 20058
rect 47400 19994 47452 20000
rect 47412 19786 47440 19994
rect 47216 19780 47268 19786
rect 47216 19722 47268 19728
rect 47400 19780 47452 19786
rect 47400 19722 47452 19728
rect 47124 19508 47176 19514
rect 47124 19450 47176 19456
rect 46848 19440 46900 19446
rect 46848 19382 46900 19388
rect 47136 19310 47164 19450
rect 47124 19304 47176 19310
rect 47124 19246 47176 19252
rect 47228 18902 47256 19722
rect 47216 18896 47268 18902
rect 47216 18838 47268 18844
rect 47308 18896 47360 18902
rect 47308 18838 47360 18844
rect 46848 18420 46900 18426
rect 46848 18362 46900 18368
rect 46860 16658 46888 18362
rect 47032 18080 47084 18086
rect 47032 18022 47084 18028
rect 47044 17746 47072 18022
rect 47320 17814 47348 18838
rect 47584 17876 47636 17882
rect 47584 17818 47636 17824
rect 47308 17808 47360 17814
rect 47308 17750 47360 17756
rect 47032 17740 47084 17746
rect 47032 17682 47084 17688
rect 47596 17542 47624 17818
rect 47584 17536 47636 17542
rect 47584 17478 47636 17484
rect 47688 16794 47716 25774
rect 47964 22574 47992 25774
rect 48424 24886 48452 26250
rect 48516 26042 48544 26250
rect 49896 26042 49924 26250
rect 48504 26036 48556 26042
rect 48504 25978 48556 25984
rect 49884 26036 49936 26042
rect 49884 25978 49936 25984
rect 49148 25900 49200 25906
rect 49148 25842 49200 25848
rect 49424 25900 49476 25906
rect 49424 25842 49476 25848
rect 48412 24880 48464 24886
rect 48464 24828 48820 24834
rect 48412 24822 48820 24828
rect 48424 24806 48820 24822
rect 48412 24744 48464 24750
rect 48412 24686 48464 24692
rect 48424 24410 48452 24686
rect 48412 24404 48464 24410
rect 48412 24346 48464 24352
rect 48504 24268 48556 24274
rect 48504 24210 48556 24216
rect 48412 24200 48464 24206
rect 48412 24142 48464 24148
rect 48424 23798 48452 24142
rect 48412 23792 48464 23798
rect 48412 23734 48464 23740
rect 48320 23724 48372 23730
rect 48320 23666 48372 23672
rect 48044 23520 48096 23526
rect 48044 23462 48096 23468
rect 48056 23186 48084 23462
rect 48332 23322 48360 23666
rect 48228 23316 48280 23322
rect 48228 23258 48280 23264
rect 48320 23316 48372 23322
rect 48320 23258 48372 23264
rect 48044 23180 48096 23186
rect 48044 23122 48096 23128
rect 48240 22778 48268 23258
rect 48228 22772 48280 22778
rect 48228 22714 48280 22720
rect 48136 22704 48188 22710
rect 48188 22652 48360 22658
rect 48136 22646 48360 22652
rect 48148 22642 48360 22646
rect 48148 22636 48372 22642
rect 48148 22630 48320 22636
rect 48320 22578 48372 22584
rect 47952 22568 48004 22574
rect 47952 22510 48004 22516
rect 48424 22522 48452 23734
rect 48516 23662 48544 24210
rect 48792 24138 48820 24806
rect 49160 24614 49188 25842
rect 49436 24818 49464 25842
rect 49424 24812 49476 24818
rect 49424 24754 49476 24760
rect 49148 24608 49200 24614
rect 49148 24550 49200 24556
rect 48780 24132 48832 24138
rect 48700 24092 48780 24120
rect 48596 24064 48648 24070
rect 48700 24018 48728 24092
rect 48780 24074 48832 24080
rect 48648 24012 48728 24018
rect 48596 24006 48728 24012
rect 48608 23990 48728 24006
rect 48504 23656 48556 23662
rect 48504 23598 48556 23604
rect 48596 23180 48648 23186
rect 48596 23122 48648 23128
rect 48608 22642 48636 23122
rect 48700 23118 48728 23990
rect 48964 23724 49016 23730
rect 48964 23666 49016 23672
rect 48688 23112 48740 23118
rect 48688 23054 48740 23060
rect 48596 22636 48648 22642
rect 48596 22578 48648 22584
rect 47768 21956 47820 21962
rect 47768 21898 47820 21904
rect 47780 21554 47808 21898
rect 47768 21548 47820 21554
rect 47768 21490 47820 21496
rect 47860 20256 47912 20262
rect 47860 20198 47912 20204
rect 47768 19848 47820 19854
rect 47768 19790 47820 19796
rect 47780 19378 47808 19790
rect 47768 19372 47820 19378
rect 47768 19314 47820 19320
rect 47872 17882 47900 20198
rect 47964 19446 47992 22510
rect 48424 22494 48544 22522
rect 48136 21888 48188 21894
rect 48136 21830 48188 21836
rect 48044 21344 48096 21350
rect 48148 21332 48176 21830
rect 48096 21304 48176 21332
rect 48044 21286 48096 21292
rect 48042 20632 48098 20641
rect 48042 20567 48098 20576
rect 47952 19440 48004 19446
rect 47952 19382 48004 19388
rect 48056 19009 48084 20567
rect 48148 19242 48176 21304
rect 48410 21040 48466 21049
rect 48410 20975 48412 20984
rect 48464 20975 48466 20984
rect 48412 20946 48464 20952
rect 48412 20392 48464 20398
rect 48412 20334 48464 20340
rect 48424 20058 48452 20334
rect 48412 20052 48464 20058
rect 48412 19994 48464 20000
rect 48516 19990 48544 22494
rect 48596 22432 48648 22438
rect 48596 22374 48648 22380
rect 48608 21010 48636 22374
rect 48596 21004 48648 21010
rect 48596 20946 48648 20952
rect 48608 20806 48636 20946
rect 48596 20800 48648 20806
rect 48596 20742 48648 20748
rect 48608 20505 48636 20742
rect 48700 20534 48728 23054
rect 48870 22536 48926 22545
rect 48870 22471 48926 22480
rect 48884 21962 48912 22471
rect 48872 21956 48924 21962
rect 48872 21898 48924 21904
rect 48872 20800 48924 20806
rect 48872 20742 48924 20748
rect 48688 20528 48740 20534
rect 48594 20496 48650 20505
rect 48688 20470 48740 20476
rect 48594 20431 48650 20440
rect 48504 19984 48556 19990
rect 48504 19926 48556 19932
rect 48596 19780 48648 19786
rect 48596 19722 48648 19728
rect 48504 19508 48556 19514
rect 48504 19450 48556 19456
rect 48228 19304 48280 19310
rect 48228 19246 48280 19252
rect 48136 19236 48188 19242
rect 48136 19178 48188 19184
rect 48042 19000 48098 19009
rect 48042 18935 48098 18944
rect 47860 17876 47912 17882
rect 47912 17836 47992 17864
rect 47860 17818 47912 17824
rect 47964 17746 47992 17836
rect 47952 17740 48004 17746
rect 47952 17682 48004 17688
rect 47768 17672 47820 17678
rect 47768 17614 47820 17620
rect 47860 17672 47912 17678
rect 47860 17614 47912 17620
rect 47780 17542 47808 17614
rect 47768 17536 47820 17542
rect 47768 17478 47820 17484
rect 47676 16788 47728 16794
rect 47676 16730 47728 16736
rect 46848 16652 46900 16658
rect 46848 16594 46900 16600
rect 45940 15830 46060 15858
rect 46112 15904 46164 15910
rect 46112 15846 46164 15852
rect 46756 15904 46808 15910
rect 46756 15846 46808 15852
rect 45940 15706 45968 15830
rect 46768 15706 46796 15846
rect 45928 15700 45980 15706
rect 45928 15642 45980 15648
rect 46756 15700 46808 15706
rect 46756 15642 46808 15648
rect 45834 15464 45890 15473
rect 45834 15399 45836 15408
rect 45888 15399 45890 15408
rect 45836 15370 45888 15376
rect 45744 14476 45796 14482
rect 45744 14418 45796 14424
rect 45940 14362 45968 15642
rect 46860 15570 46888 16594
rect 47400 16516 47452 16522
rect 47400 16458 47452 16464
rect 47308 16448 47360 16454
rect 47308 16390 47360 16396
rect 46848 15564 46900 15570
rect 46848 15506 46900 15512
rect 46664 15020 46716 15026
rect 46664 14962 46716 14968
rect 45756 14334 45968 14362
rect 46020 14340 46072 14346
rect 45756 14074 45784 14334
rect 46020 14282 46072 14288
rect 46032 14074 46060 14282
rect 46676 14249 46704 14962
rect 46756 14476 46808 14482
rect 46756 14418 46808 14424
rect 46662 14240 46718 14249
rect 46662 14175 46718 14184
rect 46768 14074 46796 14418
rect 45744 14068 45796 14074
rect 45744 14010 45796 14016
rect 46020 14068 46072 14074
rect 46020 14010 46072 14016
rect 46756 14068 46808 14074
rect 46756 14010 46808 14016
rect 45650 13424 45706 13433
rect 45650 13359 45706 13368
rect 45376 13252 45428 13258
rect 45376 13194 45428 13200
rect 45560 13184 45612 13190
rect 45560 13126 45612 13132
rect 45376 12776 45428 12782
rect 45376 12718 45428 12724
rect 45388 12442 45416 12718
rect 45204 12406 45324 12434
rect 45376 12436 45428 12442
rect 44824 11144 44876 11150
rect 44824 11086 44876 11092
rect 45204 9994 45232 12406
rect 45376 12378 45428 12384
rect 45572 12238 45600 13126
rect 45560 12232 45612 12238
rect 45560 12174 45612 12180
rect 45664 11354 45692 13359
rect 45652 11348 45704 11354
rect 45652 11290 45704 11296
rect 45652 11076 45704 11082
rect 45652 11018 45704 11024
rect 45664 10810 45692 11018
rect 45756 11014 45784 14010
rect 46768 12918 46796 14010
rect 46860 13870 46888 15506
rect 47124 14816 47176 14822
rect 47124 14758 47176 14764
rect 46940 14068 46992 14074
rect 46940 14010 46992 14016
rect 46952 13938 46980 14010
rect 46940 13932 46992 13938
rect 46940 13874 46992 13880
rect 46848 13864 46900 13870
rect 46848 13806 46900 13812
rect 47136 13802 47164 14758
rect 47320 14414 47348 16390
rect 47412 16250 47440 16458
rect 47400 16244 47452 16250
rect 47400 16186 47452 16192
rect 47492 15360 47544 15366
rect 47492 15302 47544 15308
rect 47504 14618 47532 15302
rect 47492 14612 47544 14618
rect 47492 14554 47544 14560
rect 47308 14408 47360 14414
rect 47308 14350 47360 14356
rect 47504 14278 47532 14554
rect 47780 14550 47808 17478
rect 47872 16658 47900 17614
rect 48056 17202 48084 18935
rect 48148 18630 48176 19178
rect 48240 18970 48268 19246
rect 48228 18964 48280 18970
rect 48228 18906 48280 18912
rect 48136 18624 48188 18630
rect 48136 18566 48188 18572
rect 48136 17672 48188 17678
rect 48240 17660 48268 18906
rect 48412 18760 48464 18766
rect 48412 18702 48464 18708
rect 48320 18624 48372 18630
rect 48320 18566 48372 18572
rect 48332 18358 48360 18566
rect 48320 18352 48372 18358
rect 48320 18294 48372 18300
rect 48320 18216 48372 18222
rect 48320 18158 48372 18164
rect 48188 17632 48268 17660
rect 48136 17614 48188 17620
rect 48044 17196 48096 17202
rect 48044 17138 48096 17144
rect 47860 16652 47912 16658
rect 47860 16594 47912 16600
rect 47872 16182 47900 16594
rect 48228 16584 48280 16590
rect 48332 16572 48360 18158
rect 48424 17882 48452 18702
rect 48412 17876 48464 17882
rect 48412 17818 48464 17824
rect 48280 16544 48360 16572
rect 48228 16526 48280 16532
rect 48412 16448 48464 16454
rect 48412 16390 48464 16396
rect 48424 16182 48452 16390
rect 47860 16176 47912 16182
rect 47860 16118 47912 16124
rect 48412 16176 48464 16182
rect 48412 16118 48464 16124
rect 48516 16114 48544 19450
rect 48608 16114 48636 19722
rect 48700 19446 48728 20470
rect 48884 19854 48912 20742
rect 48976 20262 49004 23666
rect 49056 23588 49108 23594
rect 49056 23530 49108 23536
rect 49068 23254 49096 23530
rect 49056 23248 49108 23254
rect 49056 23190 49108 23196
rect 49068 22094 49096 23190
rect 49160 23186 49188 24550
rect 49436 24410 49464 24754
rect 49516 24608 49568 24614
rect 49516 24550 49568 24556
rect 49424 24404 49476 24410
rect 49424 24346 49476 24352
rect 49436 24206 49464 24346
rect 49528 24274 49556 24550
rect 49516 24268 49568 24274
rect 49516 24210 49568 24216
rect 49240 24200 49292 24206
rect 49424 24200 49476 24206
rect 49292 24148 49372 24154
rect 49240 24142 49372 24148
rect 49608 24200 49660 24206
rect 49424 24142 49476 24148
rect 49528 24148 49608 24154
rect 49528 24142 49660 24148
rect 49252 24126 49372 24142
rect 49344 23866 49372 24126
rect 49528 24126 49648 24142
rect 49884 24132 49936 24138
rect 49528 24018 49556 24126
rect 49988 24120 50016 26386
rect 51184 26364 51212 26862
rect 51092 26336 51212 26364
rect 50804 26308 50856 26314
rect 50804 26250 50856 26256
rect 50528 25696 50580 25702
rect 50528 25638 50580 25644
rect 50068 24200 50120 24206
rect 50068 24142 50120 24148
rect 49936 24092 50016 24120
rect 49884 24074 49936 24080
rect 49436 23990 49556 24018
rect 49332 23860 49384 23866
rect 49332 23802 49384 23808
rect 49240 23656 49292 23662
rect 49240 23598 49292 23604
rect 49148 23180 49200 23186
rect 49148 23122 49200 23128
rect 49252 22982 49280 23598
rect 49344 23118 49372 23802
rect 49436 23662 49464 23990
rect 49424 23656 49476 23662
rect 49424 23598 49476 23604
rect 49332 23112 49384 23118
rect 49332 23054 49384 23060
rect 49884 23044 49936 23050
rect 49884 22986 49936 22992
rect 49240 22976 49292 22982
rect 49700 22976 49752 22982
rect 49240 22918 49292 22924
rect 49698 22944 49700 22953
rect 49752 22944 49754 22953
rect 49068 22066 49188 22094
rect 48964 20256 49016 20262
rect 48964 20198 49016 20204
rect 49160 20058 49188 22066
rect 49252 22030 49280 22918
rect 49698 22879 49754 22888
rect 49700 22636 49752 22642
rect 49700 22578 49752 22584
rect 49792 22636 49844 22642
rect 49792 22578 49844 22584
rect 49516 22568 49568 22574
rect 49516 22510 49568 22516
rect 49528 22438 49556 22510
rect 49516 22432 49568 22438
rect 49516 22374 49568 22380
rect 49240 22024 49292 22030
rect 49240 21966 49292 21972
rect 49332 21956 49384 21962
rect 49332 21898 49384 21904
rect 49148 20052 49200 20058
rect 49148 19994 49200 20000
rect 48780 19848 48832 19854
rect 48780 19790 48832 19796
rect 48872 19848 48924 19854
rect 48872 19790 48924 19796
rect 49056 19848 49108 19854
rect 49056 19790 49108 19796
rect 48688 19440 48740 19446
rect 48688 19382 48740 19388
rect 48792 17814 48820 19790
rect 48872 19236 48924 19242
rect 48872 19178 48924 19184
rect 48780 17808 48832 17814
rect 48780 17750 48832 17756
rect 48884 16998 48912 19178
rect 49068 18193 49096 19790
rect 49160 19378 49188 19994
rect 49148 19372 49200 19378
rect 49148 19314 49200 19320
rect 49160 18902 49188 19314
rect 49148 18896 49200 18902
rect 49148 18838 49200 18844
rect 49054 18184 49110 18193
rect 49054 18119 49110 18128
rect 49056 17196 49108 17202
rect 49056 17138 49108 17144
rect 48872 16992 48924 16998
rect 48872 16934 48924 16940
rect 48884 16590 48912 16934
rect 48872 16584 48924 16590
rect 48872 16526 48924 16532
rect 48688 16448 48740 16454
rect 48688 16390 48740 16396
rect 48504 16108 48556 16114
rect 48504 16050 48556 16056
rect 48596 16108 48648 16114
rect 48596 16050 48648 16056
rect 48136 15496 48188 15502
rect 48136 15438 48188 15444
rect 48148 15162 48176 15438
rect 48608 15366 48636 16050
rect 48700 15910 48728 16390
rect 48688 15904 48740 15910
rect 48688 15846 48740 15852
rect 48596 15360 48648 15366
rect 48596 15302 48648 15308
rect 48136 15156 48188 15162
rect 48136 15098 48188 15104
rect 48228 15156 48280 15162
rect 48228 15098 48280 15104
rect 48148 15026 48176 15098
rect 48044 15020 48096 15026
rect 48044 14962 48096 14968
rect 48136 15020 48188 15026
rect 48136 14962 48188 14968
rect 47952 14952 48004 14958
rect 47952 14894 48004 14900
rect 47860 14816 47912 14822
rect 47860 14758 47912 14764
rect 47768 14544 47820 14550
rect 47768 14486 47820 14492
rect 47584 14408 47636 14414
rect 47636 14368 47716 14396
rect 47584 14350 47636 14356
rect 47492 14272 47544 14278
rect 47492 14214 47544 14220
rect 47504 14074 47532 14214
rect 47688 14074 47716 14368
rect 47492 14068 47544 14074
rect 47492 14010 47544 14016
rect 47676 14068 47728 14074
rect 47676 14010 47728 14016
rect 47872 14006 47900 14758
rect 47964 14346 47992 14894
rect 48056 14396 48084 14962
rect 48136 14408 48188 14414
rect 48056 14368 48136 14396
rect 47952 14340 48004 14346
rect 47952 14282 48004 14288
rect 47860 14000 47912 14006
rect 47860 13942 47912 13948
rect 47124 13796 47176 13802
rect 47124 13738 47176 13744
rect 47768 13796 47820 13802
rect 47768 13738 47820 13744
rect 46940 13728 46992 13734
rect 46940 13670 46992 13676
rect 46756 12912 46808 12918
rect 46756 12854 46808 12860
rect 46848 12640 46900 12646
rect 46848 12582 46900 12588
rect 46860 12306 46888 12582
rect 46952 12442 46980 13670
rect 47780 13326 47808 13738
rect 48056 13394 48084 14368
rect 48240 14385 48268 15098
rect 48780 14816 48832 14822
rect 48780 14758 48832 14764
rect 48792 14414 48820 14758
rect 48780 14408 48832 14414
rect 48136 14350 48188 14356
rect 48226 14376 48282 14385
rect 48780 14350 48832 14356
rect 48226 14311 48282 14320
rect 48412 14272 48464 14278
rect 48412 14214 48464 14220
rect 48424 14006 48452 14214
rect 48412 14000 48464 14006
rect 48412 13942 48464 13948
rect 48044 13388 48096 13394
rect 48044 13330 48096 13336
rect 47768 13320 47820 13326
rect 47768 13262 47820 13268
rect 46940 12436 46992 12442
rect 47780 12434 47808 13262
rect 47780 12406 47900 12434
rect 46940 12378 46992 12384
rect 46848 12300 46900 12306
rect 46848 12242 46900 12248
rect 45836 11824 45888 11830
rect 45836 11766 45888 11772
rect 45744 11008 45796 11014
rect 45744 10950 45796 10956
rect 45652 10804 45704 10810
rect 45652 10746 45704 10752
rect 45284 10532 45336 10538
rect 45284 10474 45336 10480
rect 45192 9988 45244 9994
rect 45192 9930 45244 9936
rect 45296 9722 45324 10474
rect 45560 9988 45612 9994
rect 45560 9930 45612 9936
rect 45572 9722 45600 9930
rect 45284 9716 45336 9722
rect 45284 9658 45336 9664
rect 45560 9716 45612 9722
rect 45560 9658 45612 9664
rect 44730 9072 44786 9081
rect 44730 9007 44786 9016
rect 44560 8758 44680 8786
rect 44456 7540 44508 7546
rect 44456 7482 44508 7488
rect 44456 6452 44508 6458
rect 44456 6394 44508 6400
rect 44468 6322 44496 6394
rect 44456 6316 44508 6322
rect 44456 6258 44508 6264
rect 44364 5908 44416 5914
rect 44364 5850 44416 5856
rect 44560 5302 44588 8758
rect 44744 8616 44772 9007
rect 45468 8968 45520 8974
rect 45468 8910 45520 8916
rect 44916 8900 44968 8906
rect 44916 8842 44968 8848
rect 44652 8588 44772 8616
rect 44652 7410 44680 8588
rect 44928 8498 44956 8842
rect 45480 8634 45508 8910
rect 45468 8628 45520 8634
rect 45468 8570 45520 8576
rect 45376 8560 45428 8566
rect 45376 8502 45428 8508
rect 44732 8492 44784 8498
rect 44732 8434 44784 8440
rect 44916 8492 44968 8498
rect 44916 8434 44968 8440
rect 45100 8492 45152 8498
rect 45100 8434 45152 8440
rect 44640 7404 44692 7410
rect 44640 7346 44692 7352
rect 44640 6928 44692 6934
rect 44640 6870 44692 6876
rect 44652 6322 44680 6870
rect 44640 6316 44692 6322
rect 44640 6258 44692 6264
rect 44548 5296 44600 5302
rect 44548 5238 44600 5244
rect 44272 4684 44324 4690
rect 44272 4626 44324 4632
rect 44284 3670 44312 4626
rect 44560 3670 44588 5238
rect 44744 4826 44772 8434
rect 44928 8401 44956 8434
rect 44914 8392 44970 8401
rect 44914 8327 44970 8336
rect 45112 8090 45140 8434
rect 45284 8288 45336 8294
rect 45282 8256 45284 8265
rect 45336 8256 45338 8265
rect 45282 8191 45338 8200
rect 45100 8084 45152 8090
rect 45100 8026 45152 8032
rect 45388 7886 45416 8502
rect 45652 8424 45704 8430
rect 45652 8366 45704 8372
rect 45664 7886 45692 8366
rect 45376 7880 45428 7886
rect 45376 7822 45428 7828
rect 45652 7880 45704 7886
rect 45652 7822 45704 7828
rect 45744 7880 45796 7886
rect 45744 7822 45796 7828
rect 44824 7200 44876 7206
rect 44824 7142 44876 7148
rect 44836 6390 44864 7142
rect 45664 6934 45692 7822
rect 45756 7274 45784 7822
rect 45848 7818 45876 11766
rect 46572 11620 46624 11626
rect 46572 11562 46624 11568
rect 46296 11348 46348 11354
rect 46296 11290 46348 11296
rect 46112 11008 46164 11014
rect 46112 10950 46164 10956
rect 46124 10674 46152 10950
rect 46308 10742 46336 11290
rect 46584 11150 46612 11562
rect 46952 11558 46980 12378
rect 47124 12232 47176 12238
rect 47124 12174 47176 12180
rect 46940 11552 46992 11558
rect 46940 11494 46992 11500
rect 46572 11144 46624 11150
rect 46572 11086 46624 11092
rect 46296 10736 46348 10742
rect 46296 10678 46348 10684
rect 46112 10668 46164 10674
rect 46112 10610 46164 10616
rect 46124 9722 46152 10610
rect 46112 9716 46164 9722
rect 46112 9658 46164 9664
rect 45928 9580 45980 9586
rect 45928 9522 45980 9528
rect 45940 8090 45968 9522
rect 46308 9110 46336 10678
rect 46584 10674 46612 11086
rect 46664 10736 46716 10742
rect 46664 10678 46716 10684
rect 46572 10668 46624 10674
rect 46572 10610 46624 10616
rect 46676 10554 46704 10678
rect 47136 10674 47164 12174
rect 47676 12164 47728 12170
rect 47676 12106 47728 12112
rect 47688 11898 47716 12106
rect 47676 11892 47728 11898
rect 47676 11834 47728 11840
rect 47872 11762 47900 12406
rect 48320 12096 48372 12102
rect 48320 12038 48372 12044
rect 47952 11892 48004 11898
rect 47952 11834 48004 11840
rect 47964 11762 47992 11834
rect 47860 11756 47912 11762
rect 47860 11698 47912 11704
rect 47952 11756 48004 11762
rect 47952 11698 48004 11704
rect 47872 11218 47900 11698
rect 48332 11694 48360 12038
rect 48792 11914 48820 14350
rect 48884 12434 48912 16526
rect 49068 16522 49096 17138
rect 49344 16590 49372 21898
rect 49528 20262 49556 22374
rect 49712 22234 49740 22578
rect 49804 22506 49832 22578
rect 49792 22500 49844 22506
rect 49792 22442 49844 22448
rect 49700 22228 49752 22234
rect 49700 22170 49752 22176
rect 49700 22092 49752 22098
rect 49700 22034 49752 22040
rect 49792 22092 49844 22098
rect 49792 22034 49844 22040
rect 49608 22024 49660 22030
rect 49608 21966 49660 21972
rect 49516 20256 49568 20262
rect 49516 20198 49568 20204
rect 49528 19854 49556 20198
rect 49516 19848 49568 19854
rect 49516 19790 49568 19796
rect 49516 17740 49568 17746
rect 49516 17682 49568 17688
rect 49332 16584 49384 16590
rect 49332 16526 49384 16532
rect 48964 16516 49016 16522
rect 48964 16458 49016 16464
rect 49056 16516 49108 16522
rect 49056 16458 49108 16464
rect 48976 15434 49004 16458
rect 49068 16046 49096 16458
rect 49056 16040 49108 16046
rect 49056 15982 49108 15988
rect 49344 15910 49372 16526
rect 49528 16153 49556 17682
rect 49514 16144 49570 16153
rect 49514 16079 49516 16088
rect 49568 16079 49570 16088
rect 49516 16050 49568 16056
rect 49424 16040 49476 16046
rect 49424 15982 49476 15988
rect 49332 15904 49384 15910
rect 49332 15846 49384 15852
rect 48964 15428 49016 15434
rect 48964 15370 49016 15376
rect 49240 13932 49292 13938
rect 49240 13874 49292 13880
rect 48884 12406 49096 12434
rect 48792 11886 49004 11914
rect 48504 11756 48556 11762
rect 48504 11698 48556 11704
rect 48596 11756 48648 11762
rect 48596 11698 48648 11704
rect 48872 11756 48924 11762
rect 48872 11698 48924 11704
rect 48320 11688 48372 11694
rect 48320 11630 48372 11636
rect 48136 11552 48188 11558
rect 48136 11494 48188 11500
rect 47860 11212 47912 11218
rect 47860 11154 47912 11160
rect 47124 10668 47176 10674
rect 47124 10610 47176 10616
rect 46584 10526 46704 10554
rect 47032 10600 47084 10606
rect 47032 10542 47084 10548
rect 46584 9994 46612 10526
rect 47044 10130 47072 10542
rect 47872 10130 47900 11154
rect 47952 10600 48004 10606
rect 47952 10542 48004 10548
rect 47964 10266 47992 10542
rect 48148 10266 48176 11494
rect 48332 11354 48360 11630
rect 48320 11348 48372 11354
rect 48320 11290 48372 11296
rect 48228 10464 48280 10470
rect 48228 10406 48280 10412
rect 47952 10260 48004 10266
rect 47952 10202 48004 10208
rect 48136 10260 48188 10266
rect 48136 10202 48188 10208
rect 46940 10124 46992 10130
rect 46940 10066 46992 10072
rect 47032 10124 47084 10130
rect 47032 10066 47084 10072
rect 47216 10124 47268 10130
rect 47216 10066 47268 10072
rect 47860 10124 47912 10130
rect 47860 10066 47912 10072
rect 46572 9988 46624 9994
rect 46572 9930 46624 9936
rect 46296 9104 46348 9110
rect 46296 9046 46348 9052
rect 46584 8566 46612 9930
rect 46848 9376 46900 9382
rect 46848 9318 46900 9324
rect 46860 8838 46888 9318
rect 46848 8832 46900 8838
rect 46848 8774 46900 8780
rect 46572 8560 46624 8566
rect 46572 8502 46624 8508
rect 45928 8084 45980 8090
rect 45928 8026 45980 8032
rect 45836 7812 45888 7818
rect 45836 7754 45888 7760
rect 45744 7268 45796 7274
rect 45744 7210 45796 7216
rect 45652 6928 45704 6934
rect 45006 6896 45062 6905
rect 45652 6870 45704 6876
rect 45006 6831 45008 6840
rect 45060 6831 45062 6840
rect 45008 6802 45060 6808
rect 44916 6656 44968 6662
rect 44916 6598 44968 6604
rect 44928 6458 44956 6598
rect 45020 6458 45048 6802
rect 45756 6730 45784 7210
rect 45848 6866 45876 7754
rect 46480 7540 46532 7546
rect 46480 7482 46532 7488
rect 46204 6996 46256 7002
rect 46204 6938 46256 6944
rect 46296 6996 46348 7002
rect 46296 6938 46348 6944
rect 45836 6860 45888 6866
rect 45836 6802 45888 6808
rect 45560 6724 45612 6730
rect 45560 6666 45612 6672
rect 45744 6724 45796 6730
rect 45744 6666 45796 6672
rect 44916 6452 44968 6458
rect 44916 6394 44968 6400
rect 45008 6452 45060 6458
rect 45008 6394 45060 6400
rect 44824 6384 44876 6390
rect 44824 6326 44876 6332
rect 44836 4826 44864 6326
rect 45572 6322 45600 6666
rect 45848 6662 45876 6802
rect 46216 6798 46244 6938
rect 46204 6792 46256 6798
rect 46204 6734 46256 6740
rect 45836 6656 45888 6662
rect 45836 6598 45888 6604
rect 45560 6316 45612 6322
rect 45560 6258 45612 6264
rect 45100 6248 45152 6254
rect 45020 6208 45100 6236
rect 44732 4820 44784 4826
rect 44732 4762 44784 4768
rect 44824 4820 44876 4826
rect 44824 4762 44876 4768
rect 44744 4486 44772 4762
rect 44836 4622 44864 4762
rect 44824 4616 44876 4622
rect 44824 4558 44876 4564
rect 44732 4480 44784 4486
rect 44732 4422 44784 4428
rect 44744 4146 44772 4422
rect 44732 4140 44784 4146
rect 44732 4082 44784 4088
rect 44272 3664 44324 3670
rect 44272 3606 44324 3612
rect 44548 3664 44600 3670
rect 44548 3606 44600 3612
rect 43628 3460 43680 3466
rect 43628 3402 43680 3408
rect 43904 3460 43956 3466
rect 43904 3402 43956 3408
rect 44284 3194 44312 3606
rect 44560 3466 44588 3606
rect 45020 3602 45048 6208
rect 45100 6190 45152 6196
rect 45572 4622 45600 6258
rect 45652 5160 45704 5166
rect 45652 5102 45704 5108
rect 45560 4616 45612 4622
rect 45560 4558 45612 4564
rect 45664 4486 45692 5102
rect 45848 4690 45876 6598
rect 46112 6248 46164 6254
rect 46112 6190 46164 6196
rect 46124 5914 46152 6190
rect 46112 5908 46164 5914
rect 46112 5850 46164 5856
rect 45836 4684 45888 4690
rect 45836 4626 45888 4632
rect 46124 4622 46152 5850
rect 46216 5574 46244 6734
rect 46308 6118 46336 6938
rect 46492 6798 46520 7482
rect 46480 6792 46532 6798
rect 46480 6734 46532 6740
rect 46584 6390 46612 8502
rect 46860 7954 46888 8774
rect 46952 8294 46980 10066
rect 47124 9920 47176 9926
rect 47124 9862 47176 9868
rect 47136 9586 47164 9862
rect 47124 9580 47176 9586
rect 47124 9522 47176 9528
rect 47228 9518 47256 10066
rect 47676 10056 47728 10062
rect 47676 9998 47728 10004
rect 47216 9512 47268 9518
rect 47216 9454 47268 9460
rect 47228 8566 47256 9454
rect 47216 8560 47268 8566
rect 47216 8502 47268 8508
rect 47124 8424 47176 8430
rect 47124 8366 47176 8372
rect 46940 8288 46992 8294
rect 46940 8230 46992 8236
rect 47136 8090 47164 8366
rect 47124 8084 47176 8090
rect 47124 8026 47176 8032
rect 46848 7948 46900 7954
rect 46848 7890 46900 7896
rect 46860 7002 46888 7890
rect 47124 7880 47176 7886
rect 47228 7868 47256 8502
rect 47688 7886 47716 9998
rect 48044 8424 48096 8430
rect 48044 8366 48096 8372
rect 48056 7954 48084 8366
rect 48044 7948 48096 7954
rect 48044 7890 48096 7896
rect 47176 7840 47256 7868
rect 47676 7880 47728 7886
rect 47124 7822 47176 7828
rect 47676 7822 47728 7828
rect 46848 6996 46900 7002
rect 46848 6938 46900 6944
rect 46664 6860 46716 6866
rect 46664 6802 46716 6808
rect 46676 6730 46704 6802
rect 46664 6724 46716 6730
rect 46664 6666 46716 6672
rect 46756 6724 46808 6730
rect 46756 6666 46808 6672
rect 46572 6384 46624 6390
rect 46572 6326 46624 6332
rect 46296 6112 46348 6118
rect 46296 6054 46348 6060
rect 46480 6112 46532 6118
rect 46480 6054 46532 6060
rect 46204 5568 46256 5574
rect 46204 5510 46256 5516
rect 46308 5030 46336 6054
rect 46492 5778 46520 6054
rect 46480 5772 46532 5778
rect 46480 5714 46532 5720
rect 46584 5642 46612 6326
rect 46768 6254 46796 6666
rect 46756 6248 46808 6254
rect 46756 6190 46808 6196
rect 46756 6112 46808 6118
rect 46756 6054 46808 6060
rect 46768 5778 46796 6054
rect 46756 5772 46808 5778
rect 46756 5714 46808 5720
rect 46572 5636 46624 5642
rect 46572 5578 46624 5584
rect 46296 5024 46348 5030
rect 46296 4966 46348 4972
rect 46112 4616 46164 4622
rect 46112 4558 46164 4564
rect 45560 4480 45612 4486
rect 45560 4422 45612 4428
rect 45652 4480 45704 4486
rect 45652 4422 45704 4428
rect 45572 4146 45600 4422
rect 45664 4146 45692 4422
rect 45560 4140 45612 4146
rect 45560 4082 45612 4088
rect 45652 4140 45704 4146
rect 45652 4082 45704 4088
rect 46308 4010 46336 4966
rect 46848 4684 46900 4690
rect 46848 4626 46900 4632
rect 46860 4554 46888 4626
rect 46848 4548 46900 4554
rect 46848 4490 46900 4496
rect 46756 4480 46808 4486
rect 46756 4422 46808 4428
rect 46296 4004 46348 4010
rect 46296 3946 46348 3952
rect 45284 3936 45336 3942
rect 45284 3878 45336 3884
rect 45296 3602 45324 3878
rect 46768 3738 46796 4422
rect 47136 4078 47164 7822
rect 47688 7546 47716 7822
rect 47676 7540 47728 7546
rect 47676 7482 47728 7488
rect 47308 6792 47360 6798
rect 47308 6734 47360 6740
rect 47320 6458 47348 6734
rect 47308 6452 47360 6458
rect 47308 6394 47360 6400
rect 47768 6384 47820 6390
rect 47768 6326 47820 6332
rect 47400 5024 47452 5030
rect 47400 4966 47452 4972
rect 47412 4826 47440 4966
rect 47400 4820 47452 4826
rect 47400 4762 47452 4768
rect 47308 4616 47360 4622
rect 47308 4558 47360 4564
rect 47676 4616 47728 4622
rect 47676 4558 47728 4564
rect 47320 4282 47348 4558
rect 47308 4276 47360 4282
rect 47308 4218 47360 4224
rect 47688 4078 47716 4558
rect 47780 4214 47808 6326
rect 48056 6254 48084 7890
rect 48240 7818 48268 10406
rect 48332 9994 48360 11290
rect 48516 11218 48544 11698
rect 48504 11212 48556 11218
rect 48504 11154 48556 11160
rect 48516 10044 48544 11154
rect 48608 11150 48636 11698
rect 48596 11144 48648 11150
rect 48594 11112 48596 11121
rect 48648 11112 48650 11121
rect 48594 11047 48650 11056
rect 48780 11076 48832 11082
rect 48780 11018 48832 11024
rect 48688 10260 48740 10266
rect 48688 10202 48740 10208
rect 48596 10056 48648 10062
rect 48516 10016 48596 10044
rect 48596 9998 48648 10004
rect 48320 9988 48372 9994
rect 48320 9930 48372 9936
rect 48700 9654 48728 10202
rect 48688 9648 48740 9654
rect 48688 9590 48740 9596
rect 48792 8634 48820 11018
rect 48884 10810 48912 11698
rect 48872 10804 48924 10810
rect 48872 10746 48924 10752
rect 48872 10192 48924 10198
rect 48872 10134 48924 10140
rect 48884 10062 48912 10134
rect 48872 10056 48924 10062
rect 48872 9998 48924 10004
rect 48872 9376 48924 9382
rect 48872 9318 48924 9324
rect 48780 8628 48832 8634
rect 48780 8570 48832 8576
rect 48884 8498 48912 9318
rect 48976 8838 49004 11886
rect 49068 8974 49096 12406
rect 49252 12170 49280 13874
rect 49240 12164 49292 12170
rect 49240 12106 49292 12112
rect 49344 11762 49372 15846
rect 49332 11756 49384 11762
rect 49332 11698 49384 11704
rect 49344 11082 49372 11698
rect 49332 11076 49384 11082
rect 49332 11018 49384 11024
rect 49240 10804 49292 10810
rect 49240 10746 49292 10752
rect 49252 10062 49280 10746
rect 49436 10606 49464 15982
rect 49620 15638 49648 21966
rect 49712 21418 49740 22034
rect 49804 21690 49832 22034
rect 49896 21894 49924 22986
rect 49988 22506 50016 24092
rect 49976 22500 50028 22506
rect 49976 22442 50028 22448
rect 49976 22228 50028 22234
rect 49976 22170 50028 22176
rect 49884 21888 49936 21894
rect 49884 21830 49936 21836
rect 49792 21684 49844 21690
rect 49988 21672 50016 22170
rect 50080 21690 50108 24142
rect 50540 23730 50568 25638
rect 50816 24818 50844 26250
rect 51092 26042 51120 26336
rect 51276 26234 51304 26862
rect 52092 26784 52144 26790
rect 52092 26726 52144 26732
rect 51540 26580 51592 26586
rect 51540 26522 51592 26528
rect 51356 26376 51408 26382
rect 51356 26318 51408 26324
rect 51184 26206 51304 26234
rect 51080 26036 51132 26042
rect 51080 25978 51132 25984
rect 51184 25922 51212 26206
rect 51368 26042 51396 26318
rect 51448 26240 51500 26246
rect 51448 26182 51500 26188
rect 51356 26036 51408 26042
rect 51356 25978 51408 25984
rect 51184 25906 51304 25922
rect 51172 25900 51304 25906
rect 51224 25894 51304 25900
rect 51172 25842 51224 25848
rect 51172 25764 51224 25770
rect 51172 25706 51224 25712
rect 51080 25152 51132 25158
rect 51080 25094 51132 25100
rect 50896 24880 50948 24886
rect 50896 24822 50948 24828
rect 50804 24812 50856 24818
rect 50724 24772 50804 24800
rect 50724 23730 50752 24772
rect 50804 24754 50856 24760
rect 50908 24698 50936 24822
rect 50816 24670 50936 24698
rect 50528 23724 50580 23730
rect 50528 23666 50580 23672
rect 50712 23724 50764 23730
rect 50712 23666 50764 23672
rect 50252 23656 50304 23662
rect 50252 23598 50304 23604
rect 50160 22976 50212 22982
rect 50160 22918 50212 22924
rect 50172 22642 50200 22918
rect 50160 22636 50212 22642
rect 50160 22578 50212 22584
rect 50160 22432 50212 22438
rect 50160 22374 50212 22380
rect 50172 22234 50200 22374
rect 50160 22228 50212 22234
rect 50160 22170 50212 22176
rect 50160 21888 50212 21894
rect 50160 21830 50212 21836
rect 49792 21626 49844 21632
rect 49896 21644 50016 21672
rect 50068 21684 50120 21690
rect 49700 21412 49752 21418
rect 49700 21354 49752 21360
rect 49698 21312 49754 21321
rect 49698 21247 49754 21256
rect 49712 18834 49740 21247
rect 49700 18828 49752 18834
rect 49700 18770 49752 18776
rect 49712 17134 49740 18770
rect 49700 17128 49752 17134
rect 49700 17070 49752 17076
rect 49700 16516 49752 16522
rect 49700 16458 49752 16464
rect 49712 16425 49740 16458
rect 49698 16416 49754 16425
rect 49698 16351 49754 16360
rect 49712 16182 49740 16351
rect 49700 16176 49752 16182
rect 49700 16118 49752 16124
rect 49896 15706 49924 21644
rect 50068 21626 50120 21632
rect 49976 21548 50028 21554
rect 49976 21490 50028 21496
rect 50068 21548 50120 21554
rect 50068 21490 50120 21496
rect 49988 20942 50016 21490
rect 50080 21418 50108 21490
rect 50068 21412 50120 21418
rect 50068 21354 50120 21360
rect 49976 20936 50028 20942
rect 49976 20878 50028 20884
rect 49976 18760 50028 18766
rect 49976 18702 50028 18708
rect 49988 18426 50016 18702
rect 49976 18420 50028 18426
rect 49976 18362 50028 18368
rect 50080 17066 50108 21354
rect 50068 17060 50120 17066
rect 50068 17002 50120 17008
rect 49976 16788 50028 16794
rect 49976 16730 50028 16736
rect 49988 15910 50016 16730
rect 50080 16522 50108 17002
rect 50068 16516 50120 16522
rect 50068 16458 50120 16464
rect 49976 15904 50028 15910
rect 49976 15846 50028 15852
rect 49884 15700 49936 15706
rect 49884 15642 49936 15648
rect 49608 15632 49660 15638
rect 49608 15574 49660 15580
rect 49896 15570 49924 15642
rect 49884 15564 49936 15570
rect 49884 15506 49936 15512
rect 49700 14952 49752 14958
rect 49700 14894 49752 14900
rect 49516 14816 49568 14822
rect 49514 14784 49516 14793
rect 49568 14784 49570 14793
rect 49514 14719 49570 14728
rect 49424 10600 49476 10606
rect 49424 10542 49476 10548
rect 49424 10464 49476 10470
rect 49424 10406 49476 10412
rect 49332 10260 49384 10266
rect 49332 10202 49384 10208
rect 49240 10056 49292 10062
rect 49160 10016 49240 10044
rect 49160 9654 49188 10016
rect 49240 9998 49292 10004
rect 49344 9994 49372 10202
rect 49436 10130 49464 10406
rect 49424 10124 49476 10130
rect 49424 10066 49476 10072
rect 49332 9988 49384 9994
rect 49332 9930 49384 9936
rect 49148 9648 49200 9654
rect 49148 9590 49200 9596
rect 49528 9586 49556 14719
rect 49712 14482 49740 14894
rect 49896 14634 49924 15506
rect 49976 15360 50028 15366
rect 49976 15302 50028 15308
rect 49804 14606 49924 14634
rect 49700 14476 49752 14482
rect 49700 14418 49752 14424
rect 49804 12434 49832 14606
rect 49884 14476 49936 14482
rect 49884 14418 49936 14424
rect 49896 13802 49924 14418
rect 49884 13796 49936 13802
rect 49884 13738 49936 13744
rect 49712 12406 49832 12434
rect 49712 11762 49740 12406
rect 49988 11762 50016 15302
rect 49700 11756 49752 11762
rect 49700 11698 49752 11704
rect 49976 11756 50028 11762
rect 49976 11698 50028 11704
rect 49712 11354 49740 11698
rect 49884 11688 49936 11694
rect 49884 11630 49936 11636
rect 49700 11348 49752 11354
rect 49700 11290 49752 11296
rect 49608 10464 49660 10470
rect 49608 10406 49660 10412
rect 49516 9580 49568 9586
rect 49516 9522 49568 9528
rect 49528 9178 49556 9522
rect 49516 9172 49568 9178
rect 49516 9114 49568 9120
rect 49620 9042 49648 10406
rect 49700 9920 49752 9926
rect 49700 9862 49752 9868
rect 49792 9920 49844 9926
rect 49792 9862 49844 9868
rect 49712 9654 49740 9862
rect 49700 9648 49752 9654
rect 49700 9590 49752 9596
rect 49698 9344 49754 9353
rect 49698 9279 49754 9288
rect 49712 9178 49740 9279
rect 49700 9172 49752 9178
rect 49700 9114 49752 9120
rect 49698 9072 49754 9081
rect 49608 9036 49660 9042
rect 49698 9007 49700 9016
rect 49608 8978 49660 8984
rect 49752 9007 49754 9016
rect 49700 8978 49752 8984
rect 49056 8968 49108 8974
rect 49056 8910 49108 8916
rect 49698 8936 49754 8945
rect 49698 8871 49700 8880
rect 49752 8871 49754 8880
rect 49700 8842 49752 8848
rect 48964 8832 49016 8838
rect 48964 8774 49016 8780
rect 48872 8492 48924 8498
rect 48872 8434 48924 8440
rect 48976 8430 49004 8774
rect 49804 8498 49832 9862
rect 49896 9178 49924 11630
rect 50080 10266 50108 16458
rect 50172 16250 50200 21830
rect 50264 21078 50292 23598
rect 50528 23588 50580 23594
rect 50528 23530 50580 23536
rect 50344 21684 50396 21690
rect 50344 21626 50396 21632
rect 50252 21072 50304 21078
rect 50252 21014 50304 21020
rect 50252 20800 50304 20806
rect 50252 20742 50304 20748
rect 50264 19922 50292 20742
rect 50252 19916 50304 19922
rect 50252 19858 50304 19864
rect 50252 18284 50304 18290
rect 50252 18226 50304 18232
rect 50264 17814 50292 18226
rect 50252 17808 50304 17814
rect 50252 17750 50304 17756
rect 50264 17542 50292 17750
rect 50356 17610 50384 21626
rect 50436 21344 50488 21350
rect 50540 21321 50568 23530
rect 50620 23112 50672 23118
rect 50620 23054 50672 23060
rect 50632 22778 50660 23054
rect 50712 22976 50764 22982
rect 50712 22918 50764 22924
rect 50620 22772 50672 22778
rect 50620 22714 50672 22720
rect 50632 21894 50660 22714
rect 50724 22273 50752 22918
rect 50710 22264 50766 22273
rect 50710 22199 50766 22208
rect 50620 21888 50672 21894
rect 50620 21830 50672 21836
rect 50436 21286 50488 21292
rect 50526 21312 50582 21321
rect 50448 19854 50476 21286
rect 50526 21247 50582 21256
rect 50528 21004 50580 21010
rect 50528 20946 50580 20952
rect 50540 19854 50568 20946
rect 50436 19848 50488 19854
rect 50436 19790 50488 19796
rect 50528 19848 50580 19854
rect 50528 19790 50580 19796
rect 50540 19718 50568 19790
rect 50528 19712 50580 19718
rect 50528 19654 50580 19660
rect 50540 18816 50568 19654
rect 50448 18788 50568 18816
rect 50448 18290 50476 18788
rect 50528 18692 50580 18698
rect 50528 18634 50580 18640
rect 50540 18426 50568 18634
rect 50528 18420 50580 18426
rect 50528 18362 50580 18368
rect 50436 18284 50488 18290
rect 50436 18226 50488 18232
rect 50620 18216 50672 18222
rect 50620 18158 50672 18164
rect 50344 17604 50396 17610
rect 50344 17546 50396 17552
rect 50252 17536 50304 17542
rect 50252 17478 50304 17484
rect 50356 17202 50384 17546
rect 50528 17332 50580 17338
rect 50528 17274 50580 17280
rect 50344 17196 50396 17202
rect 50344 17138 50396 17144
rect 50344 16584 50396 16590
rect 50344 16526 50396 16532
rect 50250 16416 50306 16425
rect 50250 16351 50306 16360
rect 50160 16244 50212 16250
rect 50160 16186 50212 16192
rect 50264 16114 50292 16351
rect 50252 16108 50304 16114
rect 50252 16050 50304 16056
rect 50356 14396 50384 16526
rect 50434 16280 50490 16289
rect 50434 16215 50490 16224
rect 50448 16114 50476 16215
rect 50436 16108 50488 16114
rect 50436 16050 50488 16056
rect 50434 16008 50490 16017
rect 50434 15943 50436 15952
rect 50488 15943 50490 15952
rect 50436 15914 50488 15920
rect 50436 14544 50488 14550
rect 50434 14512 50436 14521
rect 50488 14512 50490 14521
rect 50434 14447 50490 14456
rect 50436 14408 50488 14414
rect 50356 14368 50436 14396
rect 50436 14350 50488 14356
rect 50252 14272 50304 14278
rect 50436 14272 50488 14278
rect 50252 14214 50304 14220
rect 50342 14240 50398 14249
rect 50160 13864 50212 13870
rect 50160 13806 50212 13812
rect 50172 13530 50200 13806
rect 50160 13524 50212 13530
rect 50160 13466 50212 13472
rect 50264 13394 50292 14214
rect 50436 14214 50488 14220
rect 50342 14175 50398 14184
rect 50252 13388 50304 13394
rect 50252 13330 50304 13336
rect 50356 12850 50384 14175
rect 50344 12844 50396 12850
rect 50344 12786 50396 12792
rect 50344 12436 50396 12442
rect 50344 12378 50396 12384
rect 50356 12170 50384 12378
rect 50344 12164 50396 12170
rect 50344 12106 50396 12112
rect 50448 11218 50476 14214
rect 50436 11212 50488 11218
rect 50436 11154 50488 11160
rect 50068 10260 50120 10266
rect 50068 10202 50120 10208
rect 50160 10124 50212 10130
rect 50160 10066 50212 10072
rect 49976 10056 50028 10062
rect 49976 9998 50028 10004
rect 49988 9722 50016 9998
rect 49976 9716 50028 9722
rect 49976 9658 50028 9664
rect 50068 9512 50120 9518
rect 50068 9454 50120 9460
rect 49976 9444 50028 9450
rect 49976 9386 50028 9392
rect 49884 9172 49936 9178
rect 49884 9114 49936 9120
rect 49792 8492 49844 8498
rect 49792 8434 49844 8440
rect 48964 8424 49016 8430
rect 48964 8366 49016 8372
rect 48504 8288 48556 8294
rect 49988 8242 50016 9386
rect 50080 8294 50108 9454
rect 50172 9382 50200 10066
rect 50344 10056 50396 10062
rect 50344 9998 50396 10004
rect 50436 10056 50488 10062
rect 50436 9998 50488 10004
rect 50356 9722 50384 9998
rect 50344 9716 50396 9722
rect 50344 9658 50396 9664
rect 50252 9648 50304 9654
rect 50252 9590 50304 9596
rect 50342 9616 50398 9625
rect 50160 9376 50212 9382
rect 50160 9318 50212 9324
rect 50158 9208 50214 9217
rect 50158 9143 50214 9152
rect 50172 8838 50200 9143
rect 50160 8832 50212 8838
rect 50160 8774 50212 8780
rect 50172 8537 50200 8774
rect 50158 8528 50214 8537
rect 50158 8463 50214 8472
rect 50264 8430 50292 9590
rect 50342 9551 50344 9560
rect 50396 9551 50398 9560
rect 50344 9522 50396 9528
rect 50448 9518 50476 9998
rect 50436 9512 50488 9518
rect 50436 9454 50488 9460
rect 50344 9444 50396 9450
rect 50344 9386 50396 9392
rect 50356 9110 50384 9386
rect 50344 9104 50396 9110
rect 50344 9046 50396 9052
rect 50344 8900 50396 8906
rect 50344 8842 50396 8848
rect 50252 8424 50304 8430
rect 50252 8366 50304 8372
rect 48504 8230 48556 8236
rect 48516 7954 48544 8230
rect 49896 8214 50016 8242
rect 50068 8288 50120 8294
rect 50068 8230 50120 8236
rect 48504 7948 48556 7954
rect 48504 7890 48556 7896
rect 48228 7812 48280 7818
rect 48228 7754 48280 7760
rect 49896 7410 49924 8214
rect 49976 8084 50028 8090
rect 49976 8026 50028 8032
rect 49988 7478 50016 8026
rect 50080 7478 50108 8230
rect 50264 8090 50292 8366
rect 50252 8084 50304 8090
rect 50252 8026 50304 8032
rect 49976 7472 50028 7478
rect 49976 7414 50028 7420
rect 50068 7472 50120 7478
rect 50068 7414 50120 7420
rect 49884 7404 49936 7410
rect 49884 7346 49936 7352
rect 49700 7200 49752 7206
rect 49700 7142 49752 7148
rect 49712 6798 49740 7142
rect 49896 6934 49924 7346
rect 49884 6928 49936 6934
rect 49884 6870 49936 6876
rect 49792 6860 49844 6866
rect 49792 6802 49844 6808
rect 49700 6792 49752 6798
rect 49700 6734 49752 6740
rect 49056 6656 49108 6662
rect 49056 6598 49108 6604
rect 49700 6656 49752 6662
rect 49700 6598 49752 6604
rect 49068 6390 49096 6598
rect 49712 6390 49740 6598
rect 49056 6384 49108 6390
rect 49056 6326 49108 6332
rect 49700 6384 49752 6390
rect 49700 6326 49752 6332
rect 48044 6248 48096 6254
rect 48044 6190 48096 6196
rect 49516 6112 49568 6118
rect 49516 6054 49568 6060
rect 49528 5574 49556 6054
rect 49516 5568 49568 5574
rect 49516 5510 49568 5516
rect 49700 5568 49752 5574
rect 49700 5510 49752 5516
rect 49528 5234 49556 5510
rect 49712 5234 49740 5510
rect 49516 5228 49568 5234
rect 49516 5170 49568 5176
rect 49700 5228 49752 5234
rect 49700 5170 49752 5176
rect 49804 5166 49832 6802
rect 49976 6384 50028 6390
rect 49976 6326 50028 6332
rect 49792 5160 49844 5166
rect 49792 5102 49844 5108
rect 49516 5024 49568 5030
rect 49516 4966 49568 4972
rect 49528 4826 49556 4966
rect 49516 4820 49568 4826
rect 49516 4762 49568 4768
rect 49988 4554 50016 6326
rect 50080 5914 50108 7414
rect 50356 7410 50384 8842
rect 50344 7404 50396 7410
rect 50344 7346 50396 7352
rect 50448 6798 50476 9454
rect 50540 8634 50568 17274
rect 50632 17270 50660 18158
rect 50724 17338 50752 22199
rect 50816 21622 50844 24670
rect 51092 24138 51120 25094
rect 51080 24132 51132 24138
rect 51080 24074 51132 24080
rect 51080 23520 51132 23526
rect 51080 23462 51132 23468
rect 50896 23316 50948 23322
rect 50896 23258 50948 23264
rect 50908 23050 50936 23258
rect 51092 23118 51120 23462
rect 51080 23112 51132 23118
rect 51080 23054 51132 23060
rect 50896 23044 50948 23050
rect 50896 22986 50948 22992
rect 51184 22642 51212 25706
rect 51276 25294 51304 25894
rect 51264 25288 51316 25294
rect 51264 25230 51316 25236
rect 51368 24818 51396 25978
rect 51460 25906 51488 26182
rect 51448 25900 51500 25906
rect 51448 25842 51500 25848
rect 51552 25838 51580 26522
rect 51816 26308 51868 26314
rect 51816 26250 51868 26256
rect 51540 25832 51592 25838
rect 51540 25774 51592 25780
rect 51552 25498 51580 25774
rect 51828 25702 51856 26250
rect 52104 25906 52132 26726
rect 52380 26466 52408 26862
rect 52736 26784 52788 26790
rect 52736 26726 52788 26732
rect 52380 26450 52500 26466
rect 52276 26444 52328 26450
rect 52380 26444 52512 26450
rect 52380 26438 52460 26444
rect 52276 26386 52328 26392
rect 52460 26386 52512 26392
rect 52288 26330 52316 26386
rect 52748 26382 52776 26726
rect 52736 26376 52788 26382
rect 52288 26314 52500 26330
rect 52736 26318 52788 26324
rect 53748 26376 53800 26382
rect 53748 26318 53800 26324
rect 52288 26308 52512 26314
rect 52288 26302 52460 26308
rect 52460 26250 52512 26256
rect 53012 26308 53064 26314
rect 53012 26250 53064 26256
rect 52552 25968 52604 25974
rect 52552 25910 52604 25916
rect 52092 25900 52144 25906
rect 52092 25842 52144 25848
rect 51816 25696 51868 25702
rect 51814 25664 51816 25673
rect 51868 25664 51870 25673
rect 51814 25599 51870 25608
rect 51540 25492 51592 25498
rect 51540 25434 51592 25440
rect 51908 25492 51960 25498
rect 51908 25434 51960 25440
rect 51724 25288 51776 25294
rect 51724 25230 51776 25236
rect 51736 24954 51764 25230
rect 51724 24948 51776 24954
rect 51724 24890 51776 24896
rect 51356 24812 51408 24818
rect 51356 24754 51408 24760
rect 51920 23322 51948 25434
rect 52368 25424 52420 25430
rect 52368 25366 52420 25372
rect 52000 25288 52052 25294
rect 52000 25230 52052 25236
rect 52012 24954 52040 25230
rect 52276 25220 52328 25226
rect 52276 25162 52328 25168
rect 52000 24948 52052 24954
rect 52000 24890 52052 24896
rect 52092 24812 52144 24818
rect 52092 24754 52144 24760
rect 52104 24342 52132 24754
rect 52092 24336 52144 24342
rect 52092 24278 52144 24284
rect 52104 23866 52132 24278
rect 52092 23860 52144 23866
rect 52092 23802 52144 23808
rect 51540 23316 51592 23322
rect 51540 23258 51592 23264
rect 51908 23316 51960 23322
rect 51908 23258 51960 23264
rect 51552 23118 51580 23258
rect 52288 23118 52316 25162
rect 52380 24818 52408 25366
rect 52368 24812 52420 24818
rect 52368 24754 52420 24760
rect 52380 24274 52408 24754
rect 52564 24750 52592 25910
rect 53024 25838 53052 26250
rect 53760 26042 53788 26318
rect 53748 26036 53800 26042
rect 53748 25978 53800 25984
rect 53012 25832 53064 25838
rect 53012 25774 53064 25780
rect 52552 24744 52604 24750
rect 52552 24686 52604 24692
rect 52368 24268 52420 24274
rect 52368 24210 52420 24216
rect 52564 24070 52592 24686
rect 53024 24682 53052 25774
rect 53656 25492 53708 25498
rect 53656 25434 53708 25440
rect 53380 25288 53432 25294
rect 53380 25230 53432 25236
rect 53472 25288 53524 25294
rect 53472 25230 53524 25236
rect 53564 25288 53616 25294
rect 53564 25230 53616 25236
rect 53196 25152 53248 25158
rect 53196 25094 53248 25100
rect 53208 24886 53236 25094
rect 53196 24880 53248 24886
rect 53196 24822 53248 24828
rect 53392 24750 53420 25230
rect 53380 24744 53432 24750
rect 53300 24704 53380 24732
rect 53012 24676 53064 24682
rect 53012 24618 53064 24624
rect 52920 24200 52972 24206
rect 52920 24142 52972 24148
rect 52552 24064 52604 24070
rect 52552 24006 52604 24012
rect 52564 23798 52592 24006
rect 52552 23792 52604 23798
rect 52552 23734 52604 23740
rect 52932 23730 52960 24142
rect 53024 24138 53052 24618
rect 53300 24410 53328 24704
rect 53380 24686 53432 24692
rect 53484 24410 53512 25230
rect 53576 24954 53604 25230
rect 53564 24948 53616 24954
rect 53564 24890 53616 24896
rect 53288 24404 53340 24410
rect 53288 24346 53340 24352
rect 53472 24404 53524 24410
rect 53472 24346 53524 24352
rect 53012 24132 53064 24138
rect 53012 24074 53064 24080
rect 52920 23724 52972 23730
rect 52920 23666 52972 23672
rect 52932 23186 52960 23666
rect 52920 23180 52972 23186
rect 52920 23122 52972 23128
rect 51540 23112 51592 23118
rect 51540 23054 51592 23060
rect 52276 23112 52328 23118
rect 53196 23112 53248 23118
rect 52328 23072 52408 23100
rect 52276 23054 52328 23060
rect 51540 22976 51592 22982
rect 51540 22918 51592 22924
rect 51552 22642 51580 22918
rect 50988 22636 51040 22642
rect 50988 22578 51040 22584
rect 51172 22636 51224 22642
rect 51172 22578 51224 22584
rect 51540 22636 51592 22642
rect 51540 22578 51592 22584
rect 51000 22098 51028 22578
rect 51356 22568 51408 22574
rect 51356 22510 51408 22516
rect 50988 22092 51040 22098
rect 50988 22034 51040 22040
rect 50804 21616 50856 21622
rect 50804 21558 50856 21564
rect 50896 21548 50948 21554
rect 50896 21490 50948 21496
rect 50804 21140 50856 21146
rect 50804 21082 50856 21088
rect 50816 20913 50844 21082
rect 50908 21078 50936 21490
rect 50896 21072 50948 21078
rect 50894 21040 50896 21049
rect 50948 21040 50950 21049
rect 50894 20975 50950 20984
rect 50896 20936 50948 20942
rect 50802 20904 50858 20913
rect 50896 20878 50948 20884
rect 50802 20839 50858 20848
rect 50804 20800 50856 20806
rect 50804 20742 50856 20748
rect 50816 20534 50844 20742
rect 50804 20528 50856 20534
rect 50804 20470 50856 20476
rect 50908 20058 50936 20878
rect 50804 20052 50856 20058
rect 50804 19994 50856 20000
rect 50896 20052 50948 20058
rect 50896 19994 50948 20000
rect 50816 19854 50844 19994
rect 50804 19848 50856 19854
rect 50804 19790 50856 19796
rect 50804 18284 50856 18290
rect 50804 18226 50856 18232
rect 50816 17882 50844 18226
rect 50804 17876 50856 17882
rect 50804 17818 50856 17824
rect 51000 17746 51028 22034
rect 51368 21690 51396 22510
rect 51356 21684 51408 21690
rect 51356 21626 51408 21632
rect 51172 21548 51224 21554
rect 51172 21490 51224 21496
rect 51184 20913 51212 21490
rect 52184 21480 52236 21486
rect 52184 21422 52236 21428
rect 51632 21412 51684 21418
rect 51632 21354 51684 21360
rect 51540 21072 51592 21078
rect 51540 21014 51592 21020
rect 51170 20904 51226 20913
rect 51170 20839 51226 20848
rect 51080 19916 51132 19922
rect 51080 19858 51132 19864
rect 51092 17882 51120 19858
rect 51080 17876 51132 17882
rect 51080 17818 51132 17824
rect 50988 17740 51040 17746
rect 50988 17682 51040 17688
rect 51080 17604 51132 17610
rect 51080 17546 51132 17552
rect 50712 17332 50764 17338
rect 50712 17274 50764 17280
rect 50620 17264 50672 17270
rect 50620 17206 50672 17212
rect 50632 16250 50660 17206
rect 50724 16590 50752 17274
rect 51092 16674 51120 17546
rect 50804 16652 50856 16658
rect 50804 16594 50856 16600
rect 51000 16646 51120 16674
rect 51184 16658 51212 20839
rect 51356 19168 51408 19174
rect 51356 19110 51408 19116
rect 51264 18828 51316 18834
rect 51264 18770 51316 18776
rect 51276 17082 51304 18770
rect 51368 18086 51396 19110
rect 51448 18624 51500 18630
rect 51448 18566 51500 18572
rect 51460 18358 51488 18566
rect 51448 18352 51500 18358
rect 51448 18294 51500 18300
rect 51356 18080 51408 18086
rect 51356 18022 51408 18028
rect 51276 17054 51396 17082
rect 51264 16992 51316 16998
rect 51264 16934 51316 16940
rect 51172 16652 51224 16658
rect 50712 16584 50764 16590
rect 50712 16526 50764 16532
rect 50816 16250 50844 16594
rect 51000 16522 51028 16646
rect 51172 16594 51224 16600
rect 51276 16522 51304 16934
rect 51368 16658 51396 17054
rect 51356 16652 51408 16658
rect 51356 16594 51408 16600
rect 51460 16590 51488 18294
rect 51448 16584 51500 16590
rect 51448 16526 51500 16532
rect 50988 16516 51040 16522
rect 50988 16458 51040 16464
rect 51264 16516 51316 16522
rect 51264 16458 51316 16464
rect 50896 16448 50948 16454
rect 50894 16416 50896 16425
rect 51080 16448 51132 16454
rect 50948 16416 50950 16425
rect 51276 16425 51304 16458
rect 51448 16448 51500 16454
rect 51080 16390 51132 16396
rect 51262 16416 51318 16425
rect 50894 16351 50950 16360
rect 50620 16244 50672 16250
rect 50620 16186 50672 16192
rect 50804 16244 50856 16250
rect 50804 16186 50856 16192
rect 50894 16144 50950 16153
rect 50894 16079 50896 16088
rect 50948 16079 50950 16088
rect 50896 16050 50948 16056
rect 50712 16040 50764 16046
rect 50712 15982 50764 15988
rect 50620 14816 50672 14822
rect 50620 14758 50672 14764
rect 50632 14278 50660 14758
rect 50620 14272 50672 14278
rect 50620 14214 50672 14220
rect 50620 13864 50672 13870
rect 50620 13806 50672 13812
rect 50632 13326 50660 13806
rect 50620 13320 50672 13326
rect 50724 13308 50752 15982
rect 50896 15632 50948 15638
rect 50896 15574 50948 15580
rect 50908 15502 50936 15574
rect 50896 15496 50948 15502
rect 50896 15438 50948 15444
rect 50908 15366 50936 15438
rect 50988 15428 51040 15434
rect 50988 15370 51040 15376
rect 50896 15360 50948 15366
rect 50896 15302 50948 15308
rect 50804 14612 50856 14618
rect 50804 14554 50856 14560
rect 50816 13870 50844 14554
rect 50804 13864 50856 13870
rect 50804 13806 50856 13812
rect 50724 13280 50844 13308
rect 50620 13262 50672 13268
rect 50712 12164 50764 12170
rect 50712 12106 50764 12112
rect 50724 11898 50752 12106
rect 50712 11892 50764 11898
rect 50712 11834 50764 11840
rect 50620 11212 50672 11218
rect 50620 11154 50672 11160
rect 50528 8628 50580 8634
rect 50528 8570 50580 8576
rect 50528 8492 50580 8498
rect 50528 8434 50580 8440
rect 50540 7274 50568 8434
rect 50632 8430 50660 11154
rect 50712 11008 50764 11014
rect 50712 10950 50764 10956
rect 50724 10062 50752 10950
rect 50816 10742 50844 13280
rect 50908 11218 50936 15302
rect 51000 14482 51028 15370
rect 51092 14618 51120 16390
rect 51448 16390 51500 16396
rect 51262 16351 51318 16360
rect 51172 16108 51224 16114
rect 51172 16050 51224 16056
rect 51356 16108 51408 16114
rect 51356 16050 51408 16056
rect 51184 15706 51212 16050
rect 51172 15700 51224 15706
rect 51172 15642 51224 15648
rect 51080 14612 51132 14618
rect 51080 14554 51132 14560
rect 51368 14550 51396 16050
rect 51356 14544 51408 14550
rect 51356 14486 51408 14492
rect 50988 14476 51040 14482
rect 50988 14418 51040 14424
rect 50988 14340 51040 14346
rect 50988 14282 51040 14288
rect 51000 14113 51028 14282
rect 51264 14272 51316 14278
rect 51262 14240 51264 14249
rect 51316 14240 51318 14249
rect 51262 14175 51318 14184
rect 50986 14104 51042 14113
rect 50986 14039 51042 14048
rect 51368 13870 51396 14486
rect 51356 13864 51408 13870
rect 51356 13806 51408 13812
rect 51172 13728 51224 13734
rect 51172 13670 51224 13676
rect 51184 13462 51212 13670
rect 51172 13456 51224 13462
rect 51172 13398 51224 13404
rect 50988 12640 51040 12646
rect 50988 12582 51040 12588
rect 51000 11898 51028 12582
rect 50988 11892 51040 11898
rect 50988 11834 51040 11840
rect 50988 11756 51040 11762
rect 50988 11698 51040 11704
rect 51000 11354 51028 11698
rect 51184 11558 51212 13398
rect 51460 12434 51488 16390
rect 51552 16114 51580 21014
rect 51644 21010 51672 21354
rect 51632 21004 51684 21010
rect 51632 20946 51684 20952
rect 51644 20058 51672 20946
rect 52196 20330 52224 21422
rect 52380 21418 52408 23072
rect 53196 23054 53248 23060
rect 52552 23044 52604 23050
rect 52552 22986 52604 22992
rect 52564 22098 52592 22986
rect 53012 22976 53064 22982
rect 53012 22918 53064 22924
rect 53024 22710 53052 22918
rect 53012 22704 53064 22710
rect 53012 22646 53064 22652
rect 52644 22568 52696 22574
rect 52644 22510 52696 22516
rect 52736 22568 52788 22574
rect 52736 22510 52788 22516
rect 52552 22092 52604 22098
rect 52552 22034 52604 22040
rect 52656 22030 52684 22510
rect 52748 22094 52776 22510
rect 53208 22234 53236 23054
rect 53196 22228 53248 22234
rect 53196 22170 53248 22176
rect 52920 22094 52972 22098
rect 52748 22092 52972 22094
rect 52748 22066 52920 22092
rect 52644 22024 52696 22030
rect 52644 21966 52696 21972
rect 52368 21412 52420 21418
rect 52368 21354 52420 21360
rect 52276 21004 52328 21010
rect 52276 20946 52328 20952
rect 52288 20398 52316 20946
rect 52748 20602 52776 22066
rect 52920 22034 52972 22040
rect 53012 22024 53064 22030
rect 53012 21966 53064 21972
rect 53378 21992 53434 22001
rect 52828 21956 52880 21962
rect 52828 21898 52880 21904
rect 52840 21622 52868 21898
rect 52828 21616 52880 21622
rect 52828 21558 52880 21564
rect 52920 21412 52972 21418
rect 52920 21354 52972 21360
rect 52932 20942 52960 21354
rect 53024 21078 53052 21966
rect 53378 21927 53380 21936
rect 53432 21927 53434 21936
rect 53380 21898 53432 21904
rect 53392 21690 53420 21898
rect 53380 21684 53432 21690
rect 53380 21626 53432 21632
rect 53012 21072 53064 21078
rect 53012 21014 53064 21020
rect 52920 20936 52972 20942
rect 52920 20878 52972 20884
rect 52828 20868 52880 20874
rect 52828 20810 52880 20816
rect 52736 20596 52788 20602
rect 52736 20538 52788 20544
rect 52748 20466 52776 20538
rect 52736 20460 52788 20466
rect 52736 20402 52788 20408
rect 52276 20392 52328 20398
rect 52276 20334 52328 20340
rect 52184 20324 52236 20330
rect 52184 20266 52236 20272
rect 51632 20052 51684 20058
rect 51632 19994 51684 20000
rect 52196 19854 52224 20266
rect 52184 19848 52236 19854
rect 52288 19836 52316 20334
rect 52840 20058 52868 20810
rect 53012 20800 53064 20806
rect 53012 20742 53064 20748
rect 53104 20800 53156 20806
rect 53104 20742 53156 20748
rect 53024 20534 53052 20742
rect 53012 20528 53064 20534
rect 53012 20470 53064 20476
rect 52828 20052 52880 20058
rect 52828 19994 52880 20000
rect 53116 19854 53144 20742
rect 52368 19848 52420 19854
rect 52288 19808 52368 19836
rect 52184 19790 52236 19796
rect 52368 19790 52420 19796
rect 53104 19848 53156 19854
rect 53104 19790 53156 19796
rect 52368 19712 52420 19718
rect 52368 19654 52420 19660
rect 52092 18896 52144 18902
rect 52144 18844 52316 18850
rect 52092 18838 52316 18844
rect 52104 18834 52316 18838
rect 52104 18828 52328 18834
rect 52104 18822 52276 18828
rect 52276 18770 52328 18776
rect 51908 18692 51960 18698
rect 51908 18634 51960 18640
rect 51920 18154 51948 18634
rect 51908 18148 51960 18154
rect 51908 18090 51960 18096
rect 51908 17672 51960 17678
rect 51908 17614 51960 17620
rect 51724 16652 51776 16658
rect 51724 16594 51776 16600
rect 51630 16144 51686 16153
rect 51540 16108 51592 16114
rect 51630 16079 51686 16088
rect 51540 16050 51592 16056
rect 51540 14884 51592 14890
rect 51540 14826 51592 14832
rect 51552 14414 51580 14826
rect 51540 14408 51592 14414
rect 51540 14350 51592 14356
rect 51540 14000 51592 14006
rect 51540 13942 51592 13948
rect 51552 13802 51580 13942
rect 51540 13796 51592 13802
rect 51540 13738 51592 13744
rect 51368 12406 51488 12434
rect 51080 11552 51132 11558
rect 51080 11494 51132 11500
rect 51172 11552 51224 11558
rect 51172 11494 51224 11500
rect 50988 11348 51040 11354
rect 50988 11290 51040 11296
rect 50896 11212 50948 11218
rect 50896 11154 50948 11160
rect 50896 11076 50948 11082
rect 50896 11018 50948 11024
rect 50804 10736 50856 10742
rect 50804 10678 50856 10684
rect 50804 10464 50856 10470
rect 50804 10406 50856 10412
rect 50816 10062 50844 10406
rect 50712 10056 50764 10062
rect 50712 9998 50764 10004
rect 50804 10056 50856 10062
rect 50804 9998 50856 10004
rect 50712 9716 50764 9722
rect 50712 9658 50764 9664
rect 50724 9110 50752 9658
rect 50908 9586 50936 11018
rect 50988 9920 51040 9926
rect 50988 9862 51040 9868
rect 50896 9580 50948 9586
rect 50896 9522 50948 9528
rect 50804 9444 50856 9450
rect 50804 9386 50856 9392
rect 50712 9104 50764 9110
rect 50712 9046 50764 9052
rect 50816 8634 50844 9386
rect 50896 9172 50948 9178
rect 50896 9114 50948 9120
rect 50908 8634 50936 9114
rect 51000 9042 51028 9862
rect 51092 9110 51120 11494
rect 51368 10810 51396 12406
rect 51552 12102 51580 13738
rect 51540 12096 51592 12102
rect 51540 12038 51592 12044
rect 51356 10804 51408 10810
rect 51356 10746 51408 10752
rect 51368 10198 51396 10746
rect 51448 10736 51500 10742
rect 51448 10678 51500 10684
rect 51356 10192 51408 10198
rect 51356 10134 51408 10140
rect 51460 10062 51488 10678
rect 51644 10198 51672 16079
rect 51736 14414 51764 16594
rect 51920 16114 51948 17614
rect 52380 17338 52408 19654
rect 52460 18964 52512 18970
rect 52460 18906 52512 18912
rect 52472 18290 52500 18906
rect 53012 18624 53064 18630
rect 53012 18566 53064 18572
rect 53024 18290 53052 18566
rect 52460 18284 52512 18290
rect 52460 18226 52512 18232
rect 53012 18284 53064 18290
rect 53012 18226 53064 18232
rect 52472 17746 52500 18226
rect 52552 17876 52604 17882
rect 52552 17818 52604 17824
rect 53196 17876 53248 17882
rect 53196 17818 53248 17824
rect 52460 17740 52512 17746
rect 52460 17682 52512 17688
rect 52368 17332 52420 17338
rect 52368 17274 52420 17280
rect 52380 16250 52408 17274
rect 52564 16640 52592 17818
rect 53208 17678 53236 17818
rect 53196 17672 53248 17678
rect 53194 17640 53196 17649
rect 53248 17640 53250 17649
rect 53012 17604 53064 17610
rect 53194 17575 53250 17584
rect 53012 17546 53064 17552
rect 53024 17338 53052 17546
rect 53012 17332 53064 17338
rect 53012 17274 53064 17280
rect 52472 16612 52592 16640
rect 52644 16652 52696 16658
rect 52368 16244 52420 16250
rect 52368 16186 52420 16192
rect 52472 16114 52500 16612
rect 52644 16594 52696 16600
rect 52552 16516 52604 16522
rect 52552 16458 52604 16464
rect 51908 16108 51960 16114
rect 51908 16050 51960 16056
rect 52276 16108 52328 16114
rect 52276 16050 52328 16056
rect 52460 16108 52512 16114
rect 52460 16050 52512 16056
rect 51816 14816 51868 14822
rect 51816 14758 51868 14764
rect 51724 14408 51776 14414
rect 51724 14350 51776 14356
rect 51736 14074 51764 14350
rect 51724 14068 51776 14074
rect 51724 14010 51776 14016
rect 51828 13734 51856 14758
rect 51920 14113 51948 16050
rect 52288 15570 52316 16050
rect 52276 15564 52328 15570
rect 52276 15506 52328 15512
rect 52564 14346 52592 16458
rect 52656 16250 52684 16594
rect 52644 16244 52696 16250
rect 52644 16186 52696 16192
rect 53392 16182 53420 21626
rect 53668 21146 53696 25434
rect 53944 25158 53972 26998
rect 54208 26920 54260 26926
rect 54208 26862 54260 26868
rect 54484 26920 54536 26926
rect 54484 26862 54536 26868
rect 54220 26586 54248 26862
rect 54208 26580 54260 26586
rect 54208 26522 54260 26528
rect 54496 26518 54524 26862
rect 54484 26512 54536 26518
rect 54484 26454 54536 26460
rect 54496 25430 54524 26454
rect 54484 25424 54536 25430
rect 54484 25366 54536 25372
rect 55588 25220 55640 25226
rect 55588 25162 55640 25168
rect 53932 25152 53984 25158
rect 53932 25094 53984 25100
rect 54484 25152 54536 25158
rect 54484 25094 54536 25100
rect 54496 24750 54524 25094
rect 55600 24954 55628 25162
rect 55772 25152 55824 25158
rect 55772 25094 55824 25100
rect 54760 24948 54812 24954
rect 54760 24890 54812 24896
rect 55588 24948 55640 24954
rect 55588 24890 55640 24896
rect 54484 24744 54536 24750
rect 54484 24686 54536 24692
rect 53748 24064 53800 24070
rect 53748 24006 53800 24012
rect 53760 23662 53788 24006
rect 53748 23656 53800 23662
rect 53748 23598 53800 23604
rect 53760 21894 53788 23598
rect 54496 23186 54524 24686
rect 54772 24206 54800 24890
rect 55784 24886 55812 25094
rect 55772 24880 55824 24886
rect 55772 24822 55824 24828
rect 55312 24812 55364 24818
rect 55312 24754 55364 24760
rect 55404 24812 55456 24818
rect 55404 24754 55456 24760
rect 55220 24608 55272 24614
rect 55220 24550 55272 24556
rect 54944 24268 54996 24274
rect 54944 24210 54996 24216
rect 54760 24200 54812 24206
rect 54760 24142 54812 24148
rect 54956 24138 54984 24210
rect 54944 24132 54996 24138
rect 54944 24074 54996 24080
rect 54956 23730 54984 24074
rect 54576 23724 54628 23730
rect 54576 23666 54628 23672
rect 54944 23724 54996 23730
rect 54944 23666 54996 23672
rect 54484 23180 54536 23186
rect 54484 23122 54536 23128
rect 54496 22710 54524 23122
rect 54588 23118 54616 23666
rect 54576 23112 54628 23118
rect 54576 23054 54628 23060
rect 54484 22704 54536 22710
rect 54484 22646 54536 22652
rect 54588 22522 54616 23054
rect 54852 22976 54904 22982
rect 54852 22918 54904 22924
rect 54864 22642 54892 22918
rect 54852 22636 54904 22642
rect 54852 22578 54904 22584
rect 54116 22500 54168 22506
rect 54116 22442 54168 22448
rect 54496 22494 54616 22522
rect 54128 22094 54156 22442
rect 54496 22438 54524 22494
rect 54484 22432 54536 22438
rect 54484 22374 54536 22380
rect 54128 22066 54340 22094
rect 53748 21888 53800 21894
rect 53748 21830 53800 21836
rect 53760 21622 53788 21830
rect 53748 21616 53800 21622
rect 53748 21558 53800 21564
rect 54208 21344 54260 21350
rect 54208 21286 54260 21292
rect 53656 21140 53708 21146
rect 53656 21082 53708 21088
rect 53668 20262 53696 21082
rect 54220 21010 54248 21286
rect 54208 21004 54260 21010
rect 54208 20946 54260 20952
rect 54220 20330 54248 20946
rect 54208 20324 54260 20330
rect 54208 20266 54260 20272
rect 53656 20256 53708 20262
rect 53656 20198 53708 20204
rect 54024 18692 54076 18698
rect 54024 18634 54076 18640
rect 54036 18426 54064 18634
rect 54024 18420 54076 18426
rect 54024 18362 54076 18368
rect 54116 18352 54168 18358
rect 54116 18294 54168 18300
rect 54024 18284 54076 18290
rect 54024 18226 54076 18232
rect 53932 18080 53984 18086
rect 53932 18022 53984 18028
rect 53944 17542 53972 18022
rect 54036 17882 54064 18226
rect 54024 17876 54076 17882
rect 54024 17818 54076 17824
rect 54128 17814 54156 18294
rect 54116 17808 54168 17814
rect 54116 17750 54168 17756
rect 54312 17762 54340 22066
rect 54496 21690 54524 22374
rect 54956 22030 54984 23666
rect 55128 23520 55180 23526
rect 55128 23462 55180 23468
rect 55140 22642 55168 23462
rect 55232 23322 55260 24550
rect 55324 23798 55352 24754
rect 55416 24410 55444 24754
rect 55404 24404 55456 24410
rect 55404 24346 55456 24352
rect 55588 24132 55640 24138
rect 55588 24074 55640 24080
rect 55312 23792 55364 23798
rect 55312 23734 55364 23740
rect 55600 23322 55628 24074
rect 55220 23316 55272 23322
rect 55220 23258 55272 23264
rect 55312 23316 55364 23322
rect 55312 23258 55364 23264
rect 55588 23316 55640 23322
rect 55588 23258 55640 23264
rect 55128 22636 55180 22642
rect 55128 22578 55180 22584
rect 55232 22506 55260 23258
rect 55324 22982 55352 23258
rect 55312 22976 55364 22982
rect 55312 22918 55364 22924
rect 55404 22976 55456 22982
rect 55404 22918 55456 22924
rect 55416 22710 55444 22918
rect 55404 22704 55456 22710
rect 55404 22646 55456 22652
rect 55220 22500 55272 22506
rect 55220 22442 55272 22448
rect 54944 22024 54996 22030
rect 54944 21966 54996 21972
rect 54484 21684 54536 21690
rect 54484 21626 54536 21632
rect 54496 21554 54524 21626
rect 54956 21554 54984 21966
rect 55312 21616 55364 21622
rect 55312 21558 55364 21564
rect 54484 21548 54536 21554
rect 54484 21490 54536 21496
rect 54852 21548 54904 21554
rect 54852 21490 54904 21496
rect 54944 21548 54996 21554
rect 54944 21490 54996 21496
rect 54576 20868 54628 20874
rect 54576 20810 54628 20816
rect 54588 19786 54616 20810
rect 54864 20466 54892 21490
rect 55128 21344 55180 21350
rect 55128 21286 55180 21292
rect 55220 21344 55272 21350
rect 55220 21286 55272 21292
rect 54944 21140 54996 21146
rect 54944 21082 54996 21088
rect 54852 20460 54904 20466
rect 54852 20402 54904 20408
rect 54864 20058 54892 20402
rect 54956 20262 54984 21082
rect 55140 21078 55168 21286
rect 55128 21072 55180 21078
rect 55128 21014 55180 21020
rect 55232 21010 55260 21286
rect 55220 21004 55272 21010
rect 55220 20946 55272 20952
rect 55324 20890 55352 21558
rect 55496 21412 55548 21418
rect 55496 21354 55548 21360
rect 55232 20862 55352 20890
rect 55508 20874 55536 21354
rect 55496 20868 55548 20874
rect 55128 20800 55180 20806
rect 55128 20742 55180 20748
rect 55140 20466 55168 20742
rect 55232 20602 55260 20862
rect 55496 20810 55548 20816
rect 55220 20596 55272 20602
rect 55220 20538 55272 20544
rect 55128 20460 55180 20466
rect 55128 20402 55180 20408
rect 55128 20324 55180 20330
rect 55128 20266 55180 20272
rect 54944 20256 54996 20262
rect 54944 20198 54996 20204
rect 54852 20052 54904 20058
rect 54852 19994 54904 20000
rect 54576 19780 54628 19786
rect 54576 19722 54628 19728
rect 54956 18902 54984 20198
rect 55140 20097 55168 20266
rect 55126 20088 55182 20097
rect 55126 20023 55182 20032
rect 54484 18896 54536 18902
rect 54484 18838 54536 18844
rect 54944 18896 54996 18902
rect 54944 18838 54996 18844
rect 54392 18760 54444 18766
rect 54392 18702 54444 18708
rect 54404 18086 54432 18702
rect 54496 18222 54524 18838
rect 54668 18760 54720 18766
rect 54668 18702 54720 18708
rect 54484 18216 54536 18222
rect 54484 18158 54536 18164
rect 54392 18080 54444 18086
rect 54392 18022 54444 18028
rect 54680 17882 54708 18702
rect 54668 17876 54720 17882
rect 54668 17818 54720 17824
rect 54312 17734 54432 17762
rect 54116 17672 54168 17678
rect 54114 17640 54116 17649
rect 54168 17640 54170 17649
rect 54114 17575 54170 17584
rect 53932 17536 53984 17542
rect 53932 17478 53984 17484
rect 54116 17536 54168 17542
rect 54116 17478 54168 17484
rect 53944 17202 53972 17478
rect 54128 17270 54156 17478
rect 54116 17264 54168 17270
rect 54116 17206 54168 17212
rect 53932 17196 53984 17202
rect 53932 17138 53984 17144
rect 54208 17196 54260 17202
rect 54208 17138 54260 17144
rect 54116 16992 54168 16998
rect 54116 16934 54168 16940
rect 53748 16448 53800 16454
rect 53748 16390 53800 16396
rect 53840 16448 53892 16454
rect 53840 16390 53892 16396
rect 53760 16289 53788 16390
rect 53746 16280 53802 16289
rect 53746 16215 53802 16224
rect 53380 16176 53432 16182
rect 53380 16118 53432 16124
rect 53392 15706 53420 16118
rect 53852 16114 53880 16390
rect 53840 16108 53892 16114
rect 53840 16050 53892 16056
rect 54024 16040 54076 16046
rect 54024 15982 54076 15988
rect 53380 15700 53432 15706
rect 53380 15642 53432 15648
rect 53392 15473 53420 15642
rect 53378 15464 53434 15473
rect 53378 15399 53434 15408
rect 53840 15428 53892 15434
rect 53010 14376 53066 14385
rect 52092 14340 52144 14346
rect 52092 14282 52144 14288
rect 52552 14340 52604 14346
rect 53010 14311 53066 14320
rect 52552 14282 52604 14288
rect 51906 14104 51962 14113
rect 51906 14039 51962 14048
rect 52104 13938 52132 14282
rect 52184 14272 52236 14278
rect 52184 14214 52236 14220
rect 52196 13938 52224 14214
rect 52276 14068 52328 14074
rect 52276 14010 52328 14016
rect 52092 13932 52144 13938
rect 52092 13874 52144 13880
rect 52184 13932 52236 13938
rect 52184 13874 52236 13880
rect 51816 13728 51868 13734
rect 51816 13670 51868 13676
rect 52288 12434 52316 14010
rect 52564 13802 52592 14282
rect 52552 13796 52604 13802
rect 52552 13738 52604 13744
rect 52368 13728 52420 13734
rect 52368 13670 52420 13676
rect 52380 13462 52408 13670
rect 52368 13456 52420 13462
rect 52368 13398 52420 13404
rect 52196 12406 52316 12434
rect 51816 12300 51868 12306
rect 51816 12242 51868 12248
rect 51724 11076 51776 11082
rect 51724 11018 51776 11024
rect 51736 10810 51764 11018
rect 51724 10804 51776 10810
rect 51724 10746 51776 10752
rect 51828 10742 51856 12242
rect 52000 11756 52052 11762
rect 52000 11698 52052 11704
rect 52012 11626 52040 11698
rect 52000 11620 52052 11626
rect 52000 11562 52052 11568
rect 51908 11552 51960 11558
rect 51908 11494 51960 11500
rect 51816 10736 51868 10742
rect 51816 10678 51868 10684
rect 51828 10266 51856 10678
rect 51816 10260 51868 10266
rect 51816 10202 51868 10208
rect 51632 10192 51684 10198
rect 51632 10134 51684 10140
rect 51264 10056 51316 10062
rect 51448 10056 51500 10062
rect 51316 10016 51396 10044
rect 51264 9998 51316 10004
rect 51264 9920 51316 9926
rect 51264 9862 51316 9868
rect 51172 9716 51224 9722
rect 51172 9658 51224 9664
rect 51184 9450 51212 9658
rect 51172 9444 51224 9450
rect 51172 9386 51224 9392
rect 51080 9104 51132 9110
rect 51080 9046 51132 9052
rect 50988 9036 51040 9042
rect 50988 8978 51040 8984
rect 51276 8974 51304 9862
rect 51368 9586 51396 10016
rect 51448 9998 51500 10004
rect 51540 10056 51592 10062
rect 51540 9998 51592 10004
rect 51724 10056 51776 10062
rect 51724 9998 51776 10004
rect 51448 9920 51500 9926
rect 51448 9862 51500 9868
rect 51356 9580 51408 9586
rect 51356 9522 51408 9528
rect 51460 9450 51488 9862
rect 51448 9444 51500 9450
rect 51448 9386 51500 9392
rect 51080 8968 51132 8974
rect 50986 8936 51042 8945
rect 51264 8968 51316 8974
rect 51132 8928 51212 8956
rect 51080 8910 51132 8916
rect 50986 8871 50988 8880
rect 51040 8871 51042 8880
rect 50988 8842 51040 8848
rect 51184 8634 51212 8928
rect 51264 8910 51316 8916
rect 51356 8832 51408 8838
rect 51356 8774 51408 8780
rect 50804 8628 50856 8634
rect 50804 8570 50856 8576
rect 50896 8628 50948 8634
rect 50896 8570 50948 8576
rect 51172 8628 51224 8634
rect 51172 8570 51224 8576
rect 50712 8560 50764 8566
rect 50712 8502 50764 8508
rect 51080 8560 51132 8566
rect 51080 8502 51132 8508
rect 50620 8424 50672 8430
rect 50620 8366 50672 8372
rect 50632 7954 50660 8366
rect 50620 7948 50672 7954
rect 50620 7890 50672 7896
rect 50528 7268 50580 7274
rect 50528 7210 50580 7216
rect 50436 6792 50488 6798
rect 50436 6734 50488 6740
rect 50448 6458 50476 6734
rect 50436 6452 50488 6458
rect 50436 6394 50488 6400
rect 50068 5908 50120 5914
rect 50068 5850 50120 5856
rect 50344 5908 50396 5914
rect 50344 5850 50396 5856
rect 50080 5642 50108 5850
rect 50356 5710 50384 5850
rect 50448 5710 50476 6394
rect 50724 6254 50752 8502
rect 51092 8378 51120 8502
rect 51264 8492 51316 8498
rect 51264 8434 51316 8440
rect 50908 8350 51120 8378
rect 51276 8362 51304 8434
rect 51264 8356 51316 8362
rect 50908 8294 50936 8350
rect 51264 8298 51316 8304
rect 50896 8288 50948 8294
rect 50896 8230 50948 8236
rect 51276 8090 51304 8298
rect 50804 8084 50856 8090
rect 50804 8026 50856 8032
rect 51264 8084 51316 8090
rect 51264 8026 51316 8032
rect 50816 7002 50844 8026
rect 51172 7404 51224 7410
rect 51172 7346 51224 7352
rect 50804 6996 50856 7002
rect 50804 6938 50856 6944
rect 50712 6248 50764 6254
rect 50712 6190 50764 6196
rect 50724 5710 50752 6190
rect 50816 5710 50844 6938
rect 50988 6860 51040 6866
rect 50988 6802 51040 6808
rect 51000 5914 51028 6802
rect 50988 5908 51040 5914
rect 51040 5868 51120 5896
rect 50988 5850 51040 5856
rect 51092 5778 51120 5868
rect 51080 5772 51132 5778
rect 51080 5714 51132 5720
rect 51184 5710 51212 7346
rect 50344 5704 50396 5710
rect 50344 5646 50396 5652
rect 50436 5704 50488 5710
rect 50436 5646 50488 5652
rect 50712 5704 50764 5710
rect 50712 5646 50764 5652
rect 50804 5704 50856 5710
rect 50804 5646 50856 5652
rect 51172 5704 51224 5710
rect 51172 5646 51224 5652
rect 50068 5636 50120 5642
rect 50068 5578 50120 5584
rect 50988 5228 51040 5234
rect 51184 5216 51212 5646
rect 51040 5188 51212 5216
rect 50988 5170 51040 5176
rect 51000 4690 51028 5170
rect 50988 4684 51040 4690
rect 50988 4626 51040 4632
rect 49976 4548 50028 4554
rect 49976 4490 50028 4496
rect 50344 4548 50396 4554
rect 50344 4490 50396 4496
rect 49056 4480 49108 4486
rect 49056 4422 49108 4428
rect 47768 4208 47820 4214
rect 47768 4150 47820 4156
rect 47124 4072 47176 4078
rect 47124 4014 47176 4020
rect 47676 4072 47728 4078
rect 47676 4014 47728 4020
rect 46756 3732 46808 3738
rect 46756 3674 46808 3680
rect 44824 3596 44876 3602
rect 44824 3538 44876 3544
rect 45008 3596 45060 3602
rect 45008 3538 45060 3544
rect 45284 3596 45336 3602
rect 45284 3538 45336 3544
rect 44548 3460 44600 3466
rect 44548 3402 44600 3408
rect 44272 3188 44324 3194
rect 44272 3130 44324 3136
rect 44836 3058 44864 3538
rect 44916 3528 44968 3534
rect 44916 3470 44968 3476
rect 44928 3126 44956 3470
rect 47780 3466 47808 4150
rect 49068 4078 49096 4422
rect 49056 4072 49108 4078
rect 49056 4014 49108 4020
rect 50356 3738 50384 4490
rect 51080 4072 51132 4078
rect 51080 4014 51132 4020
rect 50344 3732 50396 3738
rect 50344 3674 50396 3680
rect 50356 3466 50384 3674
rect 47768 3460 47820 3466
rect 47768 3402 47820 3408
rect 50344 3460 50396 3466
rect 50344 3402 50396 3408
rect 50804 3392 50856 3398
rect 50804 3334 50856 3340
rect 50988 3392 51040 3398
rect 50988 3334 51040 3340
rect 50816 3126 50844 3334
rect 44916 3120 44968 3126
rect 44916 3062 44968 3068
rect 50804 3120 50856 3126
rect 50804 3062 50856 3068
rect 44180 3052 44232 3058
rect 44180 2994 44232 3000
rect 44824 3052 44876 3058
rect 44824 2994 44876 3000
rect 45560 3052 45612 3058
rect 45560 2994 45612 3000
rect 43352 2848 43404 2854
rect 43352 2790 43404 2796
rect 43536 2848 43588 2854
rect 43536 2790 43588 2796
rect 43364 2446 43392 2790
rect 43548 2514 43576 2790
rect 44192 2650 44220 2994
rect 45008 2848 45060 2854
rect 45008 2790 45060 2796
rect 44180 2644 44232 2650
rect 44180 2586 44232 2592
rect 43536 2508 43588 2514
rect 43536 2450 43588 2456
rect 45020 2446 45048 2790
rect 45572 2650 45600 2994
rect 49792 2916 49844 2922
rect 49792 2858 49844 2864
rect 45836 2848 45888 2854
rect 45836 2790 45888 2796
rect 46480 2848 46532 2854
rect 46480 2790 46532 2796
rect 47124 2848 47176 2854
rect 47124 2790 47176 2796
rect 47768 2848 47820 2854
rect 47768 2790 47820 2796
rect 49056 2848 49108 2854
rect 49056 2790 49108 2796
rect 49700 2848 49752 2854
rect 49700 2790 49752 2796
rect 45560 2644 45612 2650
rect 45560 2586 45612 2592
rect 45100 2508 45152 2514
rect 45100 2450 45152 2456
rect 43260 2440 43312 2446
rect 43260 2382 43312 2388
rect 43352 2440 43404 2446
rect 43352 2382 43404 2388
rect 45008 2440 45060 2446
rect 45008 2382 45060 2388
rect 43364 2038 43392 2382
rect 43812 2304 43864 2310
rect 43812 2246 43864 2252
rect 43352 2032 43404 2038
rect 43352 1974 43404 1980
rect 43824 800 43852 2246
rect 44456 2100 44508 2106
rect 44456 2042 44508 2048
rect 44468 800 44496 2042
rect 45112 800 45140 2450
rect 45848 2446 45876 2790
rect 46492 2446 46520 2790
rect 47136 2446 47164 2790
rect 47780 2446 47808 2790
rect 49068 2446 49096 2790
rect 49712 2582 49740 2790
rect 49700 2576 49752 2582
rect 49700 2518 49752 2524
rect 49804 2446 49832 2858
rect 51000 2650 51028 3334
rect 51092 3058 51120 4014
rect 51368 3738 51396 8774
rect 51460 8090 51488 9386
rect 51448 8084 51500 8090
rect 51448 8026 51500 8032
rect 51552 7936 51580 9998
rect 51736 9722 51764 9998
rect 51724 9716 51776 9722
rect 51724 9658 51776 9664
rect 51632 9648 51684 9654
rect 51630 9616 51632 9625
rect 51684 9616 51686 9625
rect 51630 9551 51686 9560
rect 51632 8900 51684 8906
rect 51632 8842 51684 8848
rect 51644 8498 51672 8842
rect 51632 8492 51684 8498
rect 51632 8434 51684 8440
rect 51724 8492 51776 8498
rect 51724 8434 51776 8440
rect 51736 8378 51764 8434
rect 51460 7908 51580 7936
rect 51644 8350 51764 8378
rect 51460 5846 51488 7908
rect 51540 7812 51592 7818
rect 51540 7754 51592 7760
rect 51552 7546 51580 7754
rect 51540 7540 51592 7546
rect 51540 7482 51592 7488
rect 51644 6866 51672 8350
rect 51724 8288 51776 8294
rect 51724 8230 51776 8236
rect 51736 7410 51764 8230
rect 51828 7954 51856 10202
rect 51920 9382 51948 11494
rect 52012 11150 52040 11562
rect 52000 11144 52052 11150
rect 52000 11086 52052 11092
rect 52092 10600 52144 10606
rect 52092 10542 52144 10548
rect 52000 10192 52052 10198
rect 52000 10134 52052 10140
rect 52012 9722 52040 10134
rect 52104 10062 52132 10542
rect 52196 10198 52224 12406
rect 52644 12164 52696 12170
rect 52644 12106 52696 12112
rect 52276 12096 52328 12102
rect 52276 12038 52328 12044
rect 52288 11762 52316 12038
rect 52276 11756 52328 11762
rect 52276 11698 52328 11704
rect 52460 11552 52512 11558
rect 52460 11494 52512 11500
rect 52184 10192 52236 10198
rect 52184 10134 52236 10140
rect 52092 10056 52144 10062
rect 52092 9998 52144 10004
rect 52368 10056 52420 10062
rect 52368 9998 52420 10004
rect 52184 9988 52236 9994
rect 52184 9930 52236 9936
rect 52000 9716 52052 9722
rect 52000 9658 52052 9664
rect 51908 9376 51960 9382
rect 51908 9318 51960 9324
rect 52012 8362 52040 9658
rect 52196 8566 52224 9930
rect 52380 9450 52408 9998
rect 52368 9444 52420 9450
rect 52368 9386 52420 9392
rect 52184 8560 52236 8566
rect 52184 8502 52236 8508
rect 52000 8356 52052 8362
rect 52000 8298 52052 8304
rect 52184 8084 52236 8090
rect 52184 8026 52236 8032
rect 51816 7948 51868 7954
rect 51816 7890 51868 7896
rect 52196 7410 52224 8026
rect 51724 7404 51776 7410
rect 51724 7346 51776 7352
rect 52184 7404 52236 7410
rect 52184 7346 52236 7352
rect 51632 6860 51684 6866
rect 51632 6802 51684 6808
rect 51644 6322 51672 6802
rect 51908 6724 51960 6730
rect 51908 6666 51960 6672
rect 51632 6316 51684 6322
rect 51632 6258 51684 6264
rect 51448 5840 51500 5846
rect 51500 5800 51580 5828
rect 51448 5782 51500 5788
rect 51448 5568 51500 5574
rect 51448 5510 51500 5516
rect 51460 5302 51488 5510
rect 51448 5296 51500 5302
rect 51448 5238 51500 5244
rect 51552 4554 51580 5800
rect 51724 5636 51776 5642
rect 51724 5578 51776 5584
rect 51736 5166 51764 5578
rect 51920 5234 51948 6666
rect 52472 6118 52500 11494
rect 52656 11150 52684 12106
rect 52828 11824 52880 11830
rect 52828 11766 52880 11772
rect 52840 11150 52868 11766
rect 53024 11762 53052 14311
rect 53012 11756 53064 11762
rect 53012 11698 53064 11704
rect 52644 11144 52696 11150
rect 52644 11086 52696 11092
rect 52828 11144 52880 11150
rect 52828 11086 52880 11092
rect 53024 11082 53052 11698
rect 53012 11076 53064 11082
rect 53012 11018 53064 11024
rect 53392 10674 53420 15399
rect 53840 15370 53892 15376
rect 53564 14612 53616 14618
rect 53564 14554 53616 14560
rect 53576 14414 53604 14554
rect 53564 14408 53616 14414
rect 53564 14350 53616 14356
rect 53472 14340 53524 14346
rect 53472 14282 53524 14288
rect 53484 13938 53512 14282
rect 53472 13932 53524 13938
rect 53472 13874 53524 13880
rect 53852 13394 53880 15370
rect 54036 15026 54064 15982
rect 54024 15020 54076 15026
rect 54024 14962 54076 14968
rect 54036 14006 54064 14962
rect 54128 14804 54156 16934
rect 54220 16590 54248 17138
rect 54208 16584 54260 16590
rect 54208 16526 54260 16532
rect 54220 15502 54248 16526
rect 54404 15586 54432 17734
rect 54576 17672 54628 17678
rect 54576 17614 54628 17620
rect 54484 17264 54536 17270
rect 54484 17206 54536 17212
rect 54312 15558 54432 15586
rect 54208 15496 54260 15502
rect 54208 15438 54260 15444
rect 54208 14816 54260 14822
rect 54128 14776 54208 14804
rect 54208 14758 54260 14764
rect 54220 14550 54248 14758
rect 54208 14544 54260 14550
rect 54208 14486 54260 14492
rect 54116 14272 54168 14278
rect 54116 14214 54168 14220
rect 54024 14000 54076 14006
rect 54024 13942 54076 13948
rect 53932 13728 53984 13734
rect 53932 13670 53984 13676
rect 53944 13530 53972 13670
rect 53932 13524 53984 13530
rect 53932 13466 53984 13472
rect 53840 13388 53892 13394
rect 53840 13330 53892 13336
rect 54036 12306 54064 13942
rect 54128 13326 54156 14214
rect 54220 14074 54248 14486
rect 54312 14226 54340 15558
rect 54496 15434 54524 17206
rect 54588 17202 54616 17614
rect 54576 17196 54628 17202
rect 54628 17156 54708 17184
rect 54576 17138 54628 17144
rect 54576 16448 54628 16454
rect 54576 16390 54628 16396
rect 54588 16182 54616 16390
rect 54576 16176 54628 16182
rect 54576 16118 54628 16124
rect 54680 15502 54708 17156
rect 54760 16992 54812 16998
rect 54760 16934 54812 16940
rect 54772 16590 54800 16934
rect 54956 16590 54984 18838
rect 55036 17604 55088 17610
rect 55036 17546 55088 17552
rect 55048 16590 55076 17546
rect 54760 16584 54812 16590
rect 54760 16526 54812 16532
rect 54944 16584 54996 16590
rect 54944 16526 54996 16532
rect 55036 16584 55088 16590
rect 55036 16526 55088 16532
rect 54956 16250 54984 16526
rect 54944 16244 54996 16250
rect 54944 16186 54996 16192
rect 55048 16046 55076 16526
rect 55036 16040 55088 16046
rect 55036 15982 55088 15988
rect 54944 15564 54996 15570
rect 54944 15506 54996 15512
rect 54668 15496 54720 15502
rect 54668 15438 54720 15444
rect 54484 15428 54536 15434
rect 54484 15370 54536 15376
rect 54956 14414 54984 15506
rect 54576 14408 54628 14414
rect 54760 14408 54812 14414
rect 54576 14350 54628 14356
rect 54758 14376 54760 14385
rect 54944 14408 54996 14414
rect 54812 14376 54814 14385
rect 54312 14198 54524 14226
rect 54208 14068 54260 14074
rect 54208 14010 54260 14016
rect 54116 13320 54168 13326
rect 54116 13262 54168 13268
rect 54496 12850 54524 14198
rect 54484 12844 54536 12850
rect 54484 12786 54536 12792
rect 54024 12300 54076 12306
rect 54024 12242 54076 12248
rect 54208 12300 54260 12306
rect 54208 12242 54260 12248
rect 54116 12096 54168 12102
rect 54116 12038 54168 12044
rect 53564 11212 53616 11218
rect 54128 11200 54156 12038
rect 54220 11762 54248 12242
rect 54392 11824 54444 11830
rect 54392 11766 54444 11772
rect 54208 11756 54260 11762
rect 54208 11698 54260 11704
rect 54208 11212 54260 11218
rect 54128 11172 54208 11200
rect 53564 11154 53616 11160
rect 54208 11154 54260 11160
rect 53104 10668 53156 10674
rect 53104 10610 53156 10616
rect 53380 10668 53432 10674
rect 53380 10610 53432 10616
rect 52920 9988 52972 9994
rect 52920 9930 52972 9936
rect 52932 9722 52960 9930
rect 53012 9920 53064 9926
rect 53012 9862 53064 9868
rect 52920 9716 52972 9722
rect 52920 9658 52972 9664
rect 53024 9586 53052 9862
rect 53012 9580 53064 9586
rect 53012 9522 53064 9528
rect 52920 8356 52972 8362
rect 52920 8298 52972 8304
rect 52932 7750 52960 8298
rect 52920 7744 52972 7750
rect 52920 7686 52972 7692
rect 52552 7200 52604 7206
rect 52552 7142 52604 7148
rect 52460 6112 52512 6118
rect 52460 6054 52512 6060
rect 52092 5568 52144 5574
rect 52092 5510 52144 5516
rect 51908 5228 51960 5234
rect 51960 5188 52040 5216
rect 51908 5170 51960 5176
rect 51724 5160 51776 5166
rect 51724 5102 51776 5108
rect 52012 4622 52040 5188
rect 52104 5166 52132 5510
rect 52092 5160 52144 5166
rect 52092 5102 52144 5108
rect 52104 4690 52132 5102
rect 52564 5030 52592 7142
rect 52828 6112 52880 6118
rect 52828 6054 52880 6060
rect 52840 5234 52868 6054
rect 52932 5710 52960 7686
rect 52920 5704 52972 5710
rect 52920 5646 52972 5652
rect 52828 5228 52880 5234
rect 52828 5170 52880 5176
rect 52552 5024 52604 5030
rect 52552 4966 52604 4972
rect 52564 4758 52592 4966
rect 52552 4752 52604 4758
rect 52552 4694 52604 4700
rect 52092 4684 52144 4690
rect 52092 4626 52144 4632
rect 52000 4616 52052 4622
rect 52000 4558 52052 4564
rect 51540 4548 51592 4554
rect 51540 4490 51592 4496
rect 52104 4078 52132 4626
rect 52092 4072 52144 4078
rect 52092 4014 52144 4020
rect 51448 4004 51500 4010
rect 51448 3946 51500 3952
rect 51356 3732 51408 3738
rect 51356 3674 51408 3680
rect 51460 3058 51488 3946
rect 52932 3534 52960 5646
rect 53116 5370 53144 10610
rect 53196 9376 53248 9382
rect 53194 9344 53196 9353
rect 53248 9344 53250 9353
rect 53194 9279 53250 9288
rect 53472 8492 53524 8498
rect 53472 8434 53524 8440
rect 53288 8288 53340 8294
rect 53288 8230 53340 8236
rect 53300 7818 53328 8230
rect 53380 7948 53432 7954
rect 53380 7890 53432 7896
rect 53288 7812 53340 7818
rect 53288 7754 53340 7760
rect 53392 7274 53420 7890
rect 53484 7546 53512 8434
rect 53576 8362 53604 11154
rect 54220 10674 54248 11154
rect 54404 11150 54432 11766
rect 54484 11688 54536 11694
rect 54484 11630 54536 11636
rect 54496 11354 54524 11630
rect 54484 11348 54536 11354
rect 54484 11290 54536 11296
rect 54588 11286 54616 14350
rect 54944 14350 54996 14356
rect 54758 14311 54814 14320
rect 54944 13864 54996 13870
rect 54944 13806 54996 13812
rect 54956 12102 54984 13806
rect 54944 12096 54996 12102
rect 54944 12038 54996 12044
rect 54956 11830 54984 12038
rect 54944 11824 54996 11830
rect 54944 11766 54996 11772
rect 55036 11552 55088 11558
rect 55036 11494 55088 11500
rect 54576 11280 54628 11286
rect 54576 11222 54628 11228
rect 54392 11144 54444 11150
rect 54392 11086 54444 11092
rect 54300 11076 54352 11082
rect 54300 11018 54352 11024
rect 54312 10742 54340 11018
rect 54300 10736 54352 10742
rect 54300 10678 54352 10684
rect 54588 10674 54616 11222
rect 55048 11150 55076 11494
rect 54760 11144 54812 11150
rect 54760 11086 54812 11092
rect 55036 11144 55088 11150
rect 55036 11086 55088 11092
rect 54772 10810 54800 11086
rect 54944 11076 54996 11082
rect 54944 11018 54996 11024
rect 54760 10804 54812 10810
rect 54760 10746 54812 10752
rect 54208 10668 54260 10674
rect 54208 10610 54260 10616
rect 54576 10668 54628 10674
rect 54576 10610 54628 10616
rect 54852 10464 54904 10470
rect 54852 10406 54904 10412
rect 54864 10062 54892 10406
rect 54852 10056 54904 10062
rect 54852 9998 54904 10004
rect 54208 9988 54260 9994
rect 54208 9930 54260 9936
rect 54220 9586 54248 9930
rect 54392 9920 54444 9926
rect 54392 9862 54444 9868
rect 54208 9580 54260 9586
rect 54208 9522 54260 9528
rect 54404 9518 54432 9862
rect 54956 9738 54984 11018
rect 55048 11014 55076 11086
rect 55036 11008 55088 11014
rect 55036 10950 55088 10956
rect 54772 9722 54984 9738
rect 54772 9716 54996 9722
rect 54772 9710 54944 9716
rect 54484 9580 54536 9586
rect 54484 9522 54536 9528
rect 54668 9580 54720 9586
rect 54668 9522 54720 9528
rect 54392 9512 54444 9518
rect 54496 9489 54524 9522
rect 54392 9454 54444 9460
rect 54482 9480 54538 9489
rect 54482 9415 54538 9424
rect 53564 8356 53616 8362
rect 53564 8298 53616 8304
rect 53472 7540 53524 7546
rect 53472 7482 53524 7488
rect 53380 7268 53432 7274
rect 53380 7210 53432 7216
rect 53288 6248 53340 6254
rect 53288 6190 53340 6196
rect 53300 5914 53328 6190
rect 53288 5908 53340 5914
rect 53288 5850 53340 5856
rect 53392 5710 53420 7210
rect 53576 7206 53604 8298
rect 54680 7954 54708 9522
rect 54024 7948 54076 7954
rect 54024 7890 54076 7896
rect 54668 7948 54720 7954
rect 54668 7890 54720 7896
rect 53656 7744 53708 7750
rect 53656 7686 53708 7692
rect 53668 7410 53696 7686
rect 53748 7540 53800 7546
rect 53748 7482 53800 7488
rect 53760 7410 53788 7482
rect 53656 7404 53708 7410
rect 53656 7346 53708 7352
rect 53748 7404 53800 7410
rect 53748 7346 53800 7352
rect 53840 7404 53892 7410
rect 54036 7392 54064 7890
rect 54208 7540 54260 7546
rect 54208 7482 54260 7488
rect 53892 7364 54064 7392
rect 53840 7346 53892 7352
rect 53564 7200 53616 7206
rect 53564 7142 53616 7148
rect 53668 6322 53696 7346
rect 54036 6322 54064 7364
rect 54116 7404 54168 7410
rect 54116 7346 54168 7352
rect 54128 7002 54156 7346
rect 54220 7274 54248 7482
rect 54772 7410 54800 9710
rect 54944 9658 54996 9664
rect 54944 9580 54996 9586
rect 54944 9522 54996 9528
rect 54852 8492 54904 8498
rect 54852 8434 54904 8440
rect 54864 8090 54892 8434
rect 54852 8084 54904 8090
rect 54852 8026 54904 8032
rect 54956 7886 54984 9522
rect 55048 9489 55076 10950
rect 55034 9480 55090 9489
rect 55034 9415 55090 9424
rect 55036 9376 55088 9382
rect 55036 9318 55088 9324
rect 55048 9178 55076 9318
rect 55036 9172 55088 9178
rect 55036 9114 55088 9120
rect 54944 7880 54996 7886
rect 54944 7822 54996 7828
rect 55036 7744 55088 7750
rect 55036 7686 55088 7692
rect 55048 7546 55076 7686
rect 55036 7540 55088 7546
rect 55036 7482 55088 7488
rect 54760 7404 54812 7410
rect 54760 7346 54812 7352
rect 54208 7268 54260 7274
rect 54208 7210 54260 7216
rect 54116 6996 54168 7002
rect 54116 6938 54168 6944
rect 54220 6322 54248 7210
rect 53656 6316 53708 6322
rect 53656 6258 53708 6264
rect 54024 6316 54076 6322
rect 54024 6258 54076 6264
rect 54208 6316 54260 6322
rect 54208 6258 54260 6264
rect 53656 6112 53708 6118
rect 53656 6054 53708 6060
rect 53748 6112 53800 6118
rect 53748 6054 53800 6060
rect 53380 5704 53432 5710
rect 53380 5646 53432 5652
rect 53104 5364 53156 5370
rect 53104 5306 53156 5312
rect 53392 5166 53420 5646
rect 53564 5636 53616 5642
rect 53564 5578 53616 5584
rect 53380 5160 53432 5166
rect 53380 5102 53432 5108
rect 53576 4826 53604 5578
rect 53564 4820 53616 4826
rect 53564 4762 53616 4768
rect 53668 4622 53696 6054
rect 53760 5574 53788 6054
rect 54036 5778 54064 6258
rect 54024 5772 54076 5778
rect 54024 5714 54076 5720
rect 53748 5568 53800 5574
rect 53748 5510 53800 5516
rect 54772 4690 54800 7346
rect 55140 6458 55168 20023
rect 55232 19786 55260 20538
rect 55508 20466 55536 20810
rect 55968 20806 55996 28358
rect 66314 28316 66622 28325
rect 66314 28314 66320 28316
rect 66376 28314 66400 28316
rect 66456 28314 66480 28316
rect 66536 28314 66560 28316
rect 66616 28314 66622 28316
rect 66376 28262 66378 28314
rect 66558 28262 66560 28314
rect 66314 28260 66320 28262
rect 66376 28260 66400 28262
rect 66456 28260 66480 28262
rect 66536 28260 66560 28262
rect 66616 28260 66622 28262
rect 66314 28251 66622 28260
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 66314 27228 66622 27237
rect 66314 27226 66320 27228
rect 66376 27226 66400 27228
rect 66456 27226 66480 27228
rect 66536 27226 66560 27228
rect 66616 27226 66622 27228
rect 66376 27174 66378 27226
rect 66558 27174 66560 27226
rect 66314 27172 66320 27174
rect 66376 27172 66400 27174
rect 66456 27172 66480 27174
rect 66536 27172 66560 27174
rect 66616 27172 66622 27174
rect 66314 27163 66622 27172
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 66314 26140 66622 26149
rect 66314 26138 66320 26140
rect 66376 26138 66400 26140
rect 66456 26138 66480 26140
rect 66536 26138 66560 26140
rect 66616 26138 66622 26140
rect 66376 26086 66378 26138
rect 66558 26086 66560 26138
rect 66314 26084 66320 26086
rect 66376 26084 66400 26086
rect 66456 26084 66480 26086
rect 66536 26084 66560 26086
rect 66616 26084 66622 26086
rect 66314 26075 66622 26084
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 66314 25052 66622 25061
rect 66314 25050 66320 25052
rect 66376 25050 66400 25052
rect 66456 25050 66480 25052
rect 66536 25050 66560 25052
rect 66616 25050 66622 25052
rect 66376 24998 66378 25050
rect 66558 24998 66560 25050
rect 66314 24996 66320 24998
rect 66376 24996 66400 24998
rect 66456 24996 66480 24998
rect 66536 24996 66560 24998
rect 66616 24996 66622 24998
rect 66314 24987 66622 24996
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 66314 23964 66622 23973
rect 66314 23962 66320 23964
rect 66376 23962 66400 23964
rect 66456 23962 66480 23964
rect 66536 23962 66560 23964
rect 66616 23962 66622 23964
rect 66376 23910 66378 23962
rect 66558 23910 66560 23962
rect 66314 23908 66320 23910
rect 66376 23908 66400 23910
rect 66456 23908 66480 23910
rect 66536 23908 66560 23910
rect 66616 23908 66622 23910
rect 66314 23899 66622 23908
rect 58532 23724 58584 23730
rect 58532 23666 58584 23672
rect 56048 23588 56100 23594
rect 56048 23530 56100 23536
rect 56060 22710 56088 23530
rect 58544 23322 58572 23666
rect 78220 23520 78272 23526
rect 78220 23462 78272 23468
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 58532 23316 58584 23322
rect 58532 23258 58584 23264
rect 56232 23180 56284 23186
rect 56232 23122 56284 23128
rect 56244 23050 56272 23122
rect 57060 23112 57112 23118
rect 57060 23054 57112 23060
rect 56232 23044 56284 23050
rect 56232 22986 56284 22992
rect 56876 23044 56928 23050
rect 56876 22986 56928 22992
rect 56048 22704 56100 22710
rect 56048 22646 56100 22652
rect 56244 22624 56272 22986
rect 56888 22778 56916 22986
rect 56876 22772 56928 22778
rect 56876 22714 56928 22720
rect 56324 22636 56376 22642
rect 56244 22596 56324 22624
rect 56244 21486 56272 22596
rect 56324 22578 56376 22584
rect 56968 22094 57020 22098
rect 57072 22094 57100 23054
rect 58544 22778 58572 23258
rect 78232 23225 78260 23462
rect 78218 23216 78274 23225
rect 78218 23151 78274 23160
rect 66314 22876 66622 22885
rect 66314 22874 66320 22876
rect 66376 22874 66400 22876
rect 66456 22874 66480 22876
rect 66536 22874 66560 22876
rect 66616 22874 66622 22876
rect 66376 22822 66378 22874
rect 66558 22822 66560 22874
rect 66314 22820 66320 22822
rect 66376 22820 66400 22822
rect 66456 22820 66480 22822
rect 66536 22820 66560 22822
rect 66616 22820 66622 22822
rect 66314 22811 66622 22820
rect 58532 22772 58584 22778
rect 58532 22714 58584 22720
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 56968 22092 57100 22094
rect 57020 22066 57100 22092
rect 56968 22034 57020 22040
rect 56980 21554 57008 22034
rect 66314 21788 66622 21797
rect 66314 21786 66320 21788
rect 66376 21786 66400 21788
rect 66456 21786 66480 21788
rect 66536 21786 66560 21788
rect 66616 21786 66622 21788
rect 66376 21734 66378 21786
rect 66558 21734 66560 21786
rect 66314 21732 66320 21734
rect 66376 21732 66400 21734
rect 66456 21732 66480 21734
rect 66536 21732 66560 21734
rect 66616 21732 66622 21734
rect 66314 21723 66622 21732
rect 56968 21548 57020 21554
rect 57020 21508 57100 21536
rect 56968 21490 57020 21496
rect 56232 21480 56284 21486
rect 56232 21422 56284 21428
rect 56600 21480 56652 21486
rect 56600 21422 56652 21428
rect 55956 20800 56008 20806
rect 55956 20742 56008 20748
rect 55968 20602 55996 20742
rect 56244 20618 56272 21422
rect 56612 21146 56640 21422
rect 56600 21140 56652 21146
rect 56600 21082 56652 21088
rect 55956 20596 56008 20602
rect 56244 20590 56364 20618
rect 55956 20538 56008 20544
rect 55496 20460 55548 20466
rect 55496 20402 55548 20408
rect 55404 20256 55456 20262
rect 55404 20198 55456 20204
rect 55416 19922 55444 20198
rect 55404 19916 55456 19922
rect 55404 19858 55456 19864
rect 55220 19780 55272 19786
rect 55220 19722 55272 19728
rect 55312 16788 55364 16794
rect 55312 16730 55364 16736
rect 55220 15360 55272 15366
rect 55220 15302 55272 15308
rect 55232 15094 55260 15302
rect 55220 15088 55272 15094
rect 55220 15030 55272 15036
rect 55324 12434 55352 16730
rect 55508 15502 55536 20402
rect 56336 20262 56364 20590
rect 56048 20256 56100 20262
rect 56048 20198 56100 20204
rect 56324 20256 56376 20262
rect 56324 20198 56376 20204
rect 56060 19446 56088 20198
rect 57072 19922 57100 21508
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 66314 20700 66622 20709
rect 66314 20698 66320 20700
rect 66376 20698 66400 20700
rect 66456 20698 66480 20700
rect 66536 20698 66560 20700
rect 66616 20698 66622 20700
rect 66376 20646 66378 20698
rect 66558 20646 66560 20698
rect 66314 20644 66320 20646
rect 66376 20644 66400 20646
rect 66456 20644 66480 20646
rect 66536 20644 66560 20646
rect 66616 20644 66622 20646
rect 66314 20635 66622 20644
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 57060 19916 57112 19922
rect 57060 19858 57112 19864
rect 66314 19612 66622 19621
rect 66314 19610 66320 19612
rect 66376 19610 66400 19612
rect 66456 19610 66480 19612
rect 66536 19610 66560 19612
rect 66616 19610 66622 19612
rect 66376 19558 66378 19610
rect 66558 19558 66560 19610
rect 66314 19556 66320 19558
rect 66376 19556 66400 19558
rect 66456 19556 66480 19558
rect 66536 19556 66560 19558
rect 66616 19556 66622 19558
rect 66314 19547 66622 19556
rect 56048 19440 56100 19446
rect 56048 19382 56100 19388
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 55864 18964 55916 18970
rect 55864 18906 55916 18912
rect 55876 18358 55904 18906
rect 56416 18828 56468 18834
rect 56416 18770 56468 18776
rect 56140 18624 56192 18630
rect 56140 18566 56192 18572
rect 56152 18358 56180 18566
rect 55864 18352 55916 18358
rect 55864 18294 55916 18300
rect 56140 18352 56192 18358
rect 56140 18294 56192 18300
rect 55772 16584 55824 16590
rect 55772 16526 55824 16532
rect 55680 16516 55732 16522
rect 55680 16458 55732 16464
rect 55692 16182 55720 16458
rect 55680 16176 55732 16182
rect 55680 16118 55732 16124
rect 55496 15496 55548 15502
rect 55496 15438 55548 15444
rect 55588 15088 55640 15094
rect 55692 15076 55720 16118
rect 55784 16017 55812 16526
rect 55770 16008 55826 16017
rect 55770 15943 55826 15952
rect 55772 15564 55824 15570
rect 55772 15506 55824 15512
rect 55640 15048 55720 15076
rect 55588 15030 55640 15036
rect 55600 13938 55628 15030
rect 55588 13932 55640 13938
rect 55588 13874 55640 13880
rect 55404 13728 55456 13734
rect 55404 13670 55456 13676
rect 55416 13394 55444 13670
rect 55404 13388 55456 13394
rect 55404 13330 55456 13336
rect 55232 12406 55352 12434
rect 55128 6452 55180 6458
rect 55128 6394 55180 6400
rect 55036 5772 55088 5778
rect 55036 5714 55088 5720
rect 54760 4684 54812 4690
rect 54760 4626 54812 4632
rect 55048 4622 55076 5714
rect 55140 5234 55168 6394
rect 55128 5228 55180 5234
rect 55128 5170 55180 5176
rect 53656 4616 53708 4622
rect 53656 4558 53708 4564
rect 55036 4616 55088 4622
rect 55036 4558 55088 4564
rect 54024 4140 54076 4146
rect 54024 4082 54076 4088
rect 52920 3528 52972 3534
rect 52920 3470 52972 3476
rect 54036 3126 54064 4082
rect 54300 3528 54352 3534
rect 54300 3470 54352 3476
rect 54312 3194 54340 3470
rect 54300 3188 54352 3194
rect 54300 3130 54352 3136
rect 54024 3120 54076 3126
rect 54024 3062 54076 3068
rect 51080 3052 51132 3058
rect 51080 2994 51132 3000
rect 51448 3052 51500 3058
rect 51448 2994 51500 3000
rect 51264 2848 51316 2854
rect 51264 2790 51316 2796
rect 51632 2848 51684 2854
rect 51632 2790 51684 2796
rect 53564 2848 53616 2854
rect 53564 2790 53616 2796
rect 54116 2848 54168 2854
rect 54116 2790 54168 2796
rect 50988 2644 51040 2650
rect 50988 2586 51040 2592
rect 51276 2446 51304 2790
rect 51644 2446 51672 2790
rect 53576 2446 53604 2790
rect 54128 2446 54156 2790
rect 54312 2650 54708 2666
rect 54312 2644 54720 2650
rect 54312 2638 54668 2644
rect 54312 2582 54340 2638
rect 54668 2586 54720 2592
rect 54300 2576 54352 2582
rect 54300 2518 54352 2524
rect 54484 2508 54536 2514
rect 54484 2450 54536 2456
rect 45192 2440 45244 2446
rect 45192 2382 45244 2388
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 46480 2440 46532 2446
rect 46480 2382 46532 2388
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 47768 2440 47820 2446
rect 47768 2382 47820 2388
rect 49056 2440 49108 2446
rect 49056 2382 49108 2388
rect 49792 2440 49844 2446
rect 49792 2382 49844 2388
rect 51264 2440 51316 2446
rect 51264 2382 51316 2388
rect 51632 2440 51684 2446
rect 51632 2382 51684 2388
rect 53564 2440 53616 2446
rect 53564 2382 53616 2388
rect 54116 2440 54168 2446
rect 54116 2382 54168 2388
rect 45204 2106 45232 2382
rect 50160 2372 50212 2378
rect 50160 2314 50212 2320
rect 50252 2372 50304 2378
rect 50252 2314 50304 2320
rect 45560 2304 45612 2310
rect 45560 2246 45612 2252
rect 45744 2304 45796 2310
rect 45744 2246 45796 2252
rect 46388 2304 46440 2310
rect 46388 2246 46440 2252
rect 46480 2304 46532 2310
rect 46480 2246 46532 2252
rect 47032 2304 47084 2310
rect 47032 2246 47084 2252
rect 47676 2304 47728 2310
rect 47676 2246 47728 2252
rect 48320 2304 48372 2310
rect 48320 2246 48372 2252
rect 48964 2304 49016 2310
rect 48964 2246 49016 2252
rect 49608 2304 49660 2310
rect 49608 2246 49660 2252
rect 45572 2106 45600 2246
rect 45192 2100 45244 2106
rect 45192 2042 45244 2048
rect 45560 2100 45612 2106
rect 45560 2042 45612 2048
rect 45756 800 45784 2246
rect 46400 2038 46428 2246
rect 46388 2032 46440 2038
rect 46388 1974 46440 1980
rect 46492 1170 46520 2246
rect 46400 1142 46520 1170
rect 46400 800 46428 1142
rect 47044 800 47072 2246
rect 47688 800 47716 2246
rect 48332 800 48360 2246
rect 48976 800 49004 2246
rect 49620 800 49648 2246
rect 50172 1970 50200 2314
rect 50160 1964 50212 1970
rect 50160 1906 50212 1912
rect 50172 1834 50200 1906
rect 50160 1828 50212 1834
rect 50160 1770 50212 1776
rect 50264 800 50292 2314
rect 50896 2304 50948 2310
rect 50896 2246 50948 2252
rect 51540 2304 51592 2310
rect 51540 2246 51592 2252
rect 52184 2304 52236 2310
rect 52184 2246 52236 2252
rect 52460 2304 52512 2310
rect 52460 2246 52512 2252
rect 52828 2304 52880 2310
rect 52828 2246 52880 2252
rect 53472 2304 53524 2310
rect 53472 2246 53524 2252
rect 50908 800 50936 2246
rect 51552 800 51580 2246
rect 52196 800 52224 2246
rect 52472 1902 52500 2246
rect 52460 1896 52512 1902
rect 52460 1838 52512 1844
rect 52840 800 52868 2246
rect 53484 800 53512 2246
rect 54128 800 54156 2382
rect 54496 1970 54524 2450
rect 54852 2440 54904 2446
rect 54852 2382 54904 2388
rect 54760 2304 54812 2310
rect 54760 2246 54812 2252
rect 54484 1964 54536 1970
rect 54484 1906 54536 1912
rect 54772 800 54800 2246
rect 54864 2106 54892 2382
rect 55036 2304 55088 2310
rect 55036 2246 55088 2252
rect 55048 2106 55076 2246
rect 54852 2100 54904 2106
rect 54852 2042 54904 2048
rect 55036 2100 55088 2106
rect 55036 2042 55088 2048
rect 55232 1834 55260 12406
rect 55404 12232 55456 12238
rect 55404 12174 55456 12180
rect 55312 9580 55364 9586
rect 55312 9522 55364 9528
rect 55324 9178 55352 9522
rect 55312 9172 55364 9178
rect 55312 9114 55364 9120
rect 55312 6112 55364 6118
rect 55312 6054 55364 6060
rect 55324 3670 55352 6054
rect 55416 5642 55444 12174
rect 55784 11354 55812 15506
rect 55876 12170 55904 18294
rect 56428 18290 56456 18770
rect 66314 18524 66622 18533
rect 66314 18522 66320 18524
rect 66376 18522 66400 18524
rect 66456 18522 66480 18524
rect 66536 18522 66560 18524
rect 66616 18522 66622 18524
rect 66376 18470 66378 18522
rect 66558 18470 66560 18522
rect 66314 18468 66320 18470
rect 66376 18468 66400 18470
rect 66456 18468 66480 18470
rect 66536 18468 66560 18470
rect 66616 18468 66622 18470
rect 66314 18459 66622 18468
rect 56416 18284 56468 18290
rect 56416 18226 56468 18232
rect 56428 16658 56456 18226
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 66314 17436 66622 17445
rect 66314 17434 66320 17436
rect 66376 17434 66400 17436
rect 66456 17434 66480 17436
rect 66536 17434 66560 17436
rect 66616 17434 66622 17436
rect 66376 17382 66378 17434
rect 66558 17382 66560 17434
rect 66314 17380 66320 17382
rect 66376 17380 66400 17382
rect 66456 17380 66480 17382
rect 66536 17380 66560 17382
rect 66616 17380 66622 17382
rect 66314 17371 66622 17380
rect 77852 17196 77904 17202
rect 77852 17138 77904 17144
rect 77864 16998 77892 17138
rect 78218 17096 78274 17105
rect 78218 17031 78220 17040
rect 78272 17031 78274 17040
rect 78220 17002 78272 17008
rect 77852 16992 77904 16998
rect 77852 16934 77904 16940
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 56416 16652 56468 16658
rect 56416 16594 56468 16600
rect 77864 16590 77892 16934
rect 56140 16584 56192 16590
rect 56140 16526 56192 16532
rect 77852 16584 77904 16590
rect 77852 16526 77904 16532
rect 56152 16250 56180 16526
rect 57980 16448 58032 16454
rect 57980 16390 58032 16396
rect 57992 16250 58020 16390
rect 66314 16348 66622 16357
rect 66314 16346 66320 16348
rect 66376 16346 66400 16348
rect 66456 16346 66480 16348
rect 66536 16346 66560 16348
rect 66616 16346 66622 16348
rect 66376 16294 66378 16346
rect 66558 16294 66560 16346
rect 66314 16292 66320 16294
rect 66376 16292 66400 16294
rect 66456 16292 66480 16294
rect 66536 16292 66560 16294
rect 66616 16292 66622 16294
rect 66314 16283 66622 16292
rect 56140 16244 56192 16250
rect 56140 16186 56192 16192
rect 57980 16244 58032 16250
rect 57980 16186 58032 16192
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 55956 15496 56008 15502
rect 55956 15438 56008 15444
rect 55968 15162 55996 15438
rect 56508 15428 56560 15434
rect 56508 15370 56560 15376
rect 56520 15162 56548 15370
rect 66314 15260 66622 15269
rect 66314 15258 66320 15260
rect 66376 15258 66400 15260
rect 66456 15258 66480 15260
rect 66536 15258 66560 15260
rect 66616 15258 66622 15260
rect 66376 15206 66378 15258
rect 66558 15206 66560 15258
rect 66314 15204 66320 15206
rect 66376 15204 66400 15206
rect 66456 15204 66480 15206
rect 66536 15204 66560 15206
rect 66616 15204 66622 15206
rect 66314 15195 66622 15204
rect 55956 15156 56008 15162
rect 55956 15098 56008 15104
rect 56508 15156 56560 15162
rect 56508 15098 56560 15104
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 66314 14172 66622 14181
rect 66314 14170 66320 14172
rect 66376 14170 66400 14172
rect 66456 14170 66480 14172
rect 66536 14170 66560 14172
rect 66616 14170 66622 14172
rect 66376 14118 66378 14170
rect 66558 14118 66560 14170
rect 66314 14116 66320 14118
rect 66376 14116 66400 14118
rect 66456 14116 66480 14118
rect 66536 14116 66560 14118
rect 66616 14116 66622 14118
rect 66314 14107 66622 14116
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 66314 13084 66622 13093
rect 66314 13082 66320 13084
rect 66376 13082 66400 13084
rect 66456 13082 66480 13084
rect 66536 13082 66560 13084
rect 66616 13082 66622 13084
rect 66376 13030 66378 13082
rect 66558 13030 66560 13082
rect 66314 13028 66320 13030
rect 66376 13028 66400 13030
rect 66456 13028 66480 13030
rect 66536 13028 66560 13030
rect 66616 13028 66622 13030
rect 66314 13019 66622 13028
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 55864 12164 55916 12170
rect 55864 12106 55916 12112
rect 66314 11996 66622 12005
rect 66314 11994 66320 11996
rect 66376 11994 66400 11996
rect 66456 11994 66480 11996
rect 66536 11994 66560 11996
rect 66616 11994 66622 11996
rect 66376 11942 66378 11994
rect 66558 11942 66560 11994
rect 66314 11940 66320 11942
rect 66376 11940 66400 11942
rect 66456 11940 66480 11942
rect 66536 11940 66560 11942
rect 66616 11940 66622 11942
rect 66314 11931 66622 11940
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 55772 11348 55824 11354
rect 55772 11290 55824 11296
rect 66314 10908 66622 10917
rect 66314 10906 66320 10908
rect 66376 10906 66400 10908
rect 66456 10906 66480 10908
rect 66536 10906 66560 10908
rect 66616 10906 66622 10908
rect 66376 10854 66378 10906
rect 66558 10854 66560 10906
rect 66314 10852 66320 10854
rect 66376 10852 66400 10854
rect 66456 10852 66480 10854
rect 66536 10852 66560 10854
rect 66616 10852 66622 10854
rect 66314 10843 66622 10852
rect 56600 10600 56652 10606
rect 56600 10542 56652 10548
rect 55772 10464 55824 10470
rect 55772 10406 55824 10412
rect 55588 9988 55640 9994
rect 55588 9930 55640 9936
rect 55600 9722 55628 9930
rect 55784 9926 55812 10406
rect 56612 10130 56640 10542
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 56600 10124 56652 10130
rect 56600 10066 56652 10072
rect 55772 9920 55824 9926
rect 55772 9862 55824 9868
rect 55588 9716 55640 9722
rect 55496 9686 55548 9692
rect 55588 9658 55640 9664
rect 55496 9628 55548 9634
rect 55508 9586 55536 9628
rect 55496 9580 55548 9586
rect 55496 9522 55548 9528
rect 55496 9376 55548 9382
rect 55494 9344 55496 9353
rect 55548 9344 55550 9353
rect 55494 9279 55550 9288
rect 55784 8022 55812 9862
rect 56612 9586 56640 10066
rect 66314 9820 66622 9829
rect 66314 9818 66320 9820
rect 66376 9818 66400 9820
rect 66456 9818 66480 9820
rect 66536 9818 66560 9820
rect 66616 9818 66622 9820
rect 66376 9766 66378 9818
rect 66558 9766 66560 9818
rect 66314 9764 66320 9766
rect 66376 9764 66400 9766
rect 66456 9764 66480 9766
rect 66536 9764 66560 9766
rect 66616 9764 66622 9766
rect 66314 9755 66622 9764
rect 56600 9580 56652 9586
rect 56600 9522 56652 9528
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 66314 8732 66622 8741
rect 66314 8730 66320 8732
rect 66376 8730 66400 8732
rect 66456 8730 66480 8732
rect 66536 8730 66560 8732
rect 66616 8730 66622 8732
rect 66376 8678 66378 8730
rect 66558 8678 66560 8730
rect 66314 8676 66320 8678
rect 66376 8676 66400 8678
rect 66456 8676 66480 8678
rect 66536 8676 66560 8678
rect 66616 8676 66622 8678
rect 66314 8667 66622 8676
rect 78036 8492 78088 8498
rect 78036 8434 78088 8440
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 78048 8090 78076 8434
rect 78220 8356 78272 8362
rect 78220 8298 78272 8304
rect 78232 8265 78260 8298
rect 78218 8256 78274 8265
rect 78218 8191 78274 8200
rect 78036 8084 78088 8090
rect 78036 8026 78088 8032
rect 55772 8016 55824 8022
rect 55772 7958 55824 7964
rect 55588 7812 55640 7818
rect 55588 7754 55640 7760
rect 55600 5778 55628 7754
rect 55784 7478 55812 7958
rect 77668 7744 77720 7750
rect 77668 7686 77720 7692
rect 78404 7744 78456 7750
rect 78404 7686 78456 7692
rect 66314 7644 66622 7653
rect 66314 7642 66320 7644
rect 66376 7642 66400 7644
rect 66456 7642 66480 7644
rect 66536 7642 66560 7644
rect 66616 7642 66622 7644
rect 66376 7590 66378 7642
rect 66558 7590 66560 7642
rect 66314 7588 66320 7590
rect 66376 7588 66400 7590
rect 66456 7588 66480 7590
rect 66536 7588 66560 7590
rect 66616 7588 66622 7590
rect 66314 7579 66622 7588
rect 55772 7472 55824 7478
rect 55772 7414 55824 7420
rect 55784 7206 55812 7414
rect 77680 7410 77708 7686
rect 78416 7585 78444 7686
rect 78402 7576 78458 7585
rect 78402 7511 78458 7520
rect 77668 7404 77720 7410
rect 77668 7346 77720 7352
rect 77680 7206 77708 7346
rect 55772 7200 55824 7206
rect 55772 7142 55824 7148
rect 77668 7200 77720 7206
rect 77668 7142 77720 7148
rect 78220 7200 78272 7206
rect 78220 7142 78272 7148
rect 55588 5772 55640 5778
rect 55588 5714 55640 5720
rect 55404 5636 55456 5642
rect 55404 5578 55456 5584
rect 55416 5098 55444 5578
rect 55784 5574 55812 7142
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 66314 6556 66622 6565
rect 66314 6554 66320 6556
rect 66376 6554 66400 6556
rect 66456 6554 66480 6556
rect 66536 6554 66560 6556
rect 66616 6554 66622 6556
rect 66376 6502 66378 6554
rect 66558 6502 66560 6554
rect 66314 6500 66320 6502
rect 66376 6500 66400 6502
rect 66456 6500 66480 6502
rect 66536 6500 66560 6502
rect 66616 6500 66622 6502
rect 66314 6491 66622 6500
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 77680 5574 77708 7142
rect 78232 6905 78260 7142
rect 78218 6896 78274 6905
rect 78218 6831 78274 6840
rect 77852 6792 77904 6798
rect 77852 6734 77904 6740
rect 55772 5568 55824 5574
rect 55772 5510 55824 5516
rect 77668 5568 77720 5574
rect 77668 5510 77720 5516
rect 66314 5468 66622 5477
rect 66314 5466 66320 5468
rect 66376 5466 66400 5468
rect 66456 5466 66480 5468
rect 66536 5466 66560 5468
rect 66616 5466 66622 5468
rect 66376 5414 66378 5466
rect 66558 5414 66560 5466
rect 66314 5412 66320 5414
rect 66376 5412 66400 5414
rect 66456 5412 66480 5414
rect 66536 5412 66560 5414
rect 66616 5412 66622 5414
rect 66314 5403 66622 5412
rect 56048 5160 56100 5166
rect 56048 5102 56100 5108
rect 55404 5092 55456 5098
rect 55404 5034 55456 5040
rect 55312 3664 55364 3670
rect 55312 3606 55364 3612
rect 55404 3596 55456 3602
rect 55404 3538 55456 3544
rect 55312 2848 55364 2854
rect 55312 2790 55364 2796
rect 55324 2446 55352 2790
rect 55312 2440 55364 2446
rect 55312 2382 55364 2388
rect 55220 1828 55272 1834
rect 55220 1770 55272 1776
rect 55416 800 55444 3538
rect 55496 3528 55548 3534
rect 55496 3470 55548 3476
rect 55508 3126 55536 3470
rect 55496 3120 55548 3126
rect 55496 3062 55548 3068
rect 55508 2582 55536 3062
rect 56060 2990 56088 5102
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 66314 4380 66622 4389
rect 66314 4378 66320 4380
rect 66376 4378 66400 4380
rect 66456 4378 66480 4380
rect 66536 4378 66560 4380
rect 66616 4378 66622 4380
rect 66376 4326 66378 4378
rect 66558 4326 66560 4378
rect 66314 4324 66320 4326
rect 66376 4324 66400 4326
rect 66456 4324 66480 4326
rect 66536 4324 66560 4326
rect 66616 4324 66622 4326
rect 66314 4315 66622 4324
rect 68192 4140 68244 4146
rect 68192 4082 68244 4088
rect 59360 4072 59412 4078
rect 59360 4014 59412 4020
rect 58992 4004 59044 4010
rect 58992 3946 59044 3952
rect 56416 3936 56468 3942
rect 56416 3878 56468 3884
rect 56428 3602 56456 3878
rect 57796 3664 57848 3670
rect 57796 3606 57848 3612
rect 56416 3596 56468 3602
rect 56416 3538 56468 3544
rect 57704 3596 57756 3602
rect 57704 3538 57756 3544
rect 56784 3392 56836 3398
rect 56784 3334 56836 3340
rect 56968 3392 57020 3398
rect 56968 3334 57020 3340
rect 56796 3126 56824 3334
rect 56784 3120 56836 3126
rect 56784 3062 56836 3068
rect 56324 3052 56376 3058
rect 56324 2994 56376 3000
rect 56048 2984 56100 2990
rect 56048 2926 56100 2932
rect 55496 2576 55548 2582
rect 55496 2518 55548 2524
rect 56060 2514 56088 2926
rect 56048 2508 56100 2514
rect 56048 2450 56100 2456
rect 56060 870 56180 898
rect 56060 800 56088 870
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56152 762 56180 870
rect 56336 762 56364 2994
rect 56600 2984 56652 2990
rect 56600 2926 56652 2932
rect 56612 2378 56640 2926
rect 56692 2508 56744 2514
rect 56692 2450 56744 2456
rect 56600 2372 56652 2378
rect 56600 2314 56652 2320
rect 56704 800 56732 2450
rect 56980 2310 57008 3334
rect 57428 2848 57480 2854
rect 57428 2790 57480 2796
rect 57336 2576 57388 2582
rect 57336 2518 57388 2524
rect 56968 2304 57020 2310
rect 56968 2246 57020 2252
rect 57348 800 57376 2518
rect 57440 2514 57468 2790
rect 57428 2508 57480 2514
rect 57428 2450 57480 2456
rect 57716 2310 57744 3538
rect 57808 3398 57836 3606
rect 59004 3534 59032 3946
rect 59372 3738 59400 4014
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 59360 3732 59412 3738
rect 59360 3674 59412 3680
rect 58164 3528 58216 3534
rect 58164 3470 58216 3476
rect 58992 3528 59044 3534
rect 58992 3470 59044 3476
rect 57796 3392 57848 3398
rect 57796 3334 57848 3340
rect 57808 3058 57836 3334
rect 57796 3052 57848 3058
rect 57796 2994 57848 3000
rect 57980 2848 58032 2854
rect 57980 2790 58032 2796
rect 57992 2650 58020 2790
rect 57980 2644 58032 2650
rect 57980 2586 58032 2592
rect 58176 2514 58204 3470
rect 58256 3460 58308 3466
rect 58256 3402 58308 3408
rect 58268 3194 58296 3402
rect 58440 3392 58492 3398
rect 58440 3334 58492 3340
rect 58256 3188 58308 3194
rect 58256 3130 58308 3136
rect 58452 2990 58480 3334
rect 66314 3292 66622 3301
rect 66314 3290 66320 3292
rect 66376 3290 66400 3292
rect 66456 3290 66480 3292
rect 66536 3290 66560 3292
rect 66616 3290 66622 3292
rect 66376 3238 66378 3290
rect 66558 3238 66560 3290
rect 66314 3236 66320 3238
rect 66376 3236 66400 3238
rect 66456 3236 66480 3238
rect 66536 3236 66560 3238
rect 66616 3236 66622 3238
rect 66314 3227 66622 3236
rect 66444 3120 66496 3126
rect 66444 3062 66496 3068
rect 58716 3052 58768 3058
rect 58716 2994 58768 3000
rect 59820 3052 59872 3058
rect 59820 2994 59872 3000
rect 58348 2984 58400 2990
rect 58348 2926 58400 2932
rect 58440 2984 58492 2990
rect 58440 2926 58492 2932
rect 58164 2508 58216 2514
rect 58164 2450 58216 2456
rect 57980 2440 58032 2446
rect 57980 2382 58032 2388
rect 57704 2304 57756 2310
rect 57704 2246 57756 2252
rect 57992 800 58020 2382
rect 58360 2310 58388 2926
rect 58728 2650 58756 2994
rect 58808 2984 58860 2990
rect 58808 2926 58860 2932
rect 59636 2984 59688 2990
rect 59636 2926 59688 2932
rect 59728 2984 59780 2990
rect 59728 2926 59780 2932
rect 58716 2644 58768 2650
rect 58716 2586 58768 2592
rect 58624 2372 58676 2378
rect 58624 2314 58676 2320
rect 58348 2304 58400 2310
rect 58348 2246 58400 2252
rect 58636 800 58664 2314
rect 58820 1902 58848 2926
rect 59648 2514 59676 2926
rect 59740 2582 59768 2926
rect 59832 2650 59860 2994
rect 60004 2984 60056 2990
rect 60004 2926 60056 2932
rect 59820 2644 59872 2650
rect 59820 2586 59872 2592
rect 59728 2576 59780 2582
rect 59728 2518 59780 2524
rect 59636 2508 59688 2514
rect 59636 2450 59688 2456
rect 59268 2304 59320 2310
rect 59268 2246 59320 2252
rect 59360 2304 59412 2310
rect 59360 2246 59412 2252
rect 59912 2304 59964 2310
rect 59912 2246 59964 2252
rect 58808 1896 58860 1902
rect 58808 1838 58860 1844
rect 59280 800 59308 2246
rect 59372 1970 59400 2246
rect 59360 1964 59412 1970
rect 59360 1906 59412 1912
rect 59924 800 59952 2246
rect 60016 2106 60044 2926
rect 66456 2854 66484 3062
rect 68204 3058 68232 4082
rect 72608 3732 72660 3738
rect 72608 3674 72660 3680
rect 68928 3664 68980 3670
rect 68928 3606 68980 3612
rect 68468 3528 68520 3534
rect 68468 3470 68520 3476
rect 68192 3052 68244 3058
rect 68192 2994 68244 3000
rect 66536 2984 66588 2990
rect 66536 2926 66588 2932
rect 61752 2848 61804 2854
rect 61752 2790 61804 2796
rect 62396 2848 62448 2854
rect 62396 2790 62448 2796
rect 63224 2848 63276 2854
rect 63224 2790 63276 2796
rect 63684 2848 63736 2854
rect 63684 2790 63736 2796
rect 64328 2848 64380 2854
rect 64328 2790 64380 2796
rect 65984 2848 66036 2854
rect 65984 2790 66036 2796
rect 66444 2848 66496 2854
rect 66444 2790 66496 2796
rect 61764 2446 61792 2790
rect 62408 2446 62436 2790
rect 63236 2446 63264 2790
rect 63696 2446 63724 2790
rect 64340 2446 64368 2790
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 61752 2440 61804 2446
rect 61752 2382 61804 2388
rect 62396 2440 62448 2446
rect 62396 2382 62448 2388
rect 63224 2440 63276 2446
rect 63224 2382 63276 2388
rect 63684 2440 63736 2446
rect 63684 2382 63736 2388
rect 64328 2440 64380 2446
rect 64328 2382 64380 2388
rect 60556 2304 60608 2310
rect 60556 2246 60608 2252
rect 61200 2304 61252 2310
rect 61200 2246 61252 2252
rect 61844 2304 61896 2310
rect 61844 2246 61896 2252
rect 62488 2304 62540 2310
rect 62488 2246 62540 2252
rect 63132 2304 63184 2310
rect 63132 2246 63184 2252
rect 63776 2304 63828 2310
rect 63776 2246 63828 2252
rect 64420 2304 64472 2310
rect 64420 2246 64472 2252
rect 65064 2304 65116 2310
rect 65064 2246 65116 2252
rect 65340 2304 65392 2310
rect 65340 2246 65392 2252
rect 65708 2304 65760 2310
rect 65708 2246 65760 2252
rect 60004 2100 60056 2106
rect 60004 2042 60056 2048
rect 60568 800 60596 2246
rect 61212 800 61240 2246
rect 61856 800 61884 2246
rect 62500 800 62528 2246
rect 63144 800 63172 2246
rect 63788 800 63816 2246
rect 64432 800 64460 2246
rect 65076 800 65104 2246
rect 65352 2106 65380 2246
rect 65340 2100 65392 2106
rect 65340 2042 65392 2048
rect 65720 800 65748 2246
rect 65996 2038 66024 2790
rect 66548 2650 66576 2926
rect 68480 2922 68508 3470
rect 68940 3194 68968 3606
rect 72424 3528 72476 3534
rect 72424 3470 72476 3476
rect 72148 3392 72200 3398
rect 72148 3334 72200 3340
rect 68928 3188 68980 3194
rect 68928 3130 68980 3136
rect 68940 3058 68968 3130
rect 72160 3126 72188 3334
rect 72436 3194 72464 3470
rect 72516 3460 72568 3466
rect 72516 3402 72568 3408
rect 72528 3194 72556 3402
rect 72620 3194 72648 3674
rect 77680 3670 77708 5510
rect 77668 3664 77720 3670
rect 77668 3606 77720 3612
rect 74448 3596 74500 3602
rect 74448 3538 74500 3544
rect 73528 3528 73580 3534
rect 73528 3470 73580 3476
rect 72884 3392 72936 3398
rect 73068 3392 73120 3398
rect 72884 3334 72936 3340
rect 72988 3340 73068 3346
rect 72988 3334 73120 3340
rect 72424 3188 72476 3194
rect 72424 3130 72476 3136
rect 72516 3188 72568 3194
rect 72516 3130 72568 3136
rect 72608 3188 72660 3194
rect 72608 3130 72660 3136
rect 72148 3120 72200 3126
rect 72148 3062 72200 3068
rect 68928 3052 68980 3058
rect 68928 2994 68980 3000
rect 69020 3052 69072 3058
rect 69020 2994 69072 3000
rect 71136 3052 71188 3058
rect 71136 2994 71188 3000
rect 71228 3052 71280 3058
rect 71228 2994 71280 3000
rect 72424 3052 72476 3058
rect 72424 2994 72476 3000
rect 68468 2916 68520 2922
rect 68468 2858 68520 2864
rect 67640 2848 67692 2854
rect 67640 2790 67692 2796
rect 68652 2848 68704 2854
rect 68652 2790 68704 2796
rect 67652 2650 67680 2790
rect 66536 2644 66588 2650
rect 66536 2586 66588 2592
rect 67640 2644 67692 2650
rect 67640 2586 67692 2592
rect 68664 2446 68692 2790
rect 69032 2582 69060 2994
rect 69756 2984 69808 2990
rect 69756 2926 69808 2932
rect 69768 2650 69796 2926
rect 71148 2650 71176 2994
rect 69756 2644 69808 2650
rect 69756 2586 69808 2592
rect 71136 2644 71188 2650
rect 71136 2586 71188 2592
rect 71240 2582 71268 2994
rect 72240 2984 72292 2990
rect 72240 2926 72292 2932
rect 72252 2650 72280 2926
rect 72240 2644 72292 2650
rect 72240 2586 72292 2592
rect 69020 2576 69072 2582
rect 71228 2576 71280 2582
rect 69020 2518 69072 2524
rect 71134 2544 71190 2553
rect 71228 2518 71280 2524
rect 71134 2479 71190 2488
rect 68652 2440 68704 2446
rect 68652 2382 68704 2388
rect 71148 2310 71176 2479
rect 72056 2440 72108 2446
rect 72108 2388 72280 2394
rect 72056 2382 72280 2388
rect 72068 2378 72280 2382
rect 72068 2372 72292 2378
rect 72068 2366 72240 2372
rect 66076 2304 66128 2310
rect 66260 2304 66312 2310
rect 66076 2246 66128 2252
rect 66180 2264 66260 2292
rect 65984 2032 66036 2038
rect 65984 1974 66036 1980
rect 66088 1970 66116 2246
rect 66180 1986 66208 2264
rect 66260 2246 66312 2252
rect 66996 2304 67048 2310
rect 66996 2246 67048 2252
rect 67640 2304 67692 2310
rect 67640 2246 67692 2252
rect 68284 2304 68336 2310
rect 68284 2246 68336 2252
rect 68928 2304 68980 2310
rect 68928 2246 68980 2252
rect 69572 2304 69624 2310
rect 69572 2246 69624 2252
rect 70216 2304 70268 2310
rect 70216 2246 70268 2252
rect 70860 2304 70912 2310
rect 70860 2246 70912 2252
rect 71136 2304 71188 2310
rect 71136 2246 71188 2252
rect 71504 2304 71556 2310
rect 71504 2246 71556 2252
rect 66314 2204 66622 2213
rect 66314 2202 66320 2204
rect 66376 2202 66400 2204
rect 66456 2202 66480 2204
rect 66536 2202 66560 2204
rect 66616 2202 66622 2204
rect 66376 2150 66378 2202
rect 66558 2150 66560 2202
rect 66314 2148 66320 2150
rect 66376 2148 66400 2150
rect 66456 2148 66480 2150
rect 66536 2148 66560 2150
rect 66616 2148 66622 2150
rect 66314 2139 66622 2148
rect 66076 1964 66128 1970
rect 66180 1958 66300 1986
rect 66076 1906 66128 1912
rect 66272 1578 66300 1958
rect 66272 1550 66392 1578
rect 66364 800 66392 1550
rect 67008 800 67036 2246
rect 67652 800 67680 2246
rect 68296 800 68324 2246
rect 68940 800 68968 2246
rect 69584 800 69612 2246
rect 70228 800 70256 2246
rect 70872 800 70900 2246
rect 71516 800 71544 2246
rect 72160 800 72188 2366
rect 72240 2314 72292 2320
rect 72436 2038 72464 2994
rect 72516 2984 72568 2990
rect 72516 2926 72568 2932
rect 72424 2032 72476 2038
rect 72424 1974 72476 1980
rect 72528 1970 72556 2926
rect 72896 2446 72924 3334
rect 72988 3318 73108 3334
rect 72988 2854 73016 3318
rect 73540 3194 73568 3470
rect 73528 3188 73580 3194
rect 73528 3130 73580 3136
rect 73988 3052 74040 3058
rect 73988 2994 74040 3000
rect 74172 3052 74224 3058
rect 74172 2994 74224 3000
rect 72976 2848 73028 2854
rect 72976 2790 73028 2796
rect 74000 2774 74028 2994
rect 74000 2746 74120 2774
rect 74092 2650 74120 2746
rect 74080 2644 74132 2650
rect 74080 2586 74132 2592
rect 74184 2553 74212 2994
rect 74460 2990 74488 3538
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 76208 3058 76236 3470
rect 77760 3392 77812 3398
rect 77760 3334 77812 3340
rect 77392 3120 77444 3126
rect 77392 3062 77444 3068
rect 76196 3052 76248 3058
rect 76196 2994 76248 3000
rect 74448 2984 74500 2990
rect 74448 2926 74500 2932
rect 74264 2916 74316 2922
rect 74264 2858 74316 2864
rect 74276 2650 74304 2858
rect 76104 2848 76156 2854
rect 76104 2790 76156 2796
rect 76748 2848 76800 2854
rect 76748 2790 76800 2796
rect 76116 2650 76144 2790
rect 74264 2644 74316 2650
rect 74264 2586 74316 2592
rect 76104 2644 76156 2650
rect 76104 2586 76156 2592
rect 74170 2544 74226 2553
rect 74170 2479 74226 2488
rect 76760 2446 76788 2790
rect 77404 2650 77432 3062
rect 77772 2650 77800 3334
rect 77864 3058 77892 6734
rect 78036 6656 78088 6662
rect 78036 6598 78088 6604
rect 78048 6322 78076 6598
rect 78036 6316 78088 6322
rect 78036 6258 78088 6264
rect 78218 6216 78274 6225
rect 78218 6151 78220 6160
rect 78272 6151 78274 6160
rect 78220 6122 78272 6128
rect 78404 5568 78456 5574
rect 78402 5536 78404 5545
rect 78456 5536 78458 5545
rect 78402 5471 78458 5480
rect 78312 5228 78364 5234
rect 78312 5170 78364 5176
rect 78128 5024 78180 5030
rect 78128 4966 78180 4972
rect 78140 3466 78168 4966
rect 78324 4865 78352 5170
rect 78310 4856 78366 4865
rect 78310 4791 78366 4800
rect 78496 4616 78548 4622
rect 78496 4558 78548 4564
rect 78312 4480 78364 4486
rect 78312 4422 78364 4428
rect 78324 4078 78352 4422
rect 78508 4185 78536 4558
rect 78494 4176 78550 4185
rect 78494 4111 78550 4120
rect 78312 4072 78364 4078
rect 78312 4014 78364 4020
rect 78128 3460 78180 3466
rect 78128 3402 78180 3408
rect 77944 3392 77996 3398
rect 77944 3334 77996 3340
rect 78496 3392 78548 3398
rect 78496 3334 78548 3340
rect 77852 3052 77904 3058
rect 77852 2994 77904 3000
rect 77392 2644 77444 2650
rect 77392 2586 77444 2592
rect 77760 2644 77812 2650
rect 77760 2586 77812 2592
rect 77956 2446 77984 3334
rect 78508 3058 78536 3334
rect 78496 3052 78548 3058
rect 78496 2994 78548 3000
rect 79232 3052 79284 3058
rect 79232 2994 79284 3000
rect 78036 2848 78088 2854
rect 78036 2790 78088 2796
rect 78048 2446 78076 2790
rect 72884 2440 72936 2446
rect 72884 2382 72936 2388
rect 76748 2440 76800 2446
rect 76748 2382 76800 2388
rect 77944 2440 77996 2446
rect 77944 2382 77996 2388
rect 78036 2440 78088 2446
rect 78036 2382 78088 2388
rect 73436 2372 73488 2378
rect 73436 2314 73488 2320
rect 72792 2304 72844 2310
rect 72792 2246 72844 2252
rect 72516 1964 72568 1970
rect 72516 1906 72568 1912
rect 72804 800 72832 2246
rect 73448 800 73476 2314
rect 74080 2304 74132 2310
rect 74080 2246 74132 2252
rect 74724 2304 74776 2310
rect 74724 2246 74776 2252
rect 75368 2304 75420 2310
rect 75368 2246 75420 2252
rect 76012 2304 76064 2310
rect 76012 2246 76064 2252
rect 76656 2304 76708 2310
rect 76656 2246 76708 2252
rect 77300 2304 77352 2310
rect 77300 2246 77352 2252
rect 74092 800 74120 2246
rect 74736 800 74764 2246
rect 75380 800 75408 2246
rect 76024 800 76052 2246
rect 76668 800 76696 2246
rect 77312 800 77340 2246
rect 77956 800 77984 2382
rect 78588 2304 78640 2310
rect 78588 2246 78640 2252
rect 78600 800 78628 2246
rect 79244 800 79272 2994
rect 56152 734 56364 762
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 79874 0 79930 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 1306 36760 1362 36816
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 938 36080 994 36136
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 938 35436 940 35456
rect 940 35436 992 35456
rect 992 35436 994 35456
rect 938 35400 994 35436
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 1306 34740 1362 34776
rect 1306 34720 1308 34740
rect 1308 34720 1360 34740
rect 1360 34720 1362 34740
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 938 34076 940 34096
rect 940 34076 992 34096
rect 992 34076 994 34096
rect 938 34040 994 34076
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 938 33380 994 33416
rect 938 33360 940 33380
rect 940 33360 992 33380
rect 992 33360 994 33380
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 938 32716 940 32736
rect 940 32716 992 32736
rect 992 32716 994 32736
rect 938 32680 994 32716
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 1306 32020 1362 32056
rect 1306 32000 1308 32020
rect 1308 32000 1360 32020
rect 1360 32000 1362 32020
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 938 31320 994 31376
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 938 30640 994 30696
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 938 29996 940 30016
rect 940 29996 992 30016
rect 992 29996 994 30016
rect 938 29960 994 29996
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 1306 29300 1362 29336
rect 1306 29280 1308 29300
rect 1308 29280 1360 29300
rect 1360 29280 1362 29300
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 938 28636 940 28656
rect 940 28636 992 28656
rect 992 28636 994 28656
rect 938 28600 994 28636
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 938 27940 994 27976
rect 938 27920 940 27940
rect 940 27920 992 27940
rect 992 27920 994 27940
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 938 27276 940 27296
rect 940 27276 992 27296
rect 992 27276 994 27296
rect 938 27240 994 27276
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 1306 26580 1362 26616
rect 1306 26560 1308 26580
rect 1308 26560 1360 26580
rect 1360 26560 1362 26580
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 12530 30096 12586 30152
rect 14554 30132 14556 30152
rect 14556 30132 14608 30152
rect 14608 30132 14610 30152
rect 14554 30096 14610 30132
rect 938 25880 994 25936
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 938 25200 994 25256
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 938 24556 940 24576
rect 940 24556 992 24576
rect 992 24556 994 24576
rect 938 24520 994 24556
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 1306 23860 1362 23896
rect 1306 23840 1308 23860
rect 1308 23840 1360 23860
rect 1360 23840 1362 23860
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 1214 23196 1216 23216
rect 1216 23196 1268 23216
rect 1268 23196 1270 23216
rect 1214 23160 1270 23196
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 938 22616 994 22672
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 846 21936 902 21992
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 846 21292 848 21312
rect 848 21292 900 21312
rect 900 21292 902 21312
rect 846 21256 902 21292
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 1490 20440 1546 20496
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 846 19660 848 19680
rect 848 19660 900 19680
rect 900 19660 902 19680
rect 846 19624 902 19660
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 29826 23060 29828 23080
rect 29828 23060 29880 23080
rect 29880 23060 29882 23080
rect 29826 23024 29882 23060
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1306 15680 1362 15736
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 1398 15000 1454 15056
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1214 14356 1216 14376
rect 1216 14356 1268 14376
rect 1268 14356 1270 14376
rect 1214 14320 1270 14356
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 1398 13640 1454 13696
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19798 15680 19854 15736
rect 21086 15544 21142 15600
rect 21270 15408 21326 15464
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 22558 14048 22614 14104
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 23754 16396 23756 16416
rect 23756 16396 23808 16416
rect 23808 16396 23810 16416
rect 23754 16360 23810 16396
rect 24214 15408 24270 15464
rect 24766 14340 24822 14376
rect 24766 14320 24768 14340
rect 24768 14320 24820 14340
rect 24820 14320 24822 14340
rect 24858 13932 24914 13968
rect 24858 13912 24860 13932
rect 24860 13912 24912 13932
rect 24912 13912 24914 13932
rect 25226 15544 25282 15600
rect 25134 15408 25190 15464
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 25594 13776 25650 13832
rect 26422 13812 26424 13832
rect 26424 13812 26476 13832
rect 26476 13812 26478 13832
rect 26422 13776 26478 13812
rect 26698 16360 26754 16416
rect 27342 16360 27398 16416
rect 27526 14356 27528 14376
rect 27528 14356 27580 14376
rect 27580 14356 27582 14376
rect 27526 14320 27582 14356
rect 29458 18164 29460 18184
rect 29460 18164 29512 18184
rect 29512 18164 29514 18184
rect 29458 18128 29514 18164
rect 27710 15680 27766 15736
rect 27618 14048 27674 14104
rect 27342 13932 27398 13968
rect 27342 13912 27344 13932
rect 27344 13912 27396 13932
rect 27396 13912 27398 13932
rect 28170 14864 28226 14920
rect 28630 14320 28686 14376
rect 29826 20440 29882 20496
rect 32586 25356 32642 25392
rect 32586 25336 32588 25356
rect 32588 25336 32640 25356
rect 32640 25336 32642 25356
rect 31758 23044 31814 23080
rect 31758 23024 31760 23044
rect 31760 23024 31812 23044
rect 31812 23024 31814 23044
rect 30194 17212 30196 17232
rect 30196 17212 30248 17232
rect 30248 17212 30250 17232
rect 30194 17176 30250 17212
rect 27986 9460 27988 9480
rect 27988 9460 28040 9480
rect 28040 9460 28042 9480
rect 27986 9424 28042 9460
rect 28262 9424 28318 9480
rect 29826 8880 29882 8936
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 31758 19216 31814 19272
rect 31390 17584 31446 17640
rect 31758 17040 31814 17096
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34886 25336 34942 25392
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 34058 20304 34114 20360
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 32954 17040 33010 17096
rect 31206 11092 31208 11112
rect 31208 11092 31260 11112
rect 31260 11092 31262 11112
rect 31206 11056 31262 11092
rect 31574 9560 31630 9616
rect 31666 9288 31722 9344
rect 32402 13932 32458 13968
rect 32402 13912 32404 13932
rect 32404 13912 32456 13932
rect 32456 13912 32458 13932
rect 33138 15020 33194 15056
rect 33138 15000 33140 15020
rect 33140 15000 33192 15020
rect 33192 15000 33194 15020
rect 33598 17196 33654 17232
rect 33598 17176 33600 17196
rect 33600 17176 33652 17196
rect 33652 17176 33654 17196
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 36174 22924 36176 22944
rect 36176 22924 36228 22944
rect 36228 22924 36230 22944
rect 36174 22888 36230 22924
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 33414 13912 33470 13968
rect 34058 13932 34114 13968
rect 34058 13912 34060 13932
rect 34060 13912 34112 13932
rect 34112 13912 34114 13932
rect 32218 9016 32274 9072
rect 33230 9424 33286 9480
rect 32770 9288 32826 9344
rect 33322 9288 33378 9344
rect 33782 9288 33838 9344
rect 33414 8472 33470 8528
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 36726 19372 36782 19408
rect 36910 19660 36912 19680
rect 36912 19660 36964 19680
rect 36964 19660 36966 19680
rect 36910 19624 36966 19660
rect 36726 19352 36728 19372
rect 36728 19352 36780 19372
rect 36780 19352 36782 19372
rect 37370 19080 37426 19136
rect 37646 19352 37702 19408
rect 38382 22616 38438 22672
rect 38382 22480 38438 22536
rect 38290 19508 38346 19544
rect 38934 22344 38990 22400
rect 38290 19488 38292 19508
rect 38292 19488 38344 19508
rect 38344 19488 38346 19508
rect 36634 14356 36636 14376
rect 36636 14356 36688 14376
rect 36688 14356 36690 14376
rect 36634 14320 36690 14356
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34334 9580 34390 9616
rect 34334 9560 34336 9580
rect 34336 9560 34388 9580
rect 34388 9560 34390 9580
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 35714 9596 35716 9616
rect 35716 9596 35768 9616
rect 35768 9596 35770 9616
rect 35714 9560 35770 9596
rect 34518 9288 34574 9344
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34610 9016 34666 9072
rect 35990 9424 36046 9480
rect 35898 9324 35900 9344
rect 35900 9324 35952 9344
rect 35952 9324 35954 9344
rect 35898 9288 35954 9324
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35530 8472 35586 8528
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 36910 14320 36966 14376
rect 36358 9288 36414 9344
rect 36358 8608 36414 8664
rect 36082 8336 36138 8392
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 36726 8608 36782 8664
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 37462 12860 37464 12880
rect 37464 12860 37516 12880
rect 37516 12860 37518 12880
rect 37462 12824 37518 12860
rect 38198 17604 38254 17640
rect 38198 17584 38200 17604
rect 38200 17584 38252 17604
rect 38252 17584 38254 17604
rect 38382 18028 38384 18048
rect 38384 18028 38436 18048
rect 38436 18028 38438 18048
rect 38382 17992 38438 18028
rect 38290 12844 38346 12880
rect 38290 12824 38292 12844
rect 38292 12824 38344 12844
rect 38344 12824 38346 12844
rect 37554 9560 37610 9616
rect 39210 22344 39266 22400
rect 40406 24012 40408 24032
rect 40408 24012 40460 24032
rect 40460 24012 40462 24032
rect 40406 23976 40462 24012
rect 40222 22380 40224 22400
rect 40224 22380 40276 22400
rect 40276 22380 40278 22400
rect 40222 22344 40278 22380
rect 39302 20304 39358 20360
rect 39854 18944 39910 19000
rect 39486 17040 39542 17096
rect 39394 15136 39450 15192
rect 40314 19372 40370 19408
rect 40314 19352 40316 19372
rect 40316 19352 40368 19372
rect 40368 19352 40370 19372
rect 40038 17720 40094 17776
rect 40406 19080 40462 19136
rect 41878 22208 41934 22264
rect 40590 19352 40646 19408
rect 40774 19372 40830 19408
rect 40774 19352 40776 19372
rect 40776 19352 40828 19372
rect 40828 19352 40830 19372
rect 41786 19488 41842 19544
rect 41050 19352 41106 19408
rect 41050 19216 41106 19272
rect 41418 17060 41474 17096
rect 41418 17040 41420 17060
rect 41420 17040 41472 17060
rect 41472 17040 41474 17060
rect 41418 15136 41474 15192
rect 41050 15020 41106 15056
rect 41050 15000 41052 15020
rect 41052 15000 41104 15020
rect 41104 15000 41106 15020
rect 40590 13932 40646 13968
rect 40590 13912 40592 13932
rect 40592 13912 40644 13932
rect 40644 13912 40646 13932
rect 39670 10920 39726 10976
rect 40774 13404 40776 13424
rect 40776 13404 40828 13424
rect 40828 13404 40830 13424
rect 40774 13368 40830 13404
rect 37830 6840 37886 6896
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 42614 24928 42670 24984
rect 42890 22888 42946 22944
rect 40774 8336 40830 8392
rect 40498 6976 40554 7032
rect 41050 6704 41106 6760
rect 41326 6976 41382 7032
rect 41510 6704 41566 6760
rect 43166 22516 43168 22536
rect 43168 22516 43220 22536
rect 43220 22516 43222 22536
rect 43166 22480 43222 22516
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 66320 37018 66376 37020
rect 66400 37018 66456 37020
rect 66480 37018 66536 37020
rect 66560 37018 66616 37020
rect 66320 36966 66366 37018
rect 66366 36966 66376 37018
rect 66400 36966 66430 37018
rect 66430 36966 66442 37018
rect 66442 36966 66456 37018
rect 66480 36966 66494 37018
rect 66494 36966 66506 37018
rect 66506 36966 66536 37018
rect 66560 36966 66570 37018
rect 66570 36966 66616 37018
rect 66320 36964 66376 36966
rect 66400 36964 66456 36966
rect 66480 36964 66536 36966
rect 66560 36964 66616 36966
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 66320 35930 66376 35932
rect 66400 35930 66456 35932
rect 66480 35930 66536 35932
rect 66560 35930 66616 35932
rect 66320 35878 66366 35930
rect 66366 35878 66376 35930
rect 66400 35878 66430 35930
rect 66430 35878 66442 35930
rect 66442 35878 66456 35930
rect 66480 35878 66494 35930
rect 66494 35878 66506 35930
rect 66506 35878 66536 35930
rect 66560 35878 66570 35930
rect 66570 35878 66616 35930
rect 66320 35876 66376 35878
rect 66400 35876 66456 35878
rect 66480 35876 66536 35878
rect 66560 35876 66616 35878
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 66320 34842 66376 34844
rect 66400 34842 66456 34844
rect 66480 34842 66536 34844
rect 66560 34842 66616 34844
rect 66320 34790 66366 34842
rect 66366 34790 66376 34842
rect 66400 34790 66430 34842
rect 66430 34790 66442 34842
rect 66442 34790 66456 34842
rect 66480 34790 66494 34842
rect 66494 34790 66506 34842
rect 66506 34790 66536 34842
rect 66560 34790 66570 34842
rect 66570 34790 66616 34842
rect 66320 34788 66376 34790
rect 66400 34788 66456 34790
rect 66480 34788 66536 34790
rect 66560 34788 66616 34790
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 66320 33754 66376 33756
rect 66400 33754 66456 33756
rect 66480 33754 66536 33756
rect 66560 33754 66616 33756
rect 66320 33702 66366 33754
rect 66366 33702 66376 33754
rect 66400 33702 66430 33754
rect 66430 33702 66442 33754
rect 66442 33702 66456 33754
rect 66480 33702 66494 33754
rect 66494 33702 66506 33754
rect 66506 33702 66536 33754
rect 66560 33702 66570 33754
rect 66570 33702 66616 33754
rect 66320 33700 66376 33702
rect 66400 33700 66456 33702
rect 66480 33700 66536 33702
rect 66560 33700 66616 33702
rect 44822 29996 44824 30016
rect 44824 29996 44876 30016
rect 44876 29996 44878 30016
rect 44822 29960 44878 29996
rect 44270 24928 44326 24984
rect 43534 23976 43590 24032
rect 44270 23024 44326 23080
rect 43994 22108 43996 22128
rect 43996 22108 44048 22128
rect 44048 22108 44050 22128
rect 43994 22072 44050 22108
rect 42338 8492 42394 8528
rect 42338 8472 42340 8492
rect 42340 8472 42392 8492
rect 42392 8472 42394 8492
rect 43166 17620 43168 17640
rect 43168 17620 43220 17640
rect 43220 17620 43222 17640
rect 43166 17584 43222 17620
rect 42982 14728 43038 14784
rect 42890 9288 42946 9344
rect 42890 8492 42946 8528
rect 42890 8472 42892 8492
rect 42892 8472 42944 8492
rect 42944 8472 42946 8492
rect 43534 17176 43590 17232
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 66320 32666 66376 32668
rect 66400 32666 66456 32668
rect 66480 32666 66536 32668
rect 66560 32666 66616 32668
rect 66320 32614 66366 32666
rect 66366 32614 66376 32666
rect 66400 32614 66430 32666
rect 66430 32614 66442 32666
rect 66442 32614 66456 32666
rect 66480 32614 66494 32666
rect 66494 32614 66506 32666
rect 66506 32614 66536 32666
rect 66560 32614 66570 32666
rect 66570 32614 66616 32666
rect 66320 32612 66376 32614
rect 66400 32612 66456 32614
rect 66480 32612 66536 32614
rect 66560 32612 66616 32614
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 66320 31578 66376 31580
rect 66400 31578 66456 31580
rect 66480 31578 66536 31580
rect 66560 31578 66616 31580
rect 66320 31526 66366 31578
rect 66366 31526 66376 31578
rect 66400 31526 66430 31578
rect 66430 31526 66442 31578
rect 66442 31526 66456 31578
rect 66480 31526 66494 31578
rect 66494 31526 66506 31578
rect 66506 31526 66536 31578
rect 66560 31526 66570 31578
rect 66570 31526 66616 31578
rect 66320 31524 66376 31526
rect 66400 31524 66456 31526
rect 66480 31524 66536 31526
rect 66560 31524 66616 31526
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 66320 30490 66376 30492
rect 66400 30490 66456 30492
rect 66480 30490 66536 30492
rect 66560 30490 66616 30492
rect 66320 30438 66366 30490
rect 66366 30438 66376 30490
rect 66400 30438 66430 30490
rect 66430 30438 66442 30490
rect 66442 30438 66456 30490
rect 66480 30438 66494 30490
rect 66494 30438 66506 30490
rect 66506 30438 66536 30490
rect 66560 30438 66570 30490
rect 66570 30438 66616 30490
rect 66320 30436 66376 30438
rect 66400 30436 66456 30438
rect 66480 30436 66536 30438
rect 66560 30436 66616 30438
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 66320 29402 66376 29404
rect 66400 29402 66456 29404
rect 66480 29402 66536 29404
rect 66560 29402 66616 29404
rect 66320 29350 66366 29402
rect 66366 29350 66376 29402
rect 66400 29350 66430 29402
rect 66430 29350 66442 29402
rect 66442 29350 66456 29402
rect 66480 29350 66494 29402
rect 66494 29350 66506 29402
rect 66506 29350 66536 29402
rect 66560 29350 66570 29402
rect 66570 29350 66616 29402
rect 66320 29348 66376 29350
rect 66400 29348 66456 29350
rect 66480 29348 66536 29350
rect 66560 29348 66616 29350
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 45834 23976 45890 24032
rect 44454 22344 44510 22400
rect 44362 20032 44418 20088
rect 43810 14728 43866 14784
rect 45374 23060 45376 23080
rect 45376 23060 45428 23080
rect 45428 23060 45430 23080
rect 45374 23024 45430 23060
rect 45098 22924 45100 22944
rect 45100 22924 45152 22944
rect 45152 22924 45154 22944
rect 45098 22888 45154 22924
rect 44730 19624 44786 19680
rect 44546 17740 44602 17776
rect 44546 17720 44548 17740
rect 44548 17720 44600 17740
rect 44600 17720 44602 17740
rect 44454 16088 44510 16144
rect 43626 8880 43682 8936
rect 43718 8200 43774 8256
rect 43718 6976 43774 7032
rect 44086 8916 44088 8936
rect 44088 8916 44140 8936
rect 44140 8916 44142 8936
rect 44086 8880 44142 8916
rect 46754 22108 46756 22128
rect 46756 22108 46808 22128
rect 46808 22108 46810 22128
rect 46754 22072 46810 22108
rect 46202 19080 46258 19136
rect 45926 17604 45982 17640
rect 45926 17584 45928 17604
rect 45928 17584 45980 17604
rect 45980 17584 45982 17604
rect 45190 14340 45246 14376
rect 45190 14320 45192 14340
rect 45192 14320 45244 14340
rect 45244 14320 45246 14340
rect 45466 14864 45522 14920
rect 47214 20576 47270 20632
rect 47398 22616 47454 22672
rect 48042 20576 48098 20632
rect 48410 21004 48466 21040
rect 48410 20984 48412 21004
rect 48412 20984 48464 21004
rect 48464 20984 48466 21004
rect 48870 22480 48926 22536
rect 48594 20440 48650 20496
rect 48042 18944 48098 19000
rect 45834 15428 45890 15464
rect 45834 15408 45836 15428
rect 45836 15408 45888 15428
rect 45888 15408 45890 15428
rect 46662 14184 46718 14240
rect 45650 13368 45706 13424
rect 49698 22924 49700 22944
rect 49700 22924 49752 22944
rect 49752 22924 49754 22944
rect 49698 22888 49754 22924
rect 49054 18128 49110 18184
rect 48226 14320 48282 14376
rect 44730 9016 44786 9072
rect 44914 8336 44970 8392
rect 45282 8236 45284 8256
rect 45284 8236 45336 8256
rect 45336 8236 45338 8256
rect 45282 8200 45338 8236
rect 49514 16108 49570 16144
rect 49514 16088 49516 16108
rect 49516 16088 49568 16108
rect 49568 16088 49570 16108
rect 45006 6860 45062 6896
rect 45006 6840 45008 6860
rect 45008 6840 45060 6860
rect 45060 6840 45062 6860
rect 48594 11092 48596 11112
rect 48596 11092 48648 11112
rect 48648 11092 48650 11112
rect 48594 11056 48650 11092
rect 49698 21256 49754 21312
rect 49698 16360 49754 16416
rect 49514 14764 49516 14784
rect 49516 14764 49568 14784
rect 49568 14764 49570 14784
rect 49514 14728 49570 14764
rect 49698 9288 49754 9344
rect 49698 9036 49754 9072
rect 49698 9016 49700 9036
rect 49700 9016 49752 9036
rect 49752 9016 49754 9036
rect 49698 8900 49754 8936
rect 49698 8880 49700 8900
rect 49700 8880 49752 8900
rect 49752 8880 49754 8900
rect 50710 22208 50766 22264
rect 50526 21256 50582 21312
rect 50250 16360 50306 16416
rect 50434 16224 50490 16280
rect 50434 15972 50490 16008
rect 50434 15952 50436 15972
rect 50436 15952 50488 15972
rect 50488 15952 50490 15972
rect 50434 14492 50436 14512
rect 50436 14492 50488 14512
rect 50488 14492 50490 14512
rect 50434 14456 50490 14492
rect 50342 14184 50398 14240
rect 50158 9152 50214 9208
rect 50158 8472 50214 8528
rect 50342 9580 50398 9616
rect 50342 9560 50344 9580
rect 50344 9560 50396 9580
rect 50396 9560 50398 9580
rect 51814 25644 51816 25664
rect 51816 25644 51868 25664
rect 51868 25644 51870 25664
rect 51814 25608 51870 25644
rect 50894 21020 50896 21040
rect 50896 21020 50948 21040
rect 50948 21020 50950 21040
rect 50894 20984 50950 21020
rect 50802 20848 50858 20904
rect 51170 20848 51226 20904
rect 50894 16396 50896 16416
rect 50896 16396 50948 16416
rect 50948 16396 50950 16416
rect 50894 16360 50950 16396
rect 50894 16108 50950 16144
rect 50894 16088 50896 16108
rect 50896 16088 50948 16108
rect 50948 16088 50950 16108
rect 51262 16360 51318 16416
rect 51262 14220 51264 14240
rect 51264 14220 51316 14240
rect 51316 14220 51318 14240
rect 51262 14184 51318 14220
rect 50986 14048 51042 14104
rect 53378 21956 53434 21992
rect 53378 21936 53380 21956
rect 53380 21936 53432 21956
rect 53432 21936 53434 21956
rect 51630 16088 51686 16144
rect 53194 17620 53196 17640
rect 53196 17620 53248 17640
rect 53248 17620 53250 17640
rect 53194 17584 53250 17620
rect 55126 20032 55182 20088
rect 54114 17620 54116 17640
rect 54116 17620 54168 17640
rect 54168 17620 54170 17640
rect 54114 17584 54170 17620
rect 53746 16224 53802 16280
rect 53378 15408 53434 15464
rect 53010 14320 53066 14376
rect 51906 14048 51962 14104
rect 50986 8900 51042 8936
rect 50986 8880 50988 8900
rect 50988 8880 51040 8900
rect 51040 8880 51042 8900
rect 51630 9596 51632 9616
rect 51632 9596 51684 9616
rect 51684 9596 51686 9616
rect 51630 9560 51686 9596
rect 54758 14356 54760 14376
rect 54760 14356 54812 14376
rect 54812 14356 54814 14376
rect 53194 9324 53196 9344
rect 53196 9324 53248 9344
rect 53248 9324 53250 9344
rect 53194 9288 53250 9324
rect 54758 14320 54814 14356
rect 54482 9424 54538 9480
rect 55034 9424 55090 9480
rect 66320 28314 66376 28316
rect 66400 28314 66456 28316
rect 66480 28314 66536 28316
rect 66560 28314 66616 28316
rect 66320 28262 66366 28314
rect 66366 28262 66376 28314
rect 66400 28262 66430 28314
rect 66430 28262 66442 28314
rect 66442 28262 66456 28314
rect 66480 28262 66494 28314
rect 66494 28262 66506 28314
rect 66506 28262 66536 28314
rect 66560 28262 66570 28314
rect 66570 28262 66616 28314
rect 66320 28260 66376 28262
rect 66400 28260 66456 28262
rect 66480 28260 66536 28262
rect 66560 28260 66616 28262
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 66320 27226 66376 27228
rect 66400 27226 66456 27228
rect 66480 27226 66536 27228
rect 66560 27226 66616 27228
rect 66320 27174 66366 27226
rect 66366 27174 66376 27226
rect 66400 27174 66430 27226
rect 66430 27174 66442 27226
rect 66442 27174 66456 27226
rect 66480 27174 66494 27226
rect 66494 27174 66506 27226
rect 66506 27174 66536 27226
rect 66560 27174 66570 27226
rect 66570 27174 66616 27226
rect 66320 27172 66376 27174
rect 66400 27172 66456 27174
rect 66480 27172 66536 27174
rect 66560 27172 66616 27174
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 66320 26138 66376 26140
rect 66400 26138 66456 26140
rect 66480 26138 66536 26140
rect 66560 26138 66616 26140
rect 66320 26086 66366 26138
rect 66366 26086 66376 26138
rect 66400 26086 66430 26138
rect 66430 26086 66442 26138
rect 66442 26086 66456 26138
rect 66480 26086 66494 26138
rect 66494 26086 66506 26138
rect 66506 26086 66536 26138
rect 66560 26086 66570 26138
rect 66570 26086 66616 26138
rect 66320 26084 66376 26086
rect 66400 26084 66456 26086
rect 66480 26084 66536 26086
rect 66560 26084 66616 26086
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 66320 25050 66376 25052
rect 66400 25050 66456 25052
rect 66480 25050 66536 25052
rect 66560 25050 66616 25052
rect 66320 24998 66366 25050
rect 66366 24998 66376 25050
rect 66400 24998 66430 25050
rect 66430 24998 66442 25050
rect 66442 24998 66456 25050
rect 66480 24998 66494 25050
rect 66494 24998 66506 25050
rect 66506 24998 66536 25050
rect 66560 24998 66570 25050
rect 66570 24998 66616 25050
rect 66320 24996 66376 24998
rect 66400 24996 66456 24998
rect 66480 24996 66536 24998
rect 66560 24996 66616 24998
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 66320 23962 66376 23964
rect 66400 23962 66456 23964
rect 66480 23962 66536 23964
rect 66560 23962 66616 23964
rect 66320 23910 66366 23962
rect 66366 23910 66376 23962
rect 66400 23910 66430 23962
rect 66430 23910 66442 23962
rect 66442 23910 66456 23962
rect 66480 23910 66494 23962
rect 66494 23910 66506 23962
rect 66506 23910 66536 23962
rect 66560 23910 66570 23962
rect 66570 23910 66616 23962
rect 66320 23908 66376 23910
rect 66400 23908 66456 23910
rect 66480 23908 66536 23910
rect 66560 23908 66616 23910
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 78218 23160 78274 23216
rect 66320 22874 66376 22876
rect 66400 22874 66456 22876
rect 66480 22874 66536 22876
rect 66560 22874 66616 22876
rect 66320 22822 66366 22874
rect 66366 22822 66376 22874
rect 66400 22822 66430 22874
rect 66430 22822 66442 22874
rect 66442 22822 66456 22874
rect 66480 22822 66494 22874
rect 66494 22822 66506 22874
rect 66506 22822 66536 22874
rect 66560 22822 66570 22874
rect 66570 22822 66616 22874
rect 66320 22820 66376 22822
rect 66400 22820 66456 22822
rect 66480 22820 66536 22822
rect 66560 22820 66616 22822
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 66320 21786 66376 21788
rect 66400 21786 66456 21788
rect 66480 21786 66536 21788
rect 66560 21786 66616 21788
rect 66320 21734 66366 21786
rect 66366 21734 66376 21786
rect 66400 21734 66430 21786
rect 66430 21734 66442 21786
rect 66442 21734 66456 21786
rect 66480 21734 66494 21786
rect 66494 21734 66506 21786
rect 66506 21734 66536 21786
rect 66560 21734 66570 21786
rect 66570 21734 66616 21786
rect 66320 21732 66376 21734
rect 66400 21732 66456 21734
rect 66480 21732 66536 21734
rect 66560 21732 66616 21734
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 66320 20698 66376 20700
rect 66400 20698 66456 20700
rect 66480 20698 66536 20700
rect 66560 20698 66616 20700
rect 66320 20646 66366 20698
rect 66366 20646 66376 20698
rect 66400 20646 66430 20698
rect 66430 20646 66442 20698
rect 66442 20646 66456 20698
rect 66480 20646 66494 20698
rect 66494 20646 66506 20698
rect 66506 20646 66536 20698
rect 66560 20646 66570 20698
rect 66570 20646 66616 20698
rect 66320 20644 66376 20646
rect 66400 20644 66456 20646
rect 66480 20644 66536 20646
rect 66560 20644 66616 20646
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 66320 19610 66376 19612
rect 66400 19610 66456 19612
rect 66480 19610 66536 19612
rect 66560 19610 66616 19612
rect 66320 19558 66366 19610
rect 66366 19558 66376 19610
rect 66400 19558 66430 19610
rect 66430 19558 66442 19610
rect 66442 19558 66456 19610
rect 66480 19558 66494 19610
rect 66494 19558 66506 19610
rect 66506 19558 66536 19610
rect 66560 19558 66570 19610
rect 66570 19558 66616 19610
rect 66320 19556 66376 19558
rect 66400 19556 66456 19558
rect 66480 19556 66536 19558
rect 66560 19556 66616 19558
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 55770 15952 55826 16008
rect 66320 18522 66376 18524
rect 66400 18522 66456 18524
rect 66480 18522 66536 18524
rect 66560 18522 66616 18524
rect 66320 18470 66366 18522
rect 66366 18470 66376 18522
rect 66400 18470 66430 18522
rect 66430 18470 66442 18522
rect 66442 18470 66456 18522
rect 66480 18470 66494 18522
rect 66494 18470 66506 18522
rect 66506 18470 66536 18522
rect 66560 18470 66570 18522
rect 66570 18470 66616 18522
rect 66320 18468 66376 18470
rect 66400 18468 66456 18470
rect 66480 18468 66536 18470
rect 66560 18468 66616 18470
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 66320 17434 66376 17436
rect 66400 17434 66456 17436
rect 66480 17434 66536 17436
rect 66560 17434 66616 17436
rect 66320 17382 66366 17434
rect 66366 17382 66376 17434
rect 66400 17382 66430 17434
rect 66430 17382 66442 17434
rect 66442 17382 66456 17434
rect 66480 17382 66494 17434
rect 66494 17382 66506 17434
rect 66506 17382 66536 17434
rect 66560 17382 66570 17434
rect 66570 17382 66616 17434
rect 66320 17380 66376 17382
rect 66400 17380 66456 17382
rect 66480 17380 66536 17382
rect 66560 17380 66616 17382
rect 78218 17060 78274 17096
rect 78218 17040 78220 17060
rect 78220 17040 78272 17060
rect 78272 17040 78274 17060
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 66320 16346 66376 16348
rect 66400 16346 66456 16348
rect 66480 16346 66536 16348
rect 66560 16346 66616 16348
rect 66320 16294 66366 16346
rect 66366 16294 66376 16346
rect 66400 16294 66430 16346
rect 66430 16294 66442 16346
rect 66442 16294 66456 16346
rect 66480 16294 66494 16346
rect 66494 16294 66506 16346
rect 66506 16294 66536 16346
rect 66560 16294 66570 16346
rect 66570 16294 66616 16346
rect 66320 16292 66376 16294
rect 66400 16292 66456 16294
rect 66480 16292 66536 16294
rect 66560 16292 66616 16294
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 66320 15258 66376 15260
rect 66400 15258 66456 15260
rect 66480 15258 66536 15260
rect 66560 15258 66616 15260
rect 66320 15206 66366 15258
rect 66366 15206 66376 15258
rect 66400 15206 66430 15258
rect 66430 15206 66442 15258
rect 66442 15206 66456 15258
rect 66480 15206 66494 15258
rect 66494 15206 66506 15258
rect 66506 15206 66536 15258
rect 66560 15206 66570 15258
rect 66570 15206 66616 15258
rect 66320 15204 66376 15206
rect 66400 15204 66456 15206
rect 66480 15204 66536 15206
rect 66560 15204 66616 15206
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 66320 14170 66376 14172
rect 66400 14170 66456 14172
rect 66480 14170 66536 14172
rect 66560 14170 66616 14172
rect 66320 14118 66366 14170
rect 66366 14118 66376 14170
rect 66400 14118 66430 14170
rect 66430 14118 66442 14170
rect 66442 14118 66456 14170
rect 66480 14118 66494 14170
rect 66494 14118 66506 14170
rect 66506 14118 66536 14170
rect 66560 14118 66570 14170
rect 66570 14118 66616 14170
rect 66320 14116 66376 14118
rect 66400 14116 66456 14118
rect 66480 14116 66536 14118
rect 66560 14116 66616 14118
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 66320 13082 66376 13084
rect 66400 13082 66456 13084
rect 66480 13082 66536 13084
rect 66560 13082 66616 13084
rect 66320 13030 66366 13082
rect 66366 13030 66376 13082
rect 66400 13030 66430 13082
rect 66430 13030 66442 13082
rect 66442 13030 66456 13082
rect 66480 13030 66494 13082
rect 66494 13030 66506 13082
rect 66506 13030 66536 13082
rect 66560 13030 66570 13082
rect 66570 13030 66616 13082
rect 66320 13028 66376 13030
rect 66400 13028 66456 13030
rect 66480 13028 66536 13030
rect 66560 13028 66616 13030
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 66320 11994 66376 11996
rect 66400 11994 66456 11996
rect 66480 11994 66536 11996
rect 66560 11994 66616 11996
rect 66320 11942 66366 11994
rect 66366 11942 66376 11994
rect 66400 11942 66430 11994
rect 66430 11942 66442 11994
rect 66442 11942 66456 11994
rect 66480 11942 66494 11994
rect 66494 11942 66506 11994
rect 66506 11942 66536 11994
rect 66560 11942 66570 11994
rect 66570 11942 66616 11994
rect 66320 11940 66376 11942
rect 66400 11940 66456 11942
rect 66480 11940 66536 11942
rect 66560 11940 66616 11942
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 66320 10906 66376 10908
rect 66400 10906 66456 10908
rect 66480 10906 66536 10908
rect 66560 10906 66616 10908
rect 66320 10854 66366 10906
rect 66366 10854 66376 10906
rect 66400 10854 66430 10906
rect 66430 10854 66442 10906
rect 66442 10854 66456 10906
rect 66480 10854 66494 10906
rect 66494 10854 66506 10906
rect 66506 10854 66536 10906
rect 66560 10854 66570 10906
rect 66570 10854 66616 10906
rect 66320 10852 66376 10854
rect 66400 10852 66456 10854
rect 66480 10852 66536 10854
rect 66560 10852 66616 10854
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 55494 9324 55496 9344
rect 55496 9324 55548 9344
rect 55548 9324 55550 9344
rect 55494 9288 55550 9324
rect 66320 9818 66376 9820
rect 66400 9818 66456 9820
rect 66480 9818 66536 9820
rect 66560 9818 66616 9820
rect 66320 9766 66366 9818
rect 66366 9766 66376 9818
rect 66400 9766 66430 9818
rect 66430 9766 66442 9818
rect 66442 9766 66456 9818
rect 66480 9766 66494 9818
rect 66494 9766 66506 9818
rect 66506 9766 66536 9818
rect 66560 9766 66570 9818
rect 66570 9766 66616 9818
rect 66320 9764 66376 9766
rect 66400 9764 66456 9766
rect 66480 9764 66536 9766
rect 66560 9764 66616 9766
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 66320 8730 66376 8732
rect 66400 8730 66456 8732
rect 66480 8730 66536 8732
rect 66560 8730 66616 8732
rect 66320 8678 66366 8730
rect 66366 8678 66376 8730
rect 66400 8678 66430 8730
rect 66430 8678 66442 8730
rect 66442 8678 66456 8730
rect 66480 8678 66494 8730
rect 66494 8678 66506 8730
rect 66506 8678 66536 8730
rect 66560 8678 66570 8730
rect 66570 8678 66616 8730
rect 66320 8676 66376 8678
rect 66400 8676 66456 8678
rect 66480 8676 66536 8678
rect 66560 8676 66616 8678
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 78218 8200 78274 8256
rect 66320 7642 66376 7644
rect 66400 7642 66456 7644
rect 66480 7642 66536 7644
rect 66560 7642 66616 7644
rect 66320 7590 66366 7642
rect 66366 7590 66376 7642
rect 66400 7590 66430 7642
rect 66430 7590 66442 7642
rect 66442 7590 66456 7642
rect 66480 7590 66494 7642
rect 66494 7590 66506 7642
rect 66506 7590 66536 7642
rect 66560 7590 66570 7642
rect 66570 7590 66616 7642
rect 66320 7588 66376 7590
rect 66400 7588 66456 7590
rect 66480 7588 66536 7590
rect 66560 7588 66616 7590
rect 78402 7520 78458 7576
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 66320 6554 66376 6556
rect 66400 6554 66456 6556
rect 66480 6554 66536 6556
rect 66560 6554 66616 6556
rect 66320 6502 66366 6554
rect 66366 6502 66376 6554
rect 66400 6502 66430 6554
rect 66430 6502 66442 6554
rect 66442 6502 66456 6554
rect 66480 6502 66494 6554
rect 66494 6502 66506 6554
rect 66506 6502 66536 6554
rect 66560 6502 66570 6554
rect 66570 6502 66616 6554
rect 66320 6500 66376 6502
rect 66400 6500 66456 6502
rect 66480 6500 66536 6502
rect 66560 6500 66616 6502
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 78218 6840 78274 6896
rect 66320 5466 66376 5468
rect 66400 5466 66456 5468
rect 66480 5466 66536 5468
rect 66560 5466 66616 5468
rect 66320 5414 66366 5466
rect 66366 5414 66376 5466
rect 66400 5414 66430 5466
rect 66430 5414 66442 5466
rect 66442 5414 66456 5466
rect 66480 5414 66494 5466
rect 66494 5414 66506 5466
rect 66506 5414 66536 5466
rect 66560 5414 66570 5466
rect 66570 5414 66616 5466
rect 66320 5412 66376 5414
rect 66400 5412 66456 5414
rect 66480 5412 66536 5414
rect 66560 5412 66616 5414
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 66320 4378 66376 4380
rect 66400 4378 66456 4380
rect 66480 4378 66536 4380
rect 66560 4378 66616 4380
rect 66320 4326 66366 4378
rect 66366 4326 66376 4378
rect 66400 4326 66430 4378
rect 66430 4326 66442 4378
rect 66442 4326 66456 4378
rect 66480 4326 66494 4378
rect 66494 4326 66506 4378
rect 66506 4326 66536 4378
rect 66560 4326 66570 4378
rect 66570 4326 66616 4378
rect 66320 4324 66376 4326
rect 66400 4324 66456 4326
rect 66480 4324 66536 4326
rect 66560 4324 66616 4326
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 66320 3290 66376 3292
rect 66400 3290 66456 3292
rect 66480 3290 66536 3292
rect 66560 3290 66616 3292
rect 66320 3238 66366 3290
rect 66366 3238 66376 3290
rect 66400 3238 66430 3290
rect 66430 3238 66442 3290
rect 66442 3238 66456 3290
rect 66480 3238 66494 3290
rect 66494 3238 66506 3290
rect 66506 3238 66536 3290
rect 66560 3238 66570 3290
rect 66570 3238 66616 3290
rect 66320 3236 66376 3238
rect 66400 3236 66456 3238
rect 66480 3236 66536 3238
rect 66560 3236 66616 3238
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 71134 2488 71190 2544
rect 66320 2202 66376 2204
rect 66400 2202 66456 2204
rect 66480 2202 66536 2204
rect 66560 2202 66616 2204
rect 66320 2150 66366 2202
rect 66366 2150 66376 2202
rect 66400 2150 66430 2202
rect 66430 2150 66442 2202
rect 66442 2150 66456 2202
rect 66480 2150 66494 2202
rect 66494 2150 66506 2202
rect 66506 2150 66536 2202
rect 66560 2150 66570 2202
rect 66570 2150 66616 2202
rect 66320 2148 66376 2150
rect 66400 2148 66456 2150
rect 66480 2148 66536 2150
rect 66560 2148 66616 2150
rect 74170 2488 74226 2544
rect 78218 6180 78274 6216
rect 78218 6160 78220 6180
rect 78220 6160 78272 6180
rect 78272 6160 78274 6180
rect 78402 5516 78404 5536
rect 78404 5516 78456 5536
rect 78456 5516 78458 5536
rect 78402 5480 78458 5516
rect 78310 4800 78366 4856
rect 78494 4120 78550 4176
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 66310 37024 66626 37025
rect 66310 36960 66316 37024
rect 66380 36960 66396 37024
rect 66460 36960 66476 37024
rect 66540 36960 66556 37024
rect 66620 36960 66626 37024
rect 66310 36959 66626 36960
rect 0 36818 800 36848
rect 1301 36818 1367 36821
rect 0 36816 1367 36818
rect 0 36760 1306 36816
rect 1362 36760 1367 36816
rect 0 36758 1367 36760
rect 0 36728 800 36758
rect 1301 36755 1367 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 0 36138 800 36168
rect 933 36138 999 36141
rect 0 36136 999 36138
rect 0 36080 938 36136
rect 994 36080 999 36136
rect 0 36078 999 36080
rect 0 36048 800 36078
rect 933 36075 999 36078
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 66310 35936 66626 35937
rect 66310 35872 66316 35936
rect 66380 35872 66396 35936
rect 66460 35872 66476 35936
rect 66540 35872 66556 35936
rect 66620 35872 66626 35936
rect 66310 35871 66626 35872
rect 0 35458 800 35488
rect 933 35458 999 35461
rect 0 35456 999 35458
rect 0 35400 938 35456
rect 994 35400 999 35456
rect 0 35398 999 35400
rect 0 35368 800 35398
rect 933 35395 999 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 4870 34848 5186 34849
rect 0 34778 800 34808
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 66310 34848 66626 34849
rect 66310 34784 66316 34848
rect 66380 34784 66396 34848
rect 66460 34784 66476 34848
rect 66540 34784 66556 34848
rect 66620 34784 66626 34848
rect 66310 34783 66626 34784
rect 1301 34778 1367 34781
rect 0 34776 1367 34778
rect 0 34720 1306 34776
rect 1362 34720 1367 34776
rect 0 34718 1367 34720
rect 0 34688 800 34718
rect 1301 34715 1367 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 0 34098 800 34128
rect 933 34098 999 34101
rect 0 34096 999 34098
rect 0 34040 938 34096
rect 994 34040 999 34096
rect 0 34038 999 34040
rect 0 34008 800 34038
rect 933 34035 999 34038
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 66310 33760 66626 33761
rect 66310 33696 66316 33760
rect 66380 33696 66396 33760
rect 66460 33696 66476 33760
rect 66540 33696 66556 33760
rect 66620 33696 66626 33760
rect 66310 33695 66626 33696
rect 0 33418 800 33448
rect 933 33418 999 33421
rect 0 33416 999 33418
rect 0 33360 938 33416
rect 994 33360 999 33416
rect 0 33358 999 33360
rect 0 33328 800 33358
rect 933 33355 999 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 0 32738 800 32768
rect 933 32738 999 32741
rect 0 32736 999 32738
rect 0 32680 938 32736
rect 994 32680 999 32736
rect 0 32678 999 32680
rect 0 32648 800 32678
rect 933 32675 999 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 66310 32672 66626 32673
rect 66310 32608 66316 32672
rect 66380 32608 66396 32672
rect 66460 32608 66476 32672
rect 66540 32608 66556 32672
rect 66620 32608 66626 32672
rect 66310 32607 66626 32608
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 65650 32063 65966 32064
rect 1301 32058 1367 32061
rect 0 32056 1367 32058
rect 0 32000 1306 32056
rect 1362 32000 1367 32056
rect 0 31998 1367 32000
rect 0 31968 800 31998
rect 1301 31995 1367 31998
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 66310 31584 66626 31585
rect 66310 31520 66316 31584
rect 66380 31520 66396 31584
rect 66460 31520 66476 31584
rect 66540 31520 66556 31584
rect 66620 31520 66626 31584
rect 66310 31519 66626 31520
rect 0 31378 800 31408
rect 933 31378 999 31381
rect 0 31376 999 31378
rect 0 31320 938 31376
rect 994 31320 999 31376
rect 0 31318 999 31320
rect 0 31288 800 31318
rect 933 31315 999 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 0 30698 800 30728
rect 933 30698 999 30701
rect 0 30696 999 30698
rect 0 30640 938 30696
rect 994 30640 999 30696
rect 0 30638 999 30640
rect 0 30608 800 30638
rect 933 30635 999 30638
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 66310 30496 66626 30497
rect 66310 30432 66316 30496
rect 66380 30432 66396 30496
rect 66460 30432 66476 30496
rect 66540 30432 66556 30496
rect 66620 30432 66626 30496
rect 66310 30431 66626 30432
rect 12525 30154 12591 30157
rect 14549 30154 14615 30157
rect 12525 30152 14615 30154
rect 12525 30096 12530 30152
rect 12586 30096 14554 30152
rect 14610 30096 14615 30152
rect 12525 30094 14615 30096
rect 12525 30091 12591 30094
rect 14549 30091 14615 30094
rect 0 30018 800 30048
rect 933 30018 999 30021
rect 0 30016 999 30018
rect 0 29960 938 30016
rect 994 29960 999 30016
rect 0 29958 999 29960
rect 0 29928 800 29958
rect 933 29955 999 29958
rect 44582 29956 44588 30020
rect 44652 30018 44658 30020
rect 44817 30018 44883 30021
rect 44652 30016 44883 30018
rect 44652 29960 44822 30016
rect 44878 29960 44883 30016
rect 44652 29958 44883 29960
rect 44652 29956 44658 29958
rect 44817 29955 44883 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 4870 29408 5186 29409
rect 0 29338 800 29368
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 66310 29408 66626 29409
rect 66310 29344 66316 29408
rect 66380 29344 66396 29408
rect 66460 29344 66476 29408
rect 66540 29344 66556 29408
rect 66620 29344 66626 29408
rect 66310 29343 66626 29344
rect 1301 29338 1367 29341
rect 0 29336 1367 29338
rect 0 29280 1306 29336
rect 1362 29280 1367 29336
rect 0 29278 1367 29280
rect 0 29248 800 29278
rect 1301 29275 1367 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 0 28658 800 28688
rect 933 28658 999 28661
rect 0 28656 999 28658
rect 0 28600 938 28656
rect 994 28600 999 28656
rect 0 28598 999 28600
rect 0 28568 800 28598
rect 933 28595 999 28598
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 66310 28320 66626 28321
rect 66310 28256 66316 28320
rect 66380 28256 66396 28320
rect 66460 28256 66476 28320
rect 66540 28256 66556 28320
rect 66620 28256 66626 28320
rect 66310 28255 66626 28256
rect 0 27978 800 28008
rect 933 27978 999 27981
rect 0 27976 999 27978
rect 0 27920 938 27976
rect 994 27920 999 27976
rect 0 27918 999 27920
rect 0 27888 800 27918
rect 933 27915 999 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 0 27298 800 27328
rect 933 27298 999 27301
rect 0 27296 999 27298
rect 0 27240 938 27296
rect 994 27240 999 27296
rect 0 27238 999 27240
rect 0 27208 800 27238
rect 933 27235 999 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 66310 27232 66626 27233
rect 66310 27168 66316 27232
rect 66380 27168 66396 27232
rect 66460 27168 66476 27232
rect 66540 27168 66556 27232
rect 66620 27168 66626 27232
rect 66310 27167 66626 27168
rect 4210 26688 4526 26689
rect 0 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 1301 26618 1367 26621
rect 0 26616 1367 26618
rect 0 26560 1306 26616
rect 1362 26560 1367 26616
rect 0 26558 1367 26560
rect 0 26528 800 26558
rect 1301 26555 1367 26558
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 66310 26144 66626 26145
rect 66310 26080 66316 26144
rect 66380 26080 66396 26144
rect 66460 26080 66476 26144
rect 66540 26080 66556 26144
rect 66620 26080 66626 26144
rect 66310 26079 66626 26080
rect 0 25938 800 25968
rect 933 25938 999 25941
rect 0 25936 999 25938
rect 0 25880 938 25936
rect 994 25880 999 25936
rect 0 25878 999 25880
rect 0 25848 800 25878
rect 933 25875 999 25878
rect 51809 25666 51875 25669
rect 52494 25666 52500 25668
rect 51809 25664 52500 25666
rect 51809 25608 51814 25664
rect 51870 25608 52500 25664
rect 51809 25606 52500 25608
rect 51809 25603 51875 25606
rect 52494 25604 52500 25606
rect 52564 25604 52570 25668
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 32581 25394 32647 25397
rect 34881 25394 34947 25397
rect 32581 25392 34947 25394
rect 32581 25336 32586 25392
rect 32642 25336 34886 25392
rect 34942 25336 34947 25392
rect 32581 25334 34947 25336
rect 32581 25331 32647 25334
rect 34881 25331 34947 25334
rect 0 25258 800 25288
rect 933 25258 999 25261
rect 0 25256 999 25258
rect 0 25200 938 25256
rect 994 25200 999 25256
rect 0 25198 999 25200
rect 0 25168 800 25198
rect 933 25195 999 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 66310 25056 66626 25057
rect 66310 24992 66316 25056
rect 66380 24992 66396 25056
rect 66460 24992 66476 25056
rect 66540 24992 66556 25056
rect 66620 24992 66626 25056
rect 66310 24991 66626 24992
rect 42609 24986 42675 24989
rect 44265 24986 44331 24989
rect 42609 24984 44331 24986
rect 42609 24928 42614 24984
rect 42670 24928 44270 24984
rect 44326 24928 44331 24984
rect 42609 24926 44331 24928
rect 42609 24923 42675 24926
rect 44265 24923 44331 24926
rect 0 24578 800 24608
rect 933 24578 999 24581
rect 0 24576 999 24578
rect 0 24520 938 24576
rect 994 24520 999 24576
rect 0 24518 999 24520
rect 0 24488 800 24518
rect 933 24515 999 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 40401 24034 40467 24037
rect 43529 24034 43595 24037
rect 45829 24034 45895 24037
rect 40401 24032 45895 24034
rect 40401 23976 40406 24032
rect 40462 23976 43534 24032
rect 43590 23976 45834 24032
rect 45890 23976 45895 24032
rect 40401 23974 45895 23976
rect 40401 23971 40467 23974
rect 43529 23971 43595 23974
rect 45829 23971 45895 23974
rect 4870 23968 5186 23969
rect 0 23898 800 23928
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 66310 23968 66626 23969
rect 66310 23904 66316 23968
rect 66380 23904 66396 23968
rect 66460 23904 66476 23968
rect 66540 23904 66556 23968
rect 66620 23904 66626 23968
rect 66310 23903 66626 23904
rect 1301 23898 1367 23901
rect 0 23896 1367 23898
rect 0 23840 1306 23896
rect 1362 23840 1367 23896
rect 0 23838 1367 23840
rect 0 23808 800 23838
rect 1301 23835 1367 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 0 23218 800 23248
rect 1209 23218 1275 23221
rect 0 23216 1275 23218
rect 0 23160 1214 23216
rect 1270 23160 1275 23216
rect 0 23158 1275 23160
rect 0 23128 800 23158
rect 1209 23155 1275 23158
rect 78213 23218 78279 23221
rect 79200 23218 80000 23248
rect 78213 23216 80000 23218
rect 78213 23160 78218 23216
rect 78274 23160 80000 23216
rect 78213 23158 80000 23160
rect 78213 23155 78279 23158
rect 79200 23128 80000 23158
rect 29821 23082 29887 23085
rect 31753 23082 31819 23085
rect 29821 23080 31819 23082
rect 29821 23024 29826 23080
rect 29882 23024 31758 23080
rect 31814 23024 31819 23080
rect 29821 23022 31819 23024
rect 29821 23019 29887 23022
rect 31753 23019 31819 23022
rect 44265 23082 44331 23085
rect 45369 23082 45435 23085
rect 44265 23080 45435 23082
rect 44265 23024 44270 23080
rect 44326 23024 45374 23080
rect 45430 23024 45435 23080
rect 44265 23022 45435 23024
rect 44265 23019 44331 23022
rect 45369 23019 45435 23022
rect 36169 22946 36235 22949
rect 36302 22946 36308 22948
rect 36169 22944 36308 22946
rect 36169 22888 36174 22944
rect 36230 22888 36308 22944
rect 36169 22886 36308 22888
rect 36169 22883 36235 22886
rect 36302 22884 36308 22886
rect 36372 22884 36378 22948
rect 42885 22946 42951 22949
rect 45093 22946 45159 22949
rect 49693 22948 49759 22949
rect 49693 22946 49740 22948
rect 42885 22944 45159 22946
rect 42885 22888 42890 22944
rect 42946 22888 45098 22944
rect 45154 22888 45159 22944
rect 42885 22886 45159 22888
rect 49648 22944 49740 22946
rect 49648 22888 49698 22944
rect 49648 22886 49740 22888
rect 42885 22883 42951 22886
rect 45093 22883 45159 22886
rect 49693 22884 49740 22886
rect 49804 22884 49810 22948
rect 49693 22883 49759 22884
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 66310 22880 66626 22881
rect 66310 22816 66316 22880
rect 66380 22816 66396 22880
rect 66460 22816 66476 22880
rect 66540 22816 66556 22880
rect 66620 22816 66626 22880
rect 66310 22815 66626 22816
rect 933 22674 999 22677
rect 798 22672 999 22674
rect 798 22616 938 22672
rect 994 22616 999 22672
rect 798 22614 999 22616
rect 798 22568 858 22614
rect 933 22611 999 22614
rect 38377 22674 38443 22677
rect 47393 22674 47459 22677
rect 38377 22672 47459 22674
rect 38377 22616 38382 22672
rect 38438 22616 47398 22672
rect 47454 22616 47459 22672
rect 38377 22614 47459 22616
rect 38377 22611 38443 22614
rect 47393 22611 47459 22614
rect 0 22478 858 22568
rect 38377 22538 38443 22541
rect 43161 22538 43227 22541
rect 48865 22538 48931 22541
rect 38377 22536 48931 22538
rect 38377 22480 38382 22536
rect 38438 22480 43166 22536
rect 43222 22480 48870 22536
rect 48926 22480 48931 22536
rect 38377 22478 48931 22480
rect 0 22448 800 22478
rect 38377 22475 38443 22478
rect 43161 22475 43227 22478
rect 48865 22475 48931 22478
rect 38929 22402 38995 22405
rect 39205 22402 39271 22405
rect 38929 22400 39271 22402
rect 38929 22344 38934 22400
rect 38990 22344 39210 22400
rect 39266 22344 39271 22400
rect 38929 22342 39271 22344
rect 38929 22339 38995 22342
rect 39205 22339 39271 22342
rect 40217 22402 40283 22405
rect 44449 22402 44515 22405
rect 40217 22400 44515 22402
rect 40217 22344 40222 22400
rect 40278 22344 44454 22400
rect 44510 22344 44515 22400
rect 40217 22342 44515 22344
rect 40217 22339 40283 22342
rect 44449 22339 44515 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 41873 22266 41939 22269
rect 50705 22266 50771 22269
rect 41873 22264 50771 22266
rect 41873 22208 41878 22264
rect 41934 22208 50710 22264
rect 50766 22208 50771 22264
rect 41873 22206 50771 22208
rect 41873 22203 41939 22206
rect 50705 22203 50771 22206
rect 43989 22130 44055 22133
rect 46749 22130 46815 22133
rect 43989 22128 46815 22130
rect 43989 22072 43994 22128
rect 44050 22072 46754 22128
rect 46810 22072 46815 22128
rect 43989 22070 46815 22072
rect 43989 22067 44055 22070
rect 46749 22067 46815 22070
rect 841 21994 907 21997
rect 798 21992 907 21994
rect 798 21936 846 21992
rect 902 21936 907 21992
rect 798 21931 907 21936
rect 52494 21932 52500 21996
rect 52564 21994 52570 21996
rect 53373 21994 53439 21997
rect 52564 21992 53439 21994
rect 52564 21936 53378 21992
rect 53434 21936 53439 21992
rect 52564 21934 53439 21936
rect 52564 21932 52570 21934
rect 53373 21931 53439 21934
rect 798 21888 858 21931
rect 0 21798 858 21888
rect 0 21768 800 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 66310 21792 66626 21793
rect 66310 21728 66316 21792
rect 66380 21728 66396 21792
rect 66460 21728 66476 21792
rect 66540 21728 66556 21792
rect 66620 21728 66626 21792
rect 66310 21727 66626 21728
rect 841 21314 907 21317
rect 798 21312 907 21314
rect 798 21256 846 21312
rect 902 21256 907 21312
rect 798 21251 907 21256
rect 49693 21314 49759 21317
rect 50521 21314 50587 21317
rect 49693 21312 50587 21314
rect 49693 21256 49698 21312
rect 49754 21256 50526 21312
rect 50582 21256 50587 21312
rect 49693 21254 50587 21256
rect 49693 21251 49759 21254
rect 50521 21251 50587 21254
rect 798 21208 858 21251
rect 0 21118 858 21208
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 0 21088 800 21118
rect 48405 21042 48471 21045
rect 50889 21042 50955 21045
rect 48405 21040 50955 21042
rect 48405 20984 48410 21040
rect 48466 20984 50894 21040
rect 50950 20984 50955 21040
rect 48405 20982 50955 20984
rect 48405 20979 48471 20982
rect 50889 20979 50955 20982
rect 50797 20906 50863 20909
rect 51165 20906 51231 20909
rect 50797 20904 51231 20906
rect 50797 20848 50802 20904
rect 50858 20848 51170 20904
rect 51226 20848 51231 20904
rect 50797 20846 51231 20848
rect 50797 20843 50863 20846
rect 51165 20843 51231 20846
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 66310 20704 66626 20705
rect 66310 20640 66316 20704
rect 66380 20640 66396 20704
rect 66460 20640 66476 20704
rect 66540 20640 66556 20704
rect 66620 20640 66626 20704
rect 66310 20639 66626 20640
rect 47209 20634 47275 20637
rect 48037 20634 48103 20637
rect 49734 20634 49740 20636
rect 47209 20632 49740 20634
rect 47209 20576 47214 20632
rect 47270 20576 48042 20632
rect 48098 20576 49740 20632
rect 47209 20574 49740 20576
rect 47209 20571 47275 20574
rect 48037 20571 48103 20574
rect 49734 20572 49740 20574
rect 49804 20572 49810 20636
rect 0 20498 800 20528
rect 1485 20498 1551 20501
rect 0 20496 1551 20498
rect 0 20440 1490 20496
rect 1546 20440 1551 20496
rect 0 20438 1551 20440
rect 0 20408 800 20438
rect 1485 20435 1551 20438
rect 29821 20498 29887 20501
rect 48589 20498 48655 20501
rect 29821 20496 48655 20498
rect 29821 20440 29826 20496
rect 29882 20440 48594 20496
rect 48650 20440 48655 20496
rect 29821 20438 48655 20440
rect 29821 20435 29887 20438
rect 48589 20435 48655 20438
rect 34053 20362 34119 20365
rect 39297 20362 39363 20365
rect 34053 20360 39363 20362
rect 34053 20304 34058 20360
rect 34114 20304 39302 20360
rect 39358 20304 39363 20360
rect 34053 20302 39363 20304
rect 34053 20299 34119 20302
rect 39297 20299 39363 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 44357 20090 44423 20093
rect 44582 20090 44588 20092
rect 44357 20088 44588 20090
rect 44357 20032 44362 20088
rect 44418 20032 44588 20088
rect 44357 20030 44588 20032
rect 44357 20027 44423 20030
rect 44582 20028 44588 20030
rect 44652 20090 44658 20092
rect 55121 20090 55187 20093
rect 44652 20088 55187 20090
rect 44652 20032 55126 20088
rect 55182 20032 55187 20088
rect 44652 20030 55187 20032
rect 44652 20028 44658 20030
rect 55121 20027 55187 20030
rect 0 19818 800 19848
rect 0 19728 858 19818
rect 798 19685 858 19728
rect 798 19680 907 19685
rect 798 19624 846 19680
rect 902 19624 907 19680
rect 798 19622 907 19624
rect 841 19619 907 19622
rect 36905 19682 36971 19685
rect 44725 19682 44791 19685
rect 36905 19680 44791 19682
rect 36905 19624 36910 19680
rect 36966 19624 44730 19680
rect 44786 19624 44791 19680
rect 36905 19622 44791 19624
rect 36905 19619 36971 19622
rect 44725 19619 44791 19622
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 66310 19616 66626 19617
rect 66310 19552 66316 19616
rect 66380 19552 66396 19616
rect 66460 19552 66476 19616
rect 66540 19552 66556 19616
rect 66620 19552 66626 19616
rect 66310 19551 66626 19552
rect 38285 19546 38351 19549
rect 41781 19546 41847 19549
rect 42558 19546 42564 19548
rect 38285 19544 42564 19546
rect 38285 19488 38290 19544
rect 38346 19488 41786 19544
rect 41842 19488 42564 19544
rect 38285 19486 42564 19488
rect 38285 19483 38351 19486
rect 41781 19483 41847 19486
rect 42558 19484 42564 19486
rect 42628 19484 42634 19548
rect 36302 19348 36308 19412
rect 36372 19410 36378 19412
rect 36721 19410 36787 19413
rect 37641 19412 37707 19413
rect 36372 19408 36787 19410
rect 36372 19352 36726 19408
rect 36782 19352 36787 19408
rect 36372 19350 36787 19352
rect 36372 19348 36378 19350
rect 36721 19347 36787 19350
rect 37590 19348 37596 19412
rect 37660 19410 37707 19412
rect 40309 19410 40375 19413
rect 40585 19410 40651 19413
rect 37660 19408 37752 19410
rect 37702 19352 37752 19408
rect 37660 19350 37752 19352
rect 40309 19408 40651 19410
rect 40309 19352 40314 19408
rect 40370 19352 40590 19408
rect 40646 19352 40651 19408
rect 40309 19350 40651 19352
rect 37660 19348 37707 19350
rect 37641 19347 37707 19348
rect 40309 19347 40375 19350
rect 40585 19347 40651 19350
rect 40769 19410 40835 19413
rect 41045 19410 41111 19413
rect 40769 19408 41111 19410
rect 40769 19352 40774 19408
rect 40830 19352 41050 19408
rect 41106 19352 41111 19408
rect 40769 19350 41111 19352
rect 40769 19347 40835 19350
rect 41045 19347 41111 19350
rect 31753 19274 31819 19277
rect 41045 19274 41111 19277
rect 31753 19272 41111 19274
rect 31753 19216 31758 19272
rect 31814 19216 41050 19272
rect 41106 19216 41111 19272
rect 31753 19214 41111 19216
rect 31753 19211 31819 19214
rect 41045 19211 41111 19214
rect 37365 19138 37431 19141
rect 40401 19138 40467 19141
rect 46197 19138 46263 19141
rect 37365 19136 46263 19138
rect 37365 19080 37370 19136
rect 37426 19080 40406 19136
rect 40462 19080 46202 19136
rect 46258 19080 46263 19136
rect 37365 19078 46263 19080
rect 37365 19075 37431 19078
rect 40401 19075 40467 19078
rect 46197 19075 46263 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 39849 19002 39915 19005
rect 48037 19002 48103 19005
rect 39849 19000 48103 19002
rect 39849 18944 39854 19000
rect 39910 18944 48042 19000
rect 48098 18944 48103 19000
rect 39849 18942 48103 18944
rect 39849 18939 39915 18942
rect 48037 18939 48103 18942
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 66310 18528 66626 18529
rect 66310 18464 66316 18528
rect 66380 18464 66396 18528
rect 66460 18464 66476 18528
rect 66540 18464 66556 18528
rect 66620 18464 66626 18528
rect 66310 18463 66626 18464
rect 29453 18186 29519 18189
rect 49049 18186 49115 18189
rect 29453 18184 49115 18186
rect 29453 18128 29458 18184
rect 29514 18128 49054 18184
rect 49110 18128 49115 18184
rect 29453 18126 49115 18128
rect 29453 18123 29519 18126
rect 49049 18123 49115 18126
rect 38377 18052 38443 18053
rect 38326 18050 38332 18052
rect 38286 17990 38332 18050
rect 38396 18048 38443 18052
rect 38438 17992 38443 18048
rect 38326 17988 38332 17990
rect 38396 17988 38443 17992
rect 38377 17987 38443 17988
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 40033 17778 40099 17781
rect 44541 17778 44607 17781
rect 40033 17776 44607 17778
rect 40033 17720 40038 17776
rect 40094 17720 44546 17776
rect 44602 17720 44607 17776
rect 40033 17718 44607 17720
rect 40033 17715 40099 17718
rect 44541 17715 44607 17718
rect 31385 17642 31451 17645
rect 38193 17642 38259 17645
rect 31385 17640 38259 17642
rect 31385 17584 31390 17640
rect 31446 17584 38198 17640
rect 38254 17584 38259 17640
rect 31385 17582 38259 17584
rect 31385 17579 31451 17582
rect 38193 17579 38259 17582
rect 43161 17642 43227 17645
rect 45921 17642 45987 17645
rect 43161 17640 45987 17642
rect 43161 17584 43166 17640
rect 43222 17584 45926 17640
rect 45982 17584 45987 17640
rect 43161 17582 45987 17584
rect 43161 17579 43227 17582
rect 45921 17579 45987 17582
rect 53189 17642 53255 17645
rect 54109 17642 54175 17645
rect 53189 17640 54175 17642
rect 53189 17584 53194 17640
rect 53250 17584 54114 17640
rect 54170 17584 54175 17640
rect 53189 17582 54175 17584
rect 53189 17579 53255 17582
rect 54109 17579 54175 17582
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 66310 17440 66626 17441
rect 66310 17376 66316 17440
rect 66380 17376 66396 17440
rect 66460 17376 66476 17440
rect 66540 17376 66556 17440
rect 66620 17376 66626 17440
rect 66310 17375 66626 17376
rect 30189 17234 30255 17237
rect 33593 17234 33659 17237
rect 43529 17234 43595 17237
rect 30189 17232 43595 17234
rect 30189 17176 30194 17232
rect 30250 17176 33598 17232
rect 33654 17176 43534 17232
rect 43590 17176 43595 17232
rect 30189 17174 43595 17176
rect 30189 17171 30255 17174
rect 33593 17171 33659 17174
rect 43529 17171 43595 17174
rect 31753 17098 31819 17101
rect 32949 17098 33015 17101
rect 39481 17098 39547 17101
rect 41413 17098 41479 17101
rect 31753 17096 41479 17098
rect 31753 17040 31758 17096
rect 31814 17040 32954 17096
rect 33010 17040 39486 17096
rect 39542 17040 41418 17096
rect 41474 17040 41479 17096
rect 31753 17038 41479 17040
rect 31753 17035 31819 17038
rect 32949 17035 33015 17038
rect 39481 17035 39547 17038
rect 41413 17035 41479 17038
rect 78213 17098 78279 17101
rect 79200 17098 80000 17128
rect 78213 17096 80000 17098
rect 78213 17040 78218 17096
rect 78274 17040 80000 17096
rect 78213 17038 80000 17040
rect 78213 17035 78279 17038
rect 79200 17008 80000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 23749 16418 23815 16421
rect 26693 16418 26759 16421
rect 27337 16418 27403 16421
rect 23749 16416 27403 16418
rect 23749 16360 23754 16416
rect 23810 16360 26698 16416
rect 26754 16360 27342 16416
rect 27398 16360 27403 16416
rect 23749 16358 27403 16360
rect 23749 16355 23815 16358
rect 26693 16355 26759 16358
rect 27337 16355 27403 16358
rect 49693 16418 49759 16421
rect 49918 16418 49924 16420
rect 49693 16416 49924 16418
rect 49693 16360 49698 16416
rect 49754 16360 49924 16416
rect 49693 16358 49924 16360
rect 49693 16355 49759 16358
rect 49918 16356 49924 16358
rect 49988 16356 49994 16420
rect 50245 16418 50311 16421
rect 50889 16418 50955 16421
rect 50245 16416 50955 16418
rect 50245 16360 50250 16416
rect 50306 16360 50894 16416
rect 50950 16360 50955 16416
rect 50245 16358 50955 16360
rect 50245 16355 50311 16358
rect 50889 16355 50955 16358
rect 51257 16418 51323 16421
rect 51390 16418 51396 16420
rect 51257 16416 51396 16418
rect 51257 16360 51262 16416
rect 51318 16360 51396 16416
rect 51257 16358 51396 16360
rect 51257 16355 51323 16358
rect 51390 16356 51396 16358
rect 51460 16356 51466 16420
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 66310 16352 66626 16353
rect 66310 16288 66316 16352
rect 66380 16288 66396 16352
rect 66460 16288 66476 16352
rect 66540 16288 66556 16352
rect 66620 16288 66626 16352
rect 66310 16287 66626 16288
rect 50429 16282 50495 16285
rect 53741 16282 53807 16285
rect 50429 16280 53807 16282
rect 50429 16224 50434 16280
rect 50490 16224 53746 16280
rect 53802 16224 53807 16280
rect 50429 16222 53807 16224
rect 50429 16219 50495 16222
rect 53741 16219 53807 16222
rect 44449 16146 44515 16149
rect 44582 16146 44588 16148
rect 44449 16144 44588 16146
rect 44449 16088 44454 16144
rect 44510 16088 44588 16144
rect 44449 16086 44588 16088
rect 44449 16083 44515 16086
rect 44582 16084 44588 16086
rect 44652 16084 44658 16148
rect 49509 16146 49575 16149
rect 50889 16146 50955 16149
rect 51625 16146 51691 16149
rect 49509 16144 51691 16146
rect 49509 16088 49514 16144
rect 49570 16088 50894 16144
rect 50950 16088 51630 16144
rect 51686 16088 51691 16144
rect 49509 16086 51691 16088
rect 49509 16083 49575 16086
rect 50889 16083 50955 16086
rect 51625 16083 51691 16086
rect 50429 16010 50495 16013
rect 55765 16010 55831 16013
rect 50429 16008 55831 16010
rect 50429 15952 50434 16008
rect 50490 15952 55770 16008
rect 55826 15952 55831 16008
rect 50429 15950 55831 15952
rect 50429 15947 50495 15950
rect 55765 15947 55831 15950
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 19793 15738 19859 15741
rect 27705 15738 27771 15741
rect 19793 15736 27771 15738
rect 19793 15680 19798 15736
rect 19854 15680 27710 15736
rect 27766 15680 27771 15736
rect 19793 15678 27771 15680
rect 19793 15675 19859 15678
rect 27705 15675 27771 15678
rect 21081 15602 21147 15605
rect 25221 15602 25287 15605
rect 21081 15600 25287 15602
rect 21081 15544 21086 15600
rect 21142 15544 25226 15600
rect 25282 15544 25287 15600
rect 21081 15542 25287 15544
rect 21081 15539 21147 15542
rect 25221 15539 25287 15542
rect 21265 15466 21331 15469
rect 24209 15466 24275 15469
rect 25129 15466 25195 15469
rect 21265 15464 25195 15466
rect 21265 15408 21270 15464
rect 21326 15408 24214 15464
rect 24270 15408 25134 15464
rect 25190 15408 25195 15464
rect 21265 15406 25195 15408
rect 21265 15403 21331 15406
rect 24209 15403 24275 15406
rect 25129 15403 25195 15406
rect 45829 15466 45895 15469
rect 53373 15466 53439 15469
rect 45829 15464 53439 15466
rect 45829 15408 45834 15464
rect 45890 15408 53378 15464
rect 53434 15408 53439 15464
rect 45829 15406 53439 15408
rect 45829 15403 45895 15406
rect 53373 15403 53439 15406
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 66310 15264 66626 15265
rect 66310 15200 66316 15264
rect 66380 15200 66396 15264
rect 66460 15200 66476 15264
rect 66540 15200 66556 15264
rect 66620 15200 66626 15264
rect 66310 15199 66626 15200
rect 39389 15194 39455 15197
rect 41413 15194 41479 15197
rect 39389 15192 41479 15194
rect 39389 15136 39394 15192
rect 39450 15136 41418 15192
rect 41474 15136 41479 15192
rect 39389 15134 41479 15136
rect 39389 15131 39455 15134
rect 41413 15131 41479 15134
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 33133 15058 33199 15061
rect 41045 15058 41111 15061
rect 33133 15056 41111 15058
rect 33133 15000 33138 15056
rect 33194 15000 41050 15056
rect 41106 15000 41111 15056
rect 33133 14998 41111 15000
rect 33133 14995 33199 14998
rect 41045 14995 41111 14998
rect 28165 14922 28231 14925
rect 45461 14922 45527 14925
rect 28165 14920 45527 14922
rect 28165 14864 28170 14920
rect 28226 14864 45466 14920
rect 45522 14864 45527 14920
rect 28165 14862 45527 14864
rect 28165 14859 28231 14862
rect 45461 14859 45527 14862
rect 42977 14786 43043 14789
rect 43805 14786 43871 14789
rect 49509 14786 49575 14789
rect 42977 14784 49575 14786
rect 42977 14728 42982 14784
rect 43038 14728 43810 14784
rect 43866 14728 49514 14784
rect 49570 14728 49575 14784
rect 42977 14726 49575 14728
rect 42977 14723 43043 14726
rect 43805 14723 43871 14726
rect 49509 14723 49575 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 50429 14514 50495 14517
rect 50429 14512 51320 14514
rect 50429 14456 50434 14512
rect 50490 14456 51320 14512
rect 50429 14454 51320 14456
rect 50429 14451 50495 14454
rect 0 14378 800 14408
rect 1209 14378 1275 14381
rect 0 14376 1275 14378
rect 0 14320 1214 14376
rect 1270 14320 1275 14376
rect 0 14318 1275 14320
rect 0 14288 800 14318
rect 1209 14315 1275 14318
rect 24761 14378 24827 14381
rect 27521 14378 27587 14381
rect 28625 14378 28691 14381
rect 24761 14376 28691 14378
rect 24761 14320 24766 14376
rect 24822 14320 27526 14376
rect 27582 14320 28630 14376
rect 28686 14320 28691 14376
rect 24761 14318 28691 14320
rect 24761 14315 24827 14318
rect 27521 14315 27587 14318
rect 28625 14315 28691 14318
rect 36118 14316 36124 14380
rect 36188 14378 36194 14380
rect 36629 14378 36695 14381
rect 36905 14378 36971 14381
rect 37590 14378 37596 14380
rect 36188 14376 37596 14378
rect 36188 14320 36634 14376
rect 36690 14320 36910 14376
rect 36966 14320 37596 14376
rect 36188 14318 37596 14320
rect 36188 14316 36194 14318
rect 36629 14315 36695 14318
rect 36905 14315 36971 14318
rect 37590 14316 37596 14318
rect 37660 14316 37666 14380
rect 45185 14378 45251 14381
rect 48221 14378 48287 14381
rect 45185 14376 48287 14378
rect 45185 14320 45190 14376
rect 45246 14320 48226 14376
rect 48282 14320 48287 14376
rect 45185 14318 48287 14320
rect 45185 14315 45251 14318
rect 48221 14315 48287 14318
rect 51260 14378 51320 14454
rect 53005 14378 53071 14381
rect 54753 14378 54819 14381
rect 51260 14376 54819 14378
rect 51260 14320 53010 14376
rect 53066 14320 54758 14376
rect 54814 14320 54819 14376
rect 51260 14318 54819 14320
rect 51260 14245 51320 14318
rect 53005 14315 53071 14318
rect 54753 14315 54819 14318
rect 46657 14242 46723 14245
rect 50337 14242 50403 14245
rect 46657 14240 50403 14242
rect 46657 14184 46662 14240
rect 46718 14184 50342 14240
rect 50398 14184 50403 14240
rect 46657 14182 50403 14184
rect 46657 14179 46723 14182
rect 50337 14179 50403 14182
rect 51257 14240 51323 14245
rect 51257 14184 51262 14240
rect 51318 14184 51323 14240
rect 51257 14179 51323 14184
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 66310 14176 66626 14177
rect 66310 14112 66316 14176
rect 66380 14112 66396 14176
rect 66460 14112 66476 14176
rect 66540 14112 66556 14176
rect 66620 14112 66626 14176
rect 66310 14111 66626 14112
rect 22553 14106 22619 14109
rect 27613 14106 27679 14109
rect 22553 14104 27679 14106
rect 22553 14048 22558 14104
rect 22614 14048 27618 14104
rect 27674 14048 27679 14104
rect 22553 14046 27679 14048
rect 22553 14043 22619 14046
rect 27613 14043 27679 14046
rect 50981 14106 51047 14109
rect 51901 14106 51967 14109
rect 50981 14104 51967 14106
rect 50981 14048 50986 14104
rect 51042 14048 51906 14104
rect 51962 14048 51967 14104
rect 50981 14046 51967 14048
rect 50981 14043 51047 14046
rect 51901 14043 51967 14046
rect 24853 13970 24919 13973
rect 27337 13970 27403 13973
rect 24853 13968 27403 13970
rect 24853 13912 24858 13968
rect 24914 13912 27342 13968
rect 27398 13912 27403 13968
rect 24853 13910 27403 13912
rect 24853 13907 24919 13910
rect 27337 13907 27403 13910
rect 32397 13970 32463 13973
rect 33409 13970 33475 13973
rect 32397 13968 33475 13970
rect 32397 13912 32402 13968
rect 32458 13912 33414 13968
rect 33470 13912 33475 13968
rect 32397 13910 33475 13912
rect 32397 13907 32463 13910
rect 33409 13907 33475 13910
rect 34053 13970 34119 13973
rect 40585 13970 40651 13973
rect 34053 13968 40651 13970
rect 34053 13912 34058 13968
rect 34114 13912 40590 13968
rect 40646 13912 40651 13968
rect 34053 13910 40651 13912
rect 34053 13907 34119 13910
rect 40585 13907 40651 13910
rect 25589 13834 25655 13837
rect 26417 13834 26483 13837
rect 25589 13832 26483 13834
rect 25589 13776 25594 13832
rect 25650 13776 26422 13832
rect 26478 13776 26483 13832
rect 25589 13774 26483 13776
rect 25589 13771 25655 13774
rect 26417 13771 26483 13774
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 40769 13426 40835 13429
rect 45645 13426 45711 13429
rect 40769 13424 45711 13426
rect 40769 13368 40774 13424
rect 40830 13368 45650 13424
rect 45706 13368 45711 13424
rect 40769 13366 45711 13368
rect 40769 13363 40835 13366
rect 45645 13363 45711 13366
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 66310 13088 66626 13089
rect 66310 13024 66316 13088
rect 66380 13024 66396 13088
rect 66460 13024 66476 13088
rect 66540 13024 66556 13088
rect 66620 13024 66626 13088
rect 66310 13023 66626 13024
rect 37457 12882 37523 12885
rect 38285 12884 38351 12885
rect 37590 12882 37596 12884
rect 37457 12880 37596 12882
rect 37457 12824 37462 12880
rect 37518 12824 37596 12880
rect 37457 12822 37596 12824
rect 37457 12819 37523 12822
rect 37590 12820 37596 12822
rect 37660 12882 37666 12884
rect 38285 12882 38332 12884
rect 37660 12880 38332 12882
rect 37660 12824 38290 12880
rect 37660 12822 38332 12824
rect 37660 12820 37666 12822
rect 38285 12820 38332 12822
rect 38396 12820 38402 12884
rect 38285 12819 38351 12820
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 66310 12000 66626 12001
rect 66310 11936 66316 12000
rect 66380 11936 66396 12000
rect 66460 11936 66476 12000
rect 66540 11936 66556 12000
rect 66620 11936 66626 12000
rect 66310 11935 66626 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 31201 11114 31267 11117
rect 48589 11114 48655 11117
rect 31201 11112 48655 11114
rect 31201 11056 31206 11112
rect 31262 11056 48594 11112
rect 48650 11056 48655 11112
rect 31201 11054 48655 11056
rect 31201 11051 31267 11054
rect 48589 11051 48655 11054
rect 39665 10978 39731 10981
rect 44582 10978 44588 10980
rect 39665 10976 44588 10978
rect 39665 10920 39670 10976
rect 39726 10920 44588 10976
rect 39665 10918 44588 10920
rect 39665 10915 39731 10918
rect 44582 10916 44588 10918
rect 44652 10916 44658 10980
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 66310 10912 66626 10913
rect 66310 10848 66316 10912
rect 66380 10848 66396 10912
rect 66460 10848 66476 10912
rect 66540 10848 66556 10912
rect 66620 10848 66626 10912
rect 66310 10847 66626 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 66310 9824 66626 9825
rect 66310 9760 66316 9824
rect 66380 9760 66396 9824
rect 66460 9760 66476 9824
rect 66540 9760 66556 9824
rect 66620 9760 66626 9824
rect 66310 9759 66626 9760
rect 31569 9618 31635 9621
rect 34329 9618 34395 9621
rect 31569 9616 34395 9618
rect 31569 9560 31574 9616
rect 31630 9560 34334 9616
rect 34390 9560 34395 9616
rect 31569 9558 34395 9560
rect 31569 9555 31635 9558
rect 34329 9555 34395 9558
rect 35709 9618 35775 9621
rect 37549 9618 37615 9621
rect 50337 9618 50403 9621
rect 35709 9616 37615 9618
rect 35709 9560 35714 9616
rect 35770 9560 37554 9616
rect 37610 9560 37615 9616
rect 35709 9558 37615 9560
rect 35709 9555 35775 9558
rect 37549 9555 37615 9558
rect 50294 9616 50403 9618
rect 50294 9560 50342 9616
rect 50398 9560 50403 9616
rect 50294 9555 50403 9560
rect 51390 9556 51396 9620
rect 51460 9618 51466 9620
rect 51625 9618 51691 9621
rect 51460 9616 51691 9618
rect 51460 9560 51630 9616
rect 51686 9560 51691 9616
rect 51460 9558 51691 9560
rect 51460 9556 51466 9558
rect 51625 9555 51691 9558
rect 27981 9482 28047 9485
rect 28257 9482 28323 9485
rect 33225 9482 33291 9485
rect 35985 9482 36051 9485
rect 27981 9480 36051 9482
rect 27981 9424 27986 9480
rect 28042 9424 28262 9480
rect 28318 9424 33230 9480
rect 33286 9424 35990 9480
rect 36046 9424 36051 9480
rect 27981 9422 36051 9424
rect 27981 9419 28047 9422
rect 28257 9419 28323 9422
rect 33225 9419 33291 9422
rect 35985 9419 36051 9422
rect 31661 9346 31727 9349
rect 32765 9346 32831 9349
rect 33317 9346 33383 9349
rect 31661 9344 33383 9346
rect 31661 9288 31666 9344
rect 31722 9288 32770 9344
rect 32826 9288 33322 9344
rect 33378 9288 33383 9344
rect 31661 9286 33383 9288
rect 31661 9283 31727 9286
rect 32765 9283 32831 9286
rect 33317 9283 33383 9286
rect 33777 9346 33843 9349
rect 34513 9346 34579 9349
rect 33777 9344 34579 9346
rect 33777 9288 33782 9344
rect 33838 9288 34518 9344
rect 34574 9288 34579 9344
rect 33777 9286 34579 9288
rect 33777 9283 33843 9286
rect 34513 9283 34579 9286
rect 35893 9346 35959 9349
rect 36353 9346 36419 9349
rect 42885 9346 42951 9349
rect 35893 9344 42951 9346
rect 35893 9288 35898 9344
rect 35954 9288 36358 9344
rect 36414 9288 42890 9344
rect 42946 9288 42951 9344
rect 35893 9286 42951 9288
rect 35893 9283 35959 9286
rect 36353 9283 36419 9286
rect 42885 9283 42951 9286
rect 49693 9346 49759 9349
rect 49918 9346 49924 9348
rect 49693 9344 49924 9346
rect 49693 9288 49698 9344
rect 49754 9288 49924 9344
rect 49693 9286 49924 9288
rect 49693 9283 49759 9286
rect 49918 9284 49924 9286
rect 49988 9284 49994 9348
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 50153 9210 50219 9213
rect 50294 9210 50354 9555
rect 54477 9482 54543 9485
rect 55029 9482 55095 9485
rect 54477 9480 55095 9482
rect 54477 9424 54482 9480
rect 54538 9424 55034 9480
rect 55090 9424 55095 9480
rect 54477 9422 55095 9424
rect 54477 9419 54543 9422
rect 55029 9419 55095 9422
rect 53189 9346 53255 9349
rect 55489 9346 55555 9349
rect 53189 9344 55555 9346
rect 53189 9288 53194 9344
rect 53250 9288 55494 9344
rect 55550 9288 55555 9344
rect 53189 9286 55555 9288
rect 53189 9283 53255 9286
rect 55489 9283 55555 9286
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 50153 9208 50354 9210
rect 50153 9152 50158 9208
rect 50214 9152 50354 9208
rect 50153 9150 50354 9152
rect 50153 9147 50219 9150
rect 32213 9074 32279 9077
rect 34605 9074 34671 9077
rect 32213 9072 34671 9074
rect 32213 9016 32218 9072
rect 32274 9016 34610 9072
rect 34666 9016 34671 9072
rect 32213 9014 34671 9016
rect 32213 9011 32279 9014
rect 34605 9011 34671 9014
rect 44725 9074 44791 9077
rect 49693 9074 49759 9077
rect 44725 9072 49759 9074
rect 44725 9016 44730 9072
rect 44786 9016 49698 9072
rect 49754 9016 49759 9072
rect 44725 9014 49759 9016
rect 44725 9011 44791 9014
rect 49693 9011 49759 9014
rect 29821 8938 29887 8941
rect 43621 8938 43687 8941
rect 44081 8938 44147 8941
rect 29821 8936 44147 8938
rect 29821 8880 29826 8936
rect 29882 8880 43626 8936
rect 43682 8880 44086 8936
rect 44142 8880 44147 8936
rect 29821 8878 44147 8880
rect 29821 8875 29887 8878
rect 43621 8875 43687 8878
rect 44081 8875 44147 8878
rect 49693 8938 49759 8941
rect 49918 8938 49924 8940
rect 49693 8936 49924 8938
rect 49693 8880 49698 8936
rect 49754 8880 49924 8936
rect 49693 8878 49924 8880
rect 49693 8875 49759 8878
rect 49918 8876 49924 8878
rect 49988 8938 49994 8940
rect 50981 8938 51047 8941
rect 49988 8936 51047 8938
rect 49988 8880 50986 8936
rect 51042 8880 51047 8936
rect 49988 8878 51047 8880
rect 49988 8876 49994 8878
rect 50981 8875 51047 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 66310 8736 66626 8737
rect 66310 8672 66316 8736
rect 66380 8672 66396 8736
rect 66460 8672 66476 8736
rect 66540 8672 66556 8736
rect 66620 8672 66626 8736
rect 66310 8671 66626 8672
rect 36353 8666 36419 8669
rect 36721 8666 36787 8669
rect 37590 8666 37596 8668
rect 36353 8664 37596 8666
rect 36353 8608 36358 8664
rect 36414 8608 36726 8664
rect 36782 8608 37596 8664
rect 36353 8606 37596 8608
rect 36353 8603 36419 8606
rect 36721 8603 36787 8606
rect 37590 8604 37596 8606
rect 37660 8604 37666 8668
rect 33409 8530 33475 8533
rect 35525 8530 35591 8533
rect 33409 8528 35591 8530
rect 33409 8472 33414 8528
rect 33470 8472 35530 8528
rect 35586 8472 35591 8528
rect 33409 8470 35591 8472
rect 33409 8467 33475 8470
rect 35525 8467 35591 8470
rect 42333 8530 42399 8533
rect 42558 8530 42564 8532
rect 42333 8528 42564 8530
rect 42333 8472 42338 8528
rect 42394 8472 42564 8528
rect 42333 8470 42564 8472
rect 42333 8467 42399 8470
rect 42558 8468 42564 8470
rect 42628 8530 42634 8532
rect 42885 8530 42951 8533
rect 50153 8530 50219 8533
rect 42628 8528 50219 8530
rect 42628 8472 42890 8528
rect 42946 8472 50158 8528
rect 50214 8472 50219 8528
rect 42628 8470 50219 8472
rect 42628 8468 42634 8470
rect 42885 8467 42951 8470
rect 50153 8467 50219 8470
rect 36077 8396 36143 8397
rect 36077 8394 36124 8396
rect 36032 8392 36124 8394
rect 36032 8336 36082 8392
rect 36032 8334 36124 8336
rect 36077 8332 36124 8334
rect 36188 8332 36194 8396
rect 40769 8394 40835 8397
rect 44909 8394 44975 8397
rect 40769 8392 44975 8394
rect 40769 8336 40774 8392
rect 40830 8336 44914 8392
rect 44970 8336 44975 8392
rect 40769 8334 44975 8336
rect 36077 8331 36143 8332
rect 40769 8331 40835 8334
rect 44909 8331 44975 8334
rect 43713 8258 43779 8261
rect 45277 8258 45343 8261
rect 43713 8256 45343 8258
rect 43713 8200 43718 8256
rect 43774 8200 45282 8256
rect 45338 8200 45343 8256
rect 43713 8198 45343 8200
rect 43713 8195 43779 8198
rect 45277 8195 45343 8198
rect 78213 8258 78279 8261
rect 79200 8258 80000 8288
rect 78213 8256 80000 8258
rect 78213 8200 78218 8256
rect 78274 8200 80000 8256
rect 78213 8198 80000 8200
rect 78213 8195 78279 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 79200 8168 80000 8198
rect 65650 8127 65966 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 66310 7648 66626 7649
rect 66310 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66626 7648
rect 66310 7583 66626 7584
rect 78397 7578 78463 7581
rect 79200 7578 80000 7608
rect 78397 7576 80000 7578
rect 78397 7520 78402 7576
rect 78458 7520 80000 7576
rect 78397 7518 80000 7520
rect 78397 7515 78463 7518
rect 79200 7488 80000 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 40493 7034 40559 7037
rect 41321 7034 41387 7037
rect 43713 7034 43779 7037
rect 40493 7032 43779 7034
rect 40493 6976 40498 7032
rect 40554 6976 41326 7032
rect 41382 6976 43718 7032
rect 43774 6976 43779 7032
rect 40493 6974 43779 6976
rect 40493 6971 40559 6974
rect 41321 6971 41387 6974
rect 43713 6971 43779 6974
rect 37825 6898 37891 6901
rect 45001 6898 45067 6901
rect 37825 6896 45067 6898
rect 37825 6840 37830 6896
rect 37886 6840 45006 6896
rect 45062 6840 45067 6896
rect 37825 6838 45067 6840
rect 37825 6835 37891 6838
rect 45001 6835 45067 6838
rect 78213 6898 78279 6901
rect 79200 6898 80000 6928
rect 78213 6896 80000 6898
rect 78213 6840 78218 6896
rect 78274 6840 80000 6896
rect 78213 6838 80000 6840
rect 78213 6835 78279 6838
rect 79200 6808 80000 6838
rect 41045 6762 41111 6765
rect 41505 6762 41571 6765
rect 41045 6760 41571 6762
rect 41045 6704 41050 6760
rect 41106 6704 41510 6760
rect 41566 6704 41571 6760
rect 41045 6702 41571 6704
rect 41045 6699 41111 6702
rect 41505 6699 41571 6702
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 66310 6560 66626 6561
rect 66310 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66626 6560
rect 66310 6495 66626 6496
rect 78213 6218 78279 6221
rect 79200 6218 80000 6248
rect 78213 6216 80000 6218
rect 78213 6160 78218 6216
rect 78274 6160 80000 6216
rect 78213 6158 80000 6160
rect 78213 6155 78279 6158
rect 79200 6128 80000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 78397 5538 78463 5541
rect 79200 5538 80000 5568
rect 78397 5536 80000 5538
rect 78397 5480 78402 5536
rect 78458 5480 80000 5536
rect 78397 5478 80000 5480
rect 78397 5475 78463 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 66310 5472 66626 5473
rect 66310 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66626 5472
rect 79200 5448 80000 5478
rect 66310 5407 66626 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 78305 4858 78371 4861
rect 79200 4858 80000 4888
rect 78305 4856 80000 4858
rect 78305 4800 78310 4856
rect 78366 4800 80000 4856
rect 78305 4798 80000 4800
rect 78305 4795 78371 4798
rect 79200 4768 80000 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 66310 4384 66626 4385
rect 66310 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66626 4384
rect 66310 4319 66626 4320
rect 78489 4178 78555 4181
rect 79200 4178 80000 4208
rect 78489 4176 80000 4178
rect 78489 4120 78494 4176
rect 78550 4120 80000 4176
rect 78489 4118 80000 4120
rect 78489 4115 78555 4118
rect 79200 4088 80000 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 66310 3296 66626 3297
rect 66310 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66626 3296
rect 66310 3231 66626 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 71129 2546 71195 2549
rect 74165 2546 74231 2549
rect 71129 2544 74231 2546
rect 71129 2488 71134 2544
rect 71190 2488 74170 2544
rect 74226 2488 74231 2544
rect 71129 2486 74231 2488
rect 71129 2483 71195 2486
rect 74165 2483 74231 2486
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 66310 2208 66626 2209
rect 66310 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66626 2208
rect 66310 2143 66626 2144
rect 79200 2048 80000 2168
rect 79200 1368 80000 1488
rect 79200 688 80000 808
rect 79200 8 80000 128
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 66316 37020 66380 37024
rect 66316 36964 66320 37020
rect 66320 36964 66376 37020
rect 66376 36964 66380 37020
rect 66316 36960 66380 36964
rect 66396 37020 66460 37024
rect 66396 36964 66400 37020
rect 66400 36964 66456 37020
rect 66456 36964 66460 37020
rect 66396 36960 66460 36964
rect 66476 37020 66540 37024
rect 66476 36964 66480 37020
rect 66480 36964 66536 37020
rect 66536 36964 66540 37020
rect 66476 36960 66540 36964
rect 66556 37020 66620 37024
rect 66556 36964 66560 37020
rect 66560 36964 66616 37020
rect 66616 36964 66620 37020
rect 66556 36960 66620 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 66316 35932 66380 35936
rect 66316 35876 66320 35932
rect 66320 35876 66376 35932
rect 66376 35876 66380 35932
rect 66316 35872 66380 35876
rect 66396 35932 66460 35936
rect 66396 35876 66400 35932
rect 66400 35876 66456 35932
rect 66456 35876 66460 35932
rect 66396 35872 66460 35876
rect 66476 35932 66540 35936
rect 66476 35876 66480 35932
rect 66480 35876 66536 35932
rect 66536 35876 66540 35932
rect 66476 35872 66540 35876
rect 66556 35932 66620 35936
rect 66556 35876 66560 35932
rect 66560 35876 66616 35932
rect 66616 35876 66620 35932
rect 66556 35872 66620 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 66316 34844 66380 34848
rect 66316 34788 66320 34844
rect 66320 34788 66376 34844
rect 66376 34788 66380 34844
rect 66316 34784 66380 34788
rect 66396 34844 66460 34848
rect 66396 34788 66400 34844
rect 66400 34788 66456 34844
rect 66456 34788 66460 34844
rect 66396 34784 66460 34788
rect 66476 34844 66540 34848
rect 66476 34788 66480 34844
rect 66480 34788 66536 34844
rect 66536 34788 66540 34844
rect 66476 34784 66540 34788
rect 66556 34844 66620 34848
rect 66556 34788 66560 34844
rect 66560 34788 66616 34844
rect 66616 34788 66620 34844
rect 66556 34784 66620 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 66316 33756 66380 33760
rect 66316 33700 66320 33756
rect 66320 33700 66376 33756
rect 66376 33700 66380 33756
rect 66316 33696 66380 33700
rect 66396 33756 66460 33760
rect 66396 33700 66400 33756
rect 66400 33700 66456 33756
rect 66456 33700 66460 33756
rect 66396 33696 66460 33700
rect 66476 33756 66540 33760
rect 66476 33700 66480 33756
rect 66480 33700 66536 33756
rect 66536 33700 66540 33756
rect 66476 33696 66540 33700
rect 66556 33756 66620 33760
rect 66556 33700 66560 33756
rect 66560 33700 66616 33756
rect 66616 33700 66620 33756
rect 66556 33696 66620 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 66316 32668 66380 32672
rect 66316 32612 66320 32668
rect 66320 32612 66376 32668
rect 66376 32612 66380 32668
rect 66316 32608 66380 32612
rect 66396 32668 66460 32672
rect 66396 32612 66400 32668
rect 66400 32612 66456 32668
rect 66456 32612 66460 32668
rect 66396 32608 66460 32612
rect 66476 32668 66540 32672
rect 66476 32612 66480 32668
rect 66480 32612 66536 32668
rect 66536 32612 66540 32668
rect 66476 32608 66540 32612
rect 66556 32668 66620 32672
rect 66556 32612 66560 32668
rect 66560 32612 66616 32668
rect 66616 32612 66620 32668
rect 66556 32608 66620 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 66316 31580 66380 31584
rect 66316 31524 66320 31580
rect 66320 31524 66376 31580
rect 66376 31524 66380 31580
rect 66316 31520 66380 31524
rect 66396 31580 66460 31584
rect 66396 31524 66400 31580
rect 66400 31524 66456 31580
rect 66456 31524 66460 31580
rect 66396 31520 66460 31524
rect 66476 31580 66540 31584
rect 66476 31524 66480 31580
rect 66480 31524 66536 31580
rect 66536 31524 66540 31580
rect 66476 31520 66540 31524
rect 66556 31580 66620 31584
rect 66556 31524 66560 31580
rect 66560 31524 66616 31580
rect 66616 31524 66620 31580
rect 66556 31520 66620 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 66316 30492 66380 30496
rect 66316 30436 66320 30492
rect 66320 30436 66376 30492
rect 66376 30436 66380 30492
rect 66316 30432 66380 30436
rect 66396 30492 66460 30496
rect 66396 30436 66400 30492
rect 66400 30436 66456 30492
rect 66456 30436 66460 30492
rect 66396 30432 66460 30436
rect 66476 30492 66540 30496
rect 66476 30436 66480 30492
rect 66480 30436 66536 30492
rect 66536 30436 66540 30492
rect 66476 30432 66540 30436
rect 66556 30492 66620 30496
rect 66556 30436 66560 30492
rect 66560 30436 66616 30492
rect 66616 30436 66620 30492
rect 66556 30432 66620 30436
rect 44588 29956 44652 30020
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 66316 29404 66380 29408
rect 66316 29348 66320 29404
rect 66320 29348 66376 29404
rect 66376 29348 66380 29404
rect 66316 29344 66380 29348
rect 66396 29404 66460 29408
rect 66396 29348 66400 29404
rect 66400 29348 66456 29404
rect 66456 29348 66460 29404
rect 66396 29344 66460 29348
rect 66476 29404 66540 29408
rect 66476 29348 66480 29404
rect 66480 29348 66536 29404
rect 66536 29348 66540 29404
rect 66476 29344 66540 29348
rect 66556 29404 66620 29408
rect 66556 29348 66560 29404
rect 66560 29348 66616 29404
rect 66616 29348 66620 29404
rect 66556 29344 66620 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 66316 28316 66380 28320
rect 66316 28260 66320 28316
rect 66320 28260 66376 28316
rect 66376 28260 66380 28316
rect 66316 28256 66380 28260
rect 66396 28316 66460 28320
rect 66396 28260 66400 28316
rect 66400 28260 66456 28316
rect 66456 28260 66460 28316
rect 66396 28256 66460 28260
rect 66476 28316 66540 28320
rect 66476 28260 66480 28316
rect 66480 28260 66536 28316
rect 66536 28260 66540 28316
rect 66476 28256 66540 28260
rect 66556 28316 66620 28320
rect 66556 28260 66560 28316
rect 66560 28260 66616 28316
rect 66616 28260 66620 28316
rect 66556 28256 66620 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 66316 27228 66380 27232
rect 66316 27172 66320 27228
rect 66320 27172 66376 27228
rect 66376 27172 66380 27228
rect 66316 27168 66380 27172
rect 66396 27228 66460 27232
rect 66396 27172 66400 27228
rect 66400 27172 66456 27228
rect 66456 27172 66460 27228
rect 66396 27168 66460 27172
rect 66476 27228 66540 27232
rect 66476 27172 66480 27228
rect 66480 27172 66536 27228
rect 66536 27172 66540 27228
rect 66476 27168 66540 27172
rect 66556 27228 66620 27232
rect 66556 27172 66560 27228
rect 66560 27172 66616 27228
rect 66616 27172 66620 27228
rect 66556 27168 66620 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 66316 26140 66380 26144
rect 66316 26084 66320 26140
rect 66320 26084 66376 26140
rect 66376 26084 66380 26140
rect 66316 26080 66380 26084
rect 66396 26140 66460 26144
rect 66396 26084 66400 26140
rect 66400 26084 66456 26140
rect 66456 26084 66460 26140
rect 66396 26080 66460 26084
rect 66476 26140 66540 26144
rect 66476 26084 66480 26140
rect 66480 26084 66536 26140
rect 66536 26084 66540 26140
rect 66476 26080 66540 26084
rect 66556 26140 66620 26144
rect 66556 26084 66560 26140
rect 66560 26084 66616 26140
rect 66616 26084 66620 26140
rect 66556 26080 66620 26084
rect 52500 25604 52564 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 66316 25052 66380 25056
rect 66316 24996 66320 25052
rect 66320 24996 66376 25052
rect 66376 24996 66380 25052
rect 66316 24992 66380 24996
rect 66396 25052 66460 25056
rect 66396 24996 66400 25052
rect 66400 24996 66456 25052
rect 66456 24996 66460 25052
rect 66396 24992 66460 24996
rect 66476 25052 66540 25056
rect 66476 24996 66480 25052
rect 66480 24996 66536 25052
rect 66536 24996 66540 25052
rect 66476 24992 66540 24996
rect 66556 25052 66620 25056
rect 66556 24996 66560 25052
rect 66560 24996 66616 25052
rect 66616 24996 66620 25052
rect 66556 24992 66620 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 66316 23964 66380 23968
rect 66316 23908 66320 23964
rect 66320 23908 66376 23964
rect 66376 23908 66380 23964
rect 66316 23904 66380 23908
rect 66396 23964 66460 23968
rect 66396 23908 66400 23964
rect 66400 23908 66456 23964
rect 66456 23908 66460 23964
rect 66396 23904 66460 23908
rect 66476 23964 66540 23968
rect 66476 23908 66480 23964
rect 66480 23908 66536 23964
rect 66536 23908 66540 23964
rect 66476 23904 66540 23908
rect 66556 23964 66620 23968
rect 66556 23908 66560 23964
rect 66560 23908 66616 23964
rect 66616 23908 66620 23964
rect 66556 23904 66620 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 36308 22884 36372 22948
rect 49740 22944 49804 22948
rect 49740 22888 49754 22944
rect 49754 22888 49804 22944
rect 49740 22884 49804 22888
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 66316 22876 66380 22880
rect 66316 22820 66320 22876
rect 66320 22820 66376 22876
rect 66376 22820 66380 22876
rect 66316 22816 66380 22820
rect 66396 22876 66460 22880
rect 66396 22820 66400 22876
rect 66400 22820 66456 22876
rect 66456 22820 66460 22876
rect 66396 22816 66460 22820
rect 66476 22876 66540 22880
rect 66476 22820 66480 22876
rect 66480 22820 66536 22876
rect 66536 22820 66540 22876
rect 66476 22816 66540 22820
rect 66556 22876 66620 22880
rect 66556 22820 66560 22876
rect 66560 22820 66616 22876
rect 66616 22820 66620 22876
rect 66556 22816 66620 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 52500 21932 52564 21996
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 66316 21788 66380 21792
rect 66316 21732 66320 21788
rect 66320 21732 66376 21788
rect 66376 21732 66380 21788
rect 66316 21728 66380 21732
rect 66396 21788 66460 21792
rect 66396 21732 66400 21788
rect 66400 21732 66456 21788
rect 66456 21732 66460 21788
rect 66396 21728 66460 21732
rect 66476 21788 66540 21792
rect 66476 21732 66480 21788
rect 66480 21732 66536 21788
rect 66536 21732 66540 21788
rect 66476 21728 66540 21732
rect 66556 21788 66620 21792
rect 66556 21732 66560 21788
rect 66560 21732 66616 21788
rect 66616 21732 66620 21788
rect 66556 21728 66620 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 66316 20700 66380 20704
rect 66316 20644 66320 20700
rect 66320 20644 66376 20700
rect 66376 20644 66380 20700
rect 66316 20640 66380 20644
rect 66396 20700 66460 20704
rect 66396 20644 66400 20700
rect 66400 20644 66456 20700
rect 66456 20644 66460 20700
rect 66396 20640 66460 20644
rect 66476 20700 66540 20704
rect 66476 20644 66480 20700
rect 66480 20644 66536 20700
rect 66536 20644 66540 20700
rect 66476 20640 66540 20644
rect 66556 20700 66620 20704
rect 66556 20644 66560 20700
rect 66560 20644 66616 20700
rect 66616 20644 66620 20700
rect 66556 20640 66620 20644
rect 49740 20572 49804 20636
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 44588 20028 44652 20092
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 66316 19612 66380 19616
rect 66316 19556 66320 19612
rect 66320 19556 66376 19612
rect 66376 19556 66380 19612
rect 66316 19552 66380 19556
rect 66396 19612 66460 19616
rect 66396 19556 66400 19612
rect 66400 19556 66456 19612
rect 66456 19556 66460 19612
rect 66396 19552 66460 19556
rect 66476 19612 66540 19616
rect 66476 19556 66480 19612
rect 66480 19556 66536 19612
rect 66536 19556 66540 19612
rect 66476 19552 66540 19556
rect 66556 19612 66620 19616
rect 66556 19556 66560 19612
rect 66560 19556 66616 19612
rect 66616 19556 66620 19612
rect 66556 19552 66620 19556
rect 42564 19484 42628 19548
rect 36308 19348 36372 19412
rect 37596 19408 37660 19412
rect 37596 19352 37646 19408
rect 37646 19352 37660 19408
rect 37596 19348 37660 19352
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 66316 18524 66380 18528
rect 66316 18468 66320 18524
rect 66320 18468 66376 18524
rect 66376 18468 66380 18524
rect 66316 18464 66380 18468
rect 66396 18524 66460 18528
rect 66396 18468 66400 18524
rect 66400 18468 66456 18524
rect 66456 18468 66460 18524
rect 66396 18464 66460 18468
rect 66476 18524 66540 18528
rect 66476 18468 66480 18524
rect 66480 18468 66536 18524
rect 66536 18468 66540 18524
rect 66476 18464 66540 18468
rect 66556 18524 66620 18528
rect 66556 18468 66560 18524
rect 66560 18468 66616 18524
rect 66616 18468 66620 18524
rect 66556 18464 66620 18468
rect 38332 18048 38396 18052
rect 38332 17992 38382 18048
rect 38382 17992 38396 18048
rect 38332 17988 38396 17992
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 66316 17436 66380 17440
rect 66316 17380 66320 17436
rect 66320 17380 66376 17436
rect 66376 17380 66380 17436
rect 66316 17376 66380 17380
rect 66396 17436 66460 17440
rect 66396 17380 66400 17436
rect 66400 17380 66456 17436
rect 66456 17380 66460 17436
rect 66396 17376 66460 17380
rect 66476 17436 66540 17440
rect 66476 17380 66480 17436
rect 66480 17380 66536 17436
rect 66536 17380 66540 17436
rect 66476 17376 66540 17380
rect 66556 17436 66620 17440
rect 66556 17380 66560 17436
rect 66560 17380 66616 17436
rect 66616 17380 66620 17436
rect 66556 17376 66620 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 49924 16356 49988 16420
rect 51396 16356 51460 16420
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 66316 16348 66380 16352
rect 66316 16292 66320 16348
rect 66320 16292 66376 16348
rect 66376 16292 66380 16348
rect 66316 16288 66380 16292
rect 66396 16348 66460 16352
rect 66396 16292 66400 16348
rect 66400 16292 66456 16348
rect 66456 16292 66460 16348
rect 66396 16288 66460 16292
rect 66476 16348 66540 16352
rect 66476 16292 66480 16348
rect 66480 16292 66536 16348
rect 66536 16292 66540 16348
rect 66476 16288 66540 16292
rect 66556 16348 66620 16352
rect 66556 16292 66560 16348
rect 66560 16292 66616 16348
rect 66616 16292 66620 16348
rect 66556 16288 66620 16292
rect 44588 16084 44652 16148
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 66316 15260 66380 15264
rect 66316 15204 66320 15260
rect 66320 15204 66376 15260
rect 66376 15204 66380 15260
rect 66316 15200 66380 15204
rect 66396 15260 66460 15264
rect 66396 15204 66400 15260
rect 66400 15204 66456 15260
rect 66456 15204 66460 15260
rect 66396 15200 66460 15204
rect 66476 15260 66540 15264
rect 66476 15204 66480 15260
rect 66480 15204 66536 15260
rect 66536 15204 66540 15260
rect 66476 15200 66540 15204
rect 66556 15260 66620 15264
rect 66556 15204 66560 15260
rect 66560 15204 66616 15260
rect 66616 15204 66620 15260
rect 66556 15200 66620 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 36124 14316 36188 14380
rect 37596 14316 37660 14380
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 66316 14172 66380 14176
rect 66316 14116 66320 14172
rect 66320 14116 66376 14172
rect 66376 14116 66380 14172
rect 66316 14112 66380 14116
rect 66396 14172 66460 14176
rect 66396 14116 66400 14172
rect 66400 14116 66456 14172
rect 66456 14116 66460 14172
rect 66396 14112 66460 14116
rect 66476 14172 66540 14176
rect 66476 14116 66480 14172
rect 66480 14116 66536 14172
rect 66536 14116 66540 14172
rect 66476 14112 66540 14116
rect 66556 14172 66620 14176
rect 66556 14116 66560 14172
rect 66560 14116 66616 14172
rect 66616 14116 66620 14172
rect 66556 14112 66620 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 66316 13084 66380 13088
rect 66316 13028 66320 13084
rect 66320 13028 66376 13084
rect 66376 13028 66380 13084
rect 66316 13024 66380 13028
rect 66396 13084 66460 13088
rect 66396 13028 66400 13084
rect 66400 13028 66456 13084
rect 66456 13028 66460 13084
rect 66396 13024 66460 13028
rect 66476 13084 66540 13088
rect 66476 13028 66480 13084
rect 66480 13028 66536 13084
rect 66536 13028 66540 13084
rect 66476 13024 66540 13028
rect 66556 13084 66620 13088
rect 66556 13028 66560 13084
rect 66560 13028 66616 13084
rect 66616 13028 66620 13084
rect 66556 13024 66620 13028
rect 37596 12820 37660 12884
rect 38332 12880 38396 12884
rect 38332 12824 38346 12880
rect 38346 12824 38396 12880
rect 38332 12820 38396 12824
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 66316 11996 66380 12000
rect 66316 11940 66320 11996
rect 66320 11940 66376 11996
rect 66376 11940 66380 11996
rect 66316 11936 66380 11940
rect 66396 11996 66460 12000
rect 66396 11940 66400 11996
rect 66400 11940 66456 11996
rect 66456 11940 66460 11996
rect 66396 11936 66460 11940
rect 66476 11996 66540 12000
rect 66476 11940 66480 11996
rect 66480 11940 66536 11996
rect 66536 11940 66540 11996
rect 66476 11936 66540 11940
rect 66556 11996 66620 12000
rect 66556 11940 66560 11996
rect 66560 11940 66616 11996
rect 66616 11940 66620 11996
rect 66556 11936 66620 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 44588 10916 44652 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 66316 10908 66380 10912
rect 66316 10852 66320 10908
rect 66320 10852 66376 10908
rect 66376 10852 66380 10908
rect 66316 10848 66380 10852
rect 66396 10908 66460 10912
rect 66396 10852 66400 10908
rect 66400 10852 66456 10908
rect 66456 10852 66460 10908
rect 66396 10848 66460 10852
rect 66476 10908 66540 10912
rect 66476 10852 66480 10908
rect 66480 10852 66536 10908
rect 66536 10852 66540 10908
rect 66476 10848 66540 10852
rect 66556 10908 66620 10912
rect 66556 10852 66560 10908
rect 66560 10852 66616 10908
rect 66616 10852 66620 10908
rect 66556 10848 66620 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 66316 9820 66380 9824
rect 66316 9764 66320 9820
rect 66320 9764 66376 9820
rect 66376 9764 66380 9820
rect 66316 9760 66380 9764
rect 66396 9820 66460 9824
rect 66396 9764 66400 9820
rect 66400 9764 66456 9820
rect 66456 9764 66460 9820
rect 66396 9760 66460 9764
rect 66476 9820 66540 9824
rect 66476 9764 66480 9820
rect 66480 9764 66536 9820
rect 66536 9764 66540 9820
rect 66476 9760 66540 9764
rect 66556 9820 66620 9824
rect 66556 9764 66560 9820
rect 66560 9764 66616 9820
rect 66616 9764 66620 9820
rect 66556 9760 66620 9764
rect 51396 9556 51460 9620
rect 49924 9284 49988 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 49924 8876 49988 8940
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 66316 8732 66380 8736
rect 66316 8676 66320 8732
rect 66320 8676 66376 8732
rect 66376 8676 66380 8732
rect 66316 8672 66380 8676
rect 66396 8732 66460 8736
rect 66396 8676 66400 8732
rect 66400 8676 66456 8732
rect 66456 8676 66460 8732
rect 66396 8672 66460 8676
rect 66476 8732 66540 8736
rect 66476 8676 66480 8732
rect 66480 8676 66536 8732
rect 66536 8676 66540 8732
rect 66476 8672 66540 8676
rect 66556 8732 66620 8736
rect 66556 8676 66560 8732
rect 66560 8676 66616 8732
rect 66616 8676 66620 8732
rect 66556 8672 66620 8676
rect 37596 8604 37660 8668
rect 42564 8468 42628 8532
rect 36124 8392 36188 8396
rect 36124 8336 36138 8392
rect 36138 8336 36188 8392
rect 36124 8332 36188 8336
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 66316 7644 66380 7648
rect 66316 7588 66320 7644
rect 66320 7588 66376 7644
rect 66376 7588 66380 7644
rect 66316 7584 66380 7588
rect 66396 7644 66460 7648
rect 66396 7588 66400 7644
rect 66400 7588 66456 7644
rect 66456 7588 66460 7644
rect 66396 7584 66460 7588
rect 66476 7644 66540 7648
rect 66476 7588 66480 7644
rect 66480 7588 66536 7644
rect 66536 7588 66540 7644
rect 66476 7584 66540 7588
rect 66556 7644 66620 7648
rect 66556 7588 66560 7644
rect 66560 7588 66616 7644
rect 66616 7588 66620 7644
rect 66556 7584 66620 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 66316 6556 66380 6560
rect 66316 6500 66320 6556
rect 66320 6500 66376 6556
rect 66376 6500 66380 6556
rect 66316 6496 66380 6500
rect 66396 6556 66460 6560
rect 66396 6500 66400 6556
rect 66400 6500 66456 6556
rect 66456 6500 66460 6556
rect 66396 6496 66460 6500
rect 66476 6556 66540 6560
rect 66476 6500 66480 6556
rect 66480 6500 66536 6556
rect 66536 6500 66540 6556
rect 66476 6496 66540 6500
rect 66556 6556 66620 6560
rect 66556 6500 66560 6556
rect 66560 6500 66616 6556
rect 66616 6500 66620 6556
rect 66556 6496 66620 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 66316 5468 66380 5472
rect 66316 5412 66320 5468
rect 66320 5412 66376 5468
rect 66376 5412 66380 5468
rect 66316 5408 66380 5412
rect 66396 5468 66460 5472
rect 66396 5412 66400 5468
rect 66400 5412 66456 5468
rect 66456 5412 66460 5468
rect 66396 5408 66460 5412
rect 66476 5468 66540 5472
rect 66476 5412 66480 5468
rect 66480 5412 66536 5468
rect 66536 5412 66540 5468
rect 66476 5408 66540 5412
rect 66556 5468 66620 5472
rect 66556 5412 66560 5468
rect 66560 5412 66616 5468
rect 66616 5412 66620 5468
rect 66556 5408 66620 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 66316 4380 66380 4384
rect 66316 4324 66320 4380
rect 66320 4324 66376 4380
rect 66376 4324 66380 4380
rect 66316 4320 66380 4324
rect 66396 4380 66460 4384
rect 66396 4324 66400 4380
rect 66400 4324 66456 4380
rect 66456 4324 66460 4380
rect 66396 4320 66460 4324
rect 66476 4380 66540 4384
rect 66476 4324 66480 4380
rect 66480 4324 66536 4380
rect 66536 4324 66540 4380
rect 66476 4320 66540 4324
rect 66556 4380 66620 4384
rect 66556 4324 66560 4380
rect 66560 4324 66616 4380
rect 66616 4324 66620 4380
rect 66556 4320 66620 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 66316 3292 66380 3296
rect 66316 3236 66320 3292
rect 66320 3236 66376 3292
rect 66376 3236 66380 3292
rect 66316 3232 66380 3236
rect 66396 3292 66460 3296
rect 66396 3236 66400 3292
rect 66400 3236 66456 3292
rect 66456 3236 66460 3292
rect 66396 3232 66460 3236
rect 66476 3292 66540 3296
rect 66476 3236 66480 3292
rect 66480 3236 66536 3292
rect 66536 3236 66540 3292
rect 66476 3232 66540 3236
rect 66556 3292 66620 3296
rect 66556 3236 66560 3292
rect 66560 3236 66616 3292
rect 66616 3236 66620 3292
rect 66556 3232 66620 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
rect 66316 2204 66380 2208
rect 66316 2148 66320 2204
rect 66320 2148 66376 2204
rect 66376 2148 66380 2204
rect 66316 2144 66380 2148
rect 66396 2204 66460 2208
rect 66396 2148 66400 2204
rect 66400 2148 66456 2204
rect 66456 2148 66460 2204
rect 66396 2144 66460 2148
rect 66476 2204 66540 2208
rect 66476 2148 66480 2204
rect 66480 2148 66536 2204
rect 66536 2148 66540 2204
rect 66476 2144 66540 2148
rect 66556 2204 66620 2208
rect 66556 2148 66560 2204
rect 66560 2148 66616 2204
rect 66616 2148 66620 2204
rect 66556 2144 66620 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 37024 5188 37584
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 37024 35908 37584
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 35936 35908 36960
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 65648 37568 65968 37584
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 44587 30020 44653 30021
rect 44587 29956 44588 30020
rect 44652 29956 44653 30020
rect 44587 29955 44653 29956
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 36307 22948 36373 22949
rect 36307 22884 36308 22948
rect 36372 22884 36373 22948
rect 36307 22883 36373 22884
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 36310 19413 36370 22883
rect 44590 20093 44650 29955
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 52499 25668 52565 25669
rect 52499 25604 52500 25668
rect 52564 25604 52565 25668
rect 52499 25603 52565 25604
rect 49739 22948 49805 22949
rect 49739 22884 49740 22948
rect 49804 22884 49805 22948
rect 49739 22883 49805 22884
rect 49742 20637 49802 22883
rect 52502 21997 52562 25603
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 52499 21996 52565 21997
rect 52499 21932 52500 21996
rect 52564 21932 52565 21996
rect 52499 21931 52565 21932
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 49739 20636 49805 20637
rect 49739 20572 49740 20636
rect 49804 20572 49805 20636
rect 49739 20571 49805 20572
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 44587 20092 44653 20093
rect 44587 20028 44588 20092
rect 44652 20028 44653 20092
rect 44587 20027 44653 20028
rect 42563 19548 42629 19549
rect 42563 19484 42564 19548
rect 42628 19484 42629 19548
rect 42563 19483 42629 19484
rect 36307 19412 36373 19413
rect 36307 19348 36308 19412
rect 36372 19348 36373 19412
rect 36307 19347 36373 19348
rect 37595 19412 37661 19413
rect 37595 19348 37596 19412
rect 37660 19348 37661 19412
rect 37595 19347 37661 19348
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 37598 14381 37658 19347
rect 38331 18052 38397 18053
rect 38331 17988 38332 18052
rect 38396 17988 38397 18052
rect 38331 17987 38397 17988
rect 36123 14380 36189 14381
rect 36123 14316 36124 14380
rect 36188 14316 36189 14380
rect 36123 14315 36189 14316
rect 37595 14380 37661 14381
rect 37595 14316 37596 14380
rect 37660 14316 37661 14380
rect 37595 14315 37661 14316
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 36126 8397 36186 14315
rect 38334 12885 38394 17987
rect 37595 12884 37661 12885
rect 37595 12820 37596 12884
rect 37660 12820 37661 12884
rect 37595 12819 37661 12820
rect 38331 12884 38397 12885
rect 38331 12820 38332 12884
rect 38396 12820 38397 12884
rect 38331 12819 38397 12820
rect 37598 8669 37658 12819
rect 37595 8668 37661 8669
rect 37595 8604 37596 8668
rect 37660 8604 37661 8668
rect 37595 8603 37661 8604
rect 42566 8533 42626 19483
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 49923 16420 49989 16421
rect 49923 16356 49924 16420
rect 49988 16356 49989 16420
rect 49923 16355 49989 16356
rect 51395 16420 51461 16421
rect 51395 16356 51396 16420
rect 51460 16356 51461 16420
rect 51395 16355 51461 16356
rect 44587 16148 44653 16149
rect 44587 16084 44588 16148
rect 44652 16084 44653 16148
rect 44587 16083 44653 16084
rect 44590 10981 44650 16083
rect 44587 10980 44653 10981
rect 44587 10916 44588 10980
rect 44652 10916 44653 10980
rect 44587 10915 44653 10916
rect 49926 9349 49986 16355
rect 51398 9621 51458 16355
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 51395 9620 51461 9621
rect 51395 9556 51396 9620
rect 51460 9556 51461 9620
rect 51395 9555 51461 9556
rect 49923 9348 49989 9349
rect 49923 9284 49924 9348
rect 49988 9284 49989 9348
rect 49923 9283 49989 9284
rect 49926 8941 49986 9283
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 49923 8940 49989 8941
rect 49923 8876 49924 8940
rect 49988 8876 49989 8940
rect 49923 8875 49989 8876
rect 42563 8532 42629 8533
rect 42563 8468 42564 8532
rect 42628 8468 42629 8532
rect 42563 8467 42629 8468
rect 36123 8396 36189 8397
rect 36123 8332 36124 8396
rect 36188 8332 36189 8396
rect 36123 8331 36189 8332
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 5472 35908 6496
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
rect 66308 37024 66628 37584
rect 66308 36960 66316 37024
rect 66380 36960 66396 37024
rect 66460 36960 66476 37024
rect 66540 36960 66556 37024
rect 66620 36960 66628 37024
rect 66308 35936 66628 36960
rect 66308 35872 66316 35936
rect 66380 35872 66396 35936
rect 66460 35872 66476 35936
rect 66540 35872 66556 35936
rect 66620 35872 66628 35936
rect 66308 34848 66628 35872
rect 66308 34784 66316 34848
rect 66380 34784 66396 34848
rect 66460 34784 66476 34848
rect 66540 34784 66556 34848
rect 66620 34784 66628 34848
rect 66308 33760 66628 34784
rect 66308 33696 66316 33760
rect 66380 33696 66396 33760
rect 66460 33696 66476 33760
rect 66540 33696 66556 33760
rect 66620 33696 66628 33760
rect 66308 32672 66628 33696
rect 66308 32608 66316 32672
rect 66380 32608 66396 32672
rect 66460 32608 66476 32672
rect 66540 32608 66556 32672
rect 66620 32608 66628 32672
rect 66308 31584 66628 32608
rect 66308 31520 66316 31584
rect 66380 31520 66396 31584
rect 66460 31520 66476 31584
rect 66540 31520 66556 31584
rect 66620 31520 66628 31584
rect 66308 30496 66628 31520
rect 66308 30432 66316 30496
rect 66380 30432 66396 30496
rect 66460 30432 66476 30496
rect 66540 30432 66556 30496
rect 66620 30432 66628 30496
rect 66308 29408 66628 30432
rect 66308 29344 66316 29408
rect 66380 29344 66396 29408
rect 66460 29344 66476 29408
rect 66540 29344 66556 29408
rect 66620 29344 66628 29408
rect 66308 28320 66628 29344
rect 66308 28256 66316 28320
rect 66380 28256 66396 28320
rect 66460 28256 66476 28320
rect 66540 28256 66556 28320
rect 66620 28256 66628 28320
rect 66308 27232 66628 28256
rect 66308 27168 66316 27232
rect 66380 27168 66396 27232
rect 66460 27168 66476 27232
rect 66540 27168 66556 27232
rect 66620 27168 66628 27232
rect 66308 26144 66628 27168
rect 66308 26080 66316 26144
rect 66380 26080 66396 26144
rect 66460 26080 66476 26144
rect 66540 26080 66556 26144
rect 66620 26080 66628 26144
rect 66308 25056 66628 26080
rect 66308 24992 66316 25056
rect 66380 24992 66396 25056
rect 66460 24992 66476 25056
rect 66540 24992 66556 25056
rect 66620 24992 66628 25056
rect 66308 23968 66628 24992
rect 66308 23904 66316 23968
rect 66380 23904 66396 23968
rect 66460 23904 66476 23968
rect 66540 23904 66556 23968
rect 66620 23904 66628 23968
rect 66308 22880 66628 23904
rect 66308 22816 66316 22880
rect 66380 22816 66396 22880
rect 66460 22816 66476 22880
rect 66540 22816 66556 22880
rect 66620 22816 66628 22880
rect 66308 21792 66628 22816
rect 66308 21728 66316 21792
rect 66380 21728 66396 21792
rect 66460 21728 66476 21792
rect 66540 21728 66556 21792
rect 66620 21728 66628 21792
rect 66308 20704 66628 21728
rect 66308 20640 66316 20704
rect 66380 20640 66396 20704
rect 66460 20640 66476 20704
rect 66540 20640 66556 20704
rect 66620 20640 66628 20704
rect 66308 19616 66628 20640
rect 66308 19552 66316 19616
rect 66380 19552 66396 19616
rect 66460 19552 66476 19616
rect 66540 19552 66556 19616
rect 66620 19552 66628 19616
rect 66308 18528 66628 19552
rect 66308 18464 66316 18528
rect 66380 18464 66396 18528
rect 66460 18464 66476 18528
rect 66540 18464 66556 18528
rect 66620 18464 66628 18528
rect 66308 17440 66628 18464
rect 66308 17376 66316 17440
rect 66380 17376 66396 17440
rect 66460 17376 66476 17440
rect 66540 17376 66556 17440
rect 66620 17376 66628 17440
rect 66308 16352 66628 17376
rect 66308 16288 66316 16352
rect 66380 16288 66396 16352
rect 66460 16288 66476 16352
rect 66540 16288 66556 16352
rect 66620 16288 66628 16352
rect 66308 15264 66628 16288
rect 66308 15200 66316 15264
rect 66380 15200 66396 15264
rect 66460 15200 66476 15264
rect 66540 15200 66556 15264
rect 66620 15200 66628 15264
rect 66308 14176 66628 15200
rect 66308 14112 66316 14176
rect 66380 14112 66396 14176
rect 66460 14112 66476 14176
rect 66540 14112 66556 14176
rect 66620 14112 66628 14176
rect 66308 13088 66628 14112
rect 66308 13024 66316 13088
rect 66380 13024 66396 13088
rect 66460 13024 66476 13088
rect 66540 13024 66556 13088
rect 66620 13024 66628 13088
rect 66308 12000 66628 13024
rect 66308 11936 66316 12000
rect 66380 11936 66396 12000
rect 66460 11936 66476 12000
rect 66540 11936 66556 12000
rect 66620 11936 66628 12000
rect 66308 10912 66628 11936
rect 66308 10848 66316 10912
rect 66380 10848 66396 10912
rect 66460 10848 66476 10912
rect 66540 10848 66556 10912
rect 66620 10848 66628 10912
rect 66308 9824 66628 10848
rect 66308 9760 66316 9824
rect 66380 9760 66396 9824
rect 66460 9760 66476 9824
rect 66540 9760 66556 9824
rect 66620 9760 66628 9824
rect 66308 8736 66628 9760
rect 66308 8672 66316 8736
rect 66380 8672 66396 8736
rect 66460 8672 66476 8736
rect 66540 8672 66556 8736
rect 66620 8672 66628 8736
rect 66308 7648 66628 8672
rect 66308 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66628 7648
rect 66308 6560 66628 7584
rect 66308 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66628 6560
rect 66308 5472 66628 6496
rect 66308 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66628 5472
rect 66308 4384 66628 5408
rect 66308 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66628 4384
rect 66308 3296 66628 4320
rect 66308 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66628 3296
rect 66308 2208 66628 3232
rect 66308 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66628 2208
rect 66308 2128 66628 2144
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1
transform 1 0 48208 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1
transform -1 0 43516 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1
transform 1 0 45816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1
transform 1 0 45908 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1
transform -1 0 21620 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1
transform 1 0 17664 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1
transform 1 0 34040 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1
transform 1 0 40572 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1
transform 1 0 55292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0740_
timestamp 1
transform -1 0 66700 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0741_
timestamp 1
transform 1 0 58696 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0742_
timestamp 1
transform 1 0 54556 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0743_
timestamp 1
transform -1 0 59892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0744_
timestamp 1
transform 1 0 59892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0745_
timestamp 1
transform -1 0 73140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_1  _0746_
timestamp 1
transform 1 0 73968 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0747_
timestamp 1
transform -1 0 72772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0748_
timestamp 1
transform 1 0 70932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0749_
timestamp 1
transform 1 0 72036 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0750_
timestamp 1
transform -1 0 72680 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1
transform 1 0 58972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0752_
timestamp 1
transform -1 0 58972 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0753_
timestamp 1
transform 1 0 57868 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _0754_
timestamp 1
transform 1 0 19228 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__or4b_2  _0755_
timestamp 1
transform -1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0756_
timestamp 1
transform 1 0 23092 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1
transform 1 0 28612 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0758_
timestamp 1
transform 1 0 19228 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0759_
timestamp 1
transform -1 0 19044 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0760_
timestamp 1
transform 1 0 19688 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0762_
timestamp 1
transform 1 0 12328 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0763_
timestamp 1
transform 1 0 15640 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0764_
timestamp 1
transform 1 0 15916 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0765_
timestamp 1
transform 1 0 12788 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0766_
timestamp 1
transform 1 0 13984 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0767_
timestamp 1
transform -1 0 15640 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0768_
timestamp 1
transform 1 0 16652 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0769_
timestamp 1
transform -1 0 19136 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0770_
timestamp 1
transform 1 0 16836 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0771_
timestamp 1
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0772_
timestamp 1
transform 1 0 17756 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0773_
timestamp 1
transform 1 0 18400 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0774_
timestamp 1
transform 1 0 18124 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0775_
timestamp 1
transform 1 0 18216 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_4  _0776_
timestamp 1
transform -1 0 18400 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__a31oi_2  _0777_
timestamp 1
transform 1 0 18676 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1
transform 1 0 20792 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0779_
timestamp 1
transform 1 0 17020 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _0780_
timestamp 1
transform 1 0 7452 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1
transform -1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0782_
timestamp 1
transform -1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0783_
timestamp 1
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0784_
timestamp 1
transform 1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0785_
timestamp 1
transform 1 0 12880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0786_
timestamp 1
transform -1 0 20424 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0787_
timestamp 1
transform -1 0 17756 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0788_
timestamp 1
transform -1 0 19136 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0789_
timestamp 1
transform -1 0 16284 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _0790_
timestamp 1
transform 1 0 12696 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0791_
timestamp 1
transform 1 0 10764 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0792_
timestamp 1
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0793_
timestamp 1
transform -1 0 15640 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0794_
timestamp 1
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0795_
timestamp 1
transform 1 0 14352 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0796_
timestamp 1
transform 1 0 15088 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0797_
timestamp 1
transform 1 0 12696 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0798_
timestamp 1
transform 1 0 12880 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0799_
timestamp 1
transform -1 0 15732 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0800_
timestamp 1
transform -1 0 14536 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0801_
timestamp 1
transform 1 0 14628 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0802_
timestamp 1
transform -1 0 13432 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0803_
timestamp 1
transform 1 0 13432 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0804_
timestamp 1
transform -1 0 12604 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0805_
timestamp 1
transform 1 0 10580 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0806_
timestamp 1
transform -1 0 11132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0807_
timestamp 1
transform 1 0 10580 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0808_
timestamp 1
transform -1 0 10120 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0809_
timestamp 1
transform -1 0 10764 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0810_
timestamp 1
transform -1 0 9568 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0811_
timestamp 1
transform 1 0 12236 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0812_
timestamp 1
transform -1 0 12972 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0813_
timestamp 1
transform 1 0 12328 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0814_
timestamp 1
transform 1 0 11500 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0815_
timestamp 1
transform -1 0 12236 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0816_
timestamp 1
transform -1 0 11224 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1
transform -1 0 10856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0818_
timestamp 1
transform -1 0 10580 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0819_
timestamp 1
transform -1 0 11132 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1
transform 1 0 10948 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0821_
timestamp 1
transform 1 0 10212 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0822_
timestamp 1
transform 1 0 11132 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0823_
timestamp 1
transform -1 0 10948 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1
transform 1 0 10948 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0825_
timestamp 1
transform -1 0 12052 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0826_
timestamp 1
transform 1 0 11224 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0827_
timestamp 1
transform 1 0 10948 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0828_
timestamp 1
transform 1 0 11592 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0829_
timestamp 1
transform 1 0 12236 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0830_
timestamp 1
transform -1 0 13340 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0831_
timestamp 1
transform 1 0 13340 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0832_
timestamp 1
transform -1 0 16560 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0833_
timestamp 1
transform 1 0 15180 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0835_
timestamp 1
transform 1 0 15640 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0836_
timestamp 1
transform 1 0 15364 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0837_
timestamp 1
transform -1 0 16192 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0838_
timestamp 1
transform -1 0 15548 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0839_
timestamp 1
transform 1 0 15732 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0840_
timestamp 1
transform -1 0 15640 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0841_
timestamp 1
transform 1 0 16560 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0842_
timestamp 1
transform -1 0 17480 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0843_
timestamp 1
transform 1 0 17204 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0844_
timestamp 1
transform 1 0 17480 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0845_
timestamp 1
transform -1 0 18584 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0846_
timestamp 1
transform 1 0 18400 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0847_
timestamp 1
transform 1 0 17940 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0848_
timestamp 1
transform -1 0 19504 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0849_
timestamp 1
transform 1 0 19872 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0850_
timestamp 1
transform -1 0 20516 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0851_
timestamp 1
transform -1 0 21068 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0852_
timestamp 1
transform -1 0 20700 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0853_
timestamp 1
transform 1 0 19964 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0854_
timestamp 1
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0855_
timestamp 1
transform 1 0 21068 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0856_
timestamp 1
transform -1 0 19964 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0857_
timestamp 1
transform -1 0 20332 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0858_
timestamp 1
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0859_
timestamp 1
transform 1 0 19136 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0860_
timestamp 1
transform -1 0 17296 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0861_
timestamp 1
transform -1 0 17848 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0862_
timestamp 1
transform -1 0 17664 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0863_
timestamp 1
transform -1 0 17204 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0864_
timestamp 1
transform 1 0 17388 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0865_
timestamp 1
transform -1 0 18768 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0866_
timestamp 1
transform -1 0 17664 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _0867_
timestamp 1
transform -1 0 32200 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0868_
timestamp 1
transform 1 0 29532 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0869_
timestamp 1
transform -1 0 32844 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0870_
timestamp 1
transform 1 0 32016 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1
transform 1 0 38180 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0872_
timestamp 1
transform -1 0 36984 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0873_
timestamp 1
transform -1 0 36708 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0874_
timestamp 1
transform -1 0 35788 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1
transform 1 0 35420 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0876_
timestamp 1
transform -1 0 36616 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0877_
timestamp 1
transform -1 0 35236 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 1
transform -1 0 36524 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0879_
timestamp 1
transform -1 0 36800 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0880_
timestamp 1
transform 1 0 36064 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0881_
timestamp 1
transform 1 0 37260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0882_
timestamp 1
transform -1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0883_
timestamp 1
transform 1 0 36708 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0884_
timestamp 1
transform 1 0 39744 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0885_
timestamp 1
transform 1 0 40940 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0886_
timestamp 1
transform 1 0 40020 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0887_
timestamp 1
transform 1 0 40480 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0888_
timestamp 1
transform 1 0 40848 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0889_
timestamp 1
transform 1 0 40572 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0890_
timestamp 1
transform 1 0 41308 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0891_
timestamp 1
transform -1 0 45632 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1
transform -1 0 44712 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _0893_
timestamp 1
transform 1 0 44252 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _0894_
timestamp 1
transform -1 0 42228 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0895_
timestamp 1
transform -1 0 45632 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_4  _0896_
timestamp 1
transform -1 0 44988 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_4  _0897_
timestamp 1
transform 1 0 43700 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0898_
timestamp 1
transform -1 0 41768 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1
transform -1 0 40756 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0900_
timestamp 1
transform -1 0 41400 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0901_
timestamp 1
transform 1 0 40756 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0902_
timestamp 1
transform -1 0 40296 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0903_
timestamp 1
transform -1 0 39744 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0904_
timestamp 1
transform 1 0 38916 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0905_
timestamp 1
transform -1 0 40112 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0906_
timestamp 1
transform 1 0 36984 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0907_
timestamp 1
transform 1 0 37904 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0908_
timestamp 1
transform -1 0 45816 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0909_
timestamp 1
transform -1 0 46276 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0910_
timestamp 1
transform 1 0 44712 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0911_
timestamp 1
transform 1 0 46092 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0912_
timestamp 1
transform 1 0 46552 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0913_
timestamp 1
transform 1 0 46920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0914_
timestamp 1
transform -1 0 48024 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0915_
timestamp 1
transform -1 0 48392 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 1
transform -1 0 47288 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0917_
timestamp 1
transform 1 0 45816 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0918_
timestamp 1
transform -1 0 46828 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1
transform 1 0 46920 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0920_
timestamp 1
transform -1 0 48024 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _0921_
timestamp 1
transform 1 0 45632 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0922_
timestamp 1
transform 1 0 45908 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0923_
timestamp 1
transform 1 0 44344 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0924_
timestamp 1
transform -1 0 45448 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0925_
timestamp 1
transform -1 0 44160 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _0926_
timestamp 1
transform 1 0 43148 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0927_
timestamp 1
transform 1 0 43148 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0928_
timestamp 1
transform -1 0 53912 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0929_
timestamp 1
transform -1 0 56580 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0930_
timestamp 1
transform -1 0 57592 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0931_
timestamp 1
transform 1 0 42412 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0932_
timestamp 1
transform 1 0 46092 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0933_
timestamp 1
transform 1 0 44988 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_2  _0934_
timestamp 1
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0935_
timestamp 1
transform -1 0 20056 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _0936_
timestamp 1
transform 1 0 17756 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1
transform -1 0 21252 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0938_
timestamp 1
transform 1 0 18584 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0939_
timestamp 1
transform -1 0 23460 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0940_
timestamp 1
transform 1 0 19228 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0941_
timestamp 1
transform -1 0 23828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0942_
timestamp 1
transform -1 0 30268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1
transform 1 0 29256 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0944_
timestamp 1
transform -1 0 30268 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0945_
timestamp 1
transform 1 0 30728 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0946_
timestamp 1
transform 1 0 28888 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1
transform -1 0 29164 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1
transform 1 0 30268 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0949_
timestamp 1
transform -1 0 37076 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0950_
timestamp 1
transform 1 0 36432 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0951_
timestamp 1
transform 1 0 43332 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0952_
timestamp 1
transform -1 0 44528 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0953_
timestamp 1
transform -1 0 48944 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0954_
timestamp 1
transform 1 0 47656 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0955_
timestamp 1
transform -1 0 48484 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0956_
timestamp 1
transform 1 0 46368 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0957_
timestamp 1
transform 1 0 32936 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0958_
timestamp 1
transform 1 0 33764 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0959_
timestamp 1
transform -1 0 30176 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0960_
timestamp 1
transform 1 0 29808 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0961_
timestamp 1
transform 1 0 30452 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0962_
timestamp 1
transform -1 0 49404 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0963_
timestamp 1
transform 1 0 48576 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0964_
timestamp 1
transform -1 0 32936 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0965_
timestamp 1
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0966_
timestamp 1
transform -1 0 39100 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0967_
timestamp 1
transform -1 0 38548 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0968_
timestamp 1
transform 1 0 41400 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0969_
timestamp 1
transform 1 0 41860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0970_
timestamp 1
transform -1 0 49220 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0971_
timestamp 1
transform 1 0 47932 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0972_
timestamp 1
transform 1 0 47656 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0973_
timestamp 1
transform 1 0 48392 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0974_
timestamp 1
transform 1 0 31280 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0975_
timestamp 1
transform 1 0 31372 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0976_
timestamp 1
transform -1 0 30544 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0977_
timestamp 1
transform 1 0 29532 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0978_
timestamp 1
transform 1 0 50324 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0979_
timestamp 1
transform 1 0 50600 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0980_
timestamp 1
transform -1 0 34500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0981_
timestamp 1
transform 1 0 33672 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0982_
timestamp 1
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0983_
timestamp 1
transform -1 0 41584 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0984_
timestamp 1
transform -1 0 43056 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0985_
timestamp 1
transform 1 0 40756 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0986_
timestamp 1
transform -1 0 49312 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0987_
timestamp 1
transform 1 0 48576 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0988_
timestamp 1
transform -1 0 50784 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0989_
timestamp 1
transform 1 0 50140 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0990_
timestamp 1
transform 1 0 32016 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0991_
timestamp 1
transform 1 0 32844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0992_
timestamp 1
transform -1 0 33396 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0993_
timestamp 1
transform 1 0 32108 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0994_
timestamp 1
transform 1 0 52256 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0995_
timestamp 1
transform 1 0 52716 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0996_
timestamp 1
transform -1 0 36248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0997_
timestamp 1
transform 1 0 35420 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0998_
timestamp 1
transform 1 0 42964 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0999_
timestamp 1
transform 1 0 43148 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1000_
timestamp 1
transform -1 0 41676 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1001_
timestamp 1
transform 1 0 40388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1002_
timestamp 1
transform -1 0 50324 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1003_
timestamp 1
transform 1 0 49312 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1004_
timestamp 1
transform 1 0 51060 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1005_
timestamp 1
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1006_
timestamp 1
transform -1 0 31556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1007_
timestamp 1
transform 1 0 30176 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1008_
timestamp 1
transform 1 0 30084 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1009_
timestamp 1
transform 1 0 30728 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1010_
timestamp 1
transform 1 0 54372 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1011_
timestamp 1
transform -1 0 55476 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1012_
timestamp 1
transform -1 0 37996 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1013_
timestamp 1
transform 1 0 37720 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1014_
timestamp 1
transform 1 0 40848 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1015_
timestamp 1
transform -1 0 42964 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1016_
timestamp 1
transform 1 0 42412 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1017_
timestamp 1
transform 1 0 42964 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1018_
timestamp 1
transform -1 0 50876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1019_
timestamp 1
transform 1 0 49496 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1020_
timestamp 1
transform -1 0 55108 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1021_
timestamp 1
transform 1 0 53820 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1022_
timestamp 1
transform -1 0 32108 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1023_
timestamp 1
transform 1 0 30728 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1024_
timestamp 1
transform -1 0 31740 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1025_
timestamp 1
transform 1 0 30360 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1026_
timestamp 1
transform 1 0 54556 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1027_
timestamp 1
transform -1 0 56672 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1028_
timestamp 1
transform 1 0 39468 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1029_
timestamp 1
transform 1 0 40204 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1030_
timestamp 1
transform 1 0 39468 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1031_
timestamp 1
transform 1 0 39652 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1032_
timestamp 1
transform 1 0 40480 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1033_
timestamp 1
transform -1 0 42504 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1034_
timestamp 1
transform 1 0 50876 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1035_
timestamp 1
transform 1 0 51704 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1036_
timestamp 1
transform 1 0 54280 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1037_
timestamp 1
transform 1 0 55292 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1038_
timestamp 1
transform -1 0 31924 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1039_
timestamp 1
transform 1 0 30912 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1040_
timestamp 1
transform -1 0 31648 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1041_
timestamp 1
transform 1 0 30544 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1042_
timestamp 1
transform 1 0 52716 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1043_
timestamp 1
transform 1 0 52900 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1044_
timestamp 1
transform 1 0 41400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1045_
timestamp 1
transform 1 0 42412 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1046_
timestamp 1
transform 1 0 37996 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1047_
timestamp 1
transform -1 0 39744 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1048_
timestamp 1
transform -1 0 42136 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1049_
timestamp 1
transform 1 0 40480 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1050_
timestamp 1
transform -1 0 54188 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1051_
timestamp 1
transform 1 0 53360 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1052_
timestamp 1
transform 1 0 51888 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1053_
timestamp 1
transform 1 0 52716 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1054_
timestamp 1
transform 1 0 34684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1055_
timestamp 1
transform 1 0 35052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1056_
timestamp 1
transform -1 0 33028 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1057_
timestamp 1
transform -1 0 32752 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1058_
timestamp 1
transform 1 0 54280 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1059_
timestamp 1
transform -1 0 55476 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1060_
timestamp 1
transform 1 0 43332 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1061_
timestamp 1
transform 1 0 44068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1062_
timestamp 1
transform -1 0 37904 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1063_
timestamp 1
transform 1 0 36432 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1064_
timestamp 1
transform -1 0 42320 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1065_
timestamp 1
transform 1 0 41032 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1066_
timestamp 1
transform -1 0 55936 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1067_
timestamp 1
transform -1 0 55016 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1068_
timestamp 1
transform 1 0 53820 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1069_
timestamp 1
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1070_
timestamp 1
transform 1 0 33028 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1071_
timestamp 1
transform -1 0 34132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1072_
timestamp 1
transform -1 0 35328 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1073_
timestamp 1
transform 1 0 33304 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1074_
timestamp 1
transform 1 0 55292 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1075_
timestamp 1
transform -1 0 55752 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1076_
timestamp 1
transform 1 0 44988 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1077_
timestamp 1
transform 1 0 45264 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1078_
timestamp 1
transform 1 0 34868 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1079_
timestamp 1
transform 1 0 34684 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1080_
timestamp 1
transform -1 0 43332 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1081_
timestamp 1
transform 1 0 43332 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1082_
timestamp 1
transform -1 0 54188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1083_
timestamp 1
transform 1 0 53268 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1084_
timestamp 1
transform 1 0 53912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1085_
timestamp 1
transform -1 0 54924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1086_
timestamp 1
transform -1 0 34224 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1087_
timestamp 1
transform 1 0 32936 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1088_
timestamp 1
transform -1 0 35328 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1089_
timestamp 1
transform 1 0 33948 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1090_
timestamp 1
transform 1 0 52808 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1091_
timestamp 1
transform 1 0 53176 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1092_
timestamp 1
transform 1 0 42228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1093_
timestamp 1
transform 1 0 42780 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1094_
timestamp 1
transform -1 0 35328 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1095_
timestamp 1
transform 1 0 33304 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1096_
timestamp 1
transform 1 0 44988 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1097_
timestamp 1
transform 1 0 45080 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1098_
timestamp 1
transform 1 0 51244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1099_
timestamp 1
transform 1 0 51520 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1100_
timestamp 1
transform 1 0 52716 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1101_
timestamp 1
transform -1 0 54280 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1102_
timestamp 1
transform 1 0 34684 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1103_
timestamp 1
transform 1 0 35236 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1104_
timestamp 1
transform -1 0 35328 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1105_
timestamp 1
transform 1 0 33856 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1106_
timestamp 1
transform 1 0 50784 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1107_
timestamp 1
transform 1 0 51428 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1108_
timestamp 1
transform 1 0 39744 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1109_
timestamp 1
transform 1 0 40388 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1110_
timestamp 1
transform 1 0 33212 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1111_
timestamp 1
transform 1 0 33856 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1112_
timestamp 1
transform 1 0 46644 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1113_
timestamp 1
transform -1 0 47932 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1114_
timestamp 1
transform 1 0 51888 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1115_
timestamp 1
transform 1 0 52808 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1116_
timestamp 1
transform 1 0 50232 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1117_
timestamp 1
transform 1 0 50968 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1118_
timestamp 1
transform -1 0 36708 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1119_
timestamp 1
transform 1 0 36156 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1120_
timestamp 1
transform -1 0 35880 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1121_
timestamp 1
transform 1 0 35144 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1122_
timestamp 1
transform 1 0 52716 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1123_
timestamp 1
transform -1 0 54096 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1124_
timestamp 1
transform 1 0 37720 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1125_
timestamp 1
transform 1 0 38180 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1126_
timestamp 1
transform -1 0 35328 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1127_
timestamp 1
transform 1 0 34224 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1128_
timestamp 1
transform 1 0 44436 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1129_
timestamp 1
transform -1 0 46736 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1130_
timestamp 1
transform 1 0 54464 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1131_
timestamp 1
transform -1 0 55752 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1132_
timestamp 1
transform 1 0 47748 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1133_
timestamp 1
transform 1 0 48208 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1134_
timestamp 1
transform 1 0 36616 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1135_
timestamp 1
transform 1 0 37260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1136_
timestamp 1
transform 1 0 36340 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1137_
timestamp 1
transform 1 0 36616 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1138_
timestamp 1
transform 1 0 50876 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1139_
timestamp 1
transform 1 0 51060 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1140_
timestamp 1
transform -1 0 37168 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1141_
timestamp 1
transform 1 0 36248 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1142_
timestamp 1
transform -1 0 33028 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1143_
timestamp 1
transform 1 0 32108 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1144_
timestamp 1
transform 1 0 46368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1145_
timestamp 1
transform -1 0 47656 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1146_
timestamp 1
transform 1 0 54188 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1147_
timestamp 1
transform 1 0 54464 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1148_
timestamp 1
transform 1 0 45724 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1149_
timestamp 1
transform 1 0 45816 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1150_
timestamp 1
transform -1 0 38824 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1151_
timestamp 1
transform 1 0 38272 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1152_
timestamp 1
transform 1 0 37996 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1153_
timestamp 1
transform 1 0 38088 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1154_
timestamp 1
transform 1 0 49312 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1155_
timestamp 1
transform 1 0 49128 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1156_
timestamp 1
transform 1 0 34960 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1157_
timestamp 1
transform 1 0 34868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1158_
timestamp 1
transform 1 0 32108 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1159_
timestamp 1
transform 1 0 32108 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1160_
timestamp 1
transform 1 0 45356 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1161_
timestamp 1
transform 1 0 45632 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1162_
timestamp 1
transform 1 0 51980 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1163_
timestamp 1
transform 1 0 52624 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1164_
timestamp 1
transform -1 0 47104 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1165_
timestamp 1
transform 1 0 44988 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1166_
timestamp 1
transform 1 0 38180 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1167_
timestamp 1
transform 1 0 38180 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1168_
timestamp 1
transform 1 0 37536 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1169_
timestamp 1
transform 1 0 38180 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1170_
timestamp 1
transform -1 0 49680 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1171_
timestamp 1
transform 1 0 48392 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1172_
timestamp 1
transform 1 0 33028 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1173_
timestamp 1
transform 1 0 33764 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1174_
timestamp 1
transform -1 0 33304 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1175_
timestamp 1
transform 1 0 31096 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1176_
timestamp 1
transform -1 0 47840 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1177_
timestamp 1
transform -1 0 47380 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1178_
timestamp 1
transform -1 0 51796 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1179_
timestamp 1
transform 1 0 50692 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1180_
timestamp 1
transform 1 0 45816 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1181_
timestamp 1
transform -1 0 46828 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1182_
timestamp 1
transform -1 0 39468 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1183_
timestamp 1
transform -1 0 39008 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1184_
timestamp 1
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1185_
timestamp 1
transform 1 0 36432 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1186_
timestamp 1
transform -1 0 49588 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1187_
timestamp 1
transform 1 0 48024 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1188_
timestamp 1
transform 1 0 31004 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1189_
timestamp 1
transform 1 0 31464 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_4  _1190_
timestamp 1
transform 1 0 19596 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1191_
timestamp 1
transform -1 0 20608 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1192_
timestamp 1
transform 1 0 20240 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1193_
timestamp 1
transform 1 0 18032 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _1194_
timestamp 1
transform 1 0 44068 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1195_
timestamp 1
transform 1 0 40848 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1196_
timestamp 1
transform 1 0 43884 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1197_
timestamp 1
transform 1 0 45080 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a2111oi_1  _1198_
timestamp 1
transform -1 0 46460 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1199_
timestamp 1
transform 1 0 45448 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1200_
timestamp 1
transform 1 0 46092 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1201_
timestamp 1
transform -1 0 46368 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1202_
timestamp 1
transform -1 0 46736 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1203_
timestamp 1
transform -1 0 46368 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1204_
timestamp 1
transform 1 0 43700 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1205_
timestamp 1
transform -1 0 48392 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1206_
timestamp 1
transform 1 0 48484 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1207_
timestamp 1
transform 1 0 44620 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1208_
timestamp 1
transform 1 0 44988 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1209_
timestamp 1
transform 1 0 44344 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1210_
timestamp 1
transform -1 0 44528 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1211_
timestamp 1
transform -1 0 44068 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1212_
timestamp 1
transform -1 0 48392 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1213_
timestamp 1
transform 1 0 46092 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1214_
timestamp 1
transform -1 0 43240 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _1215_
timestamp 1
transform 1 0 45816 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1216_
timestamp 1
transform 1 0 42504 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1217_
timestamp 1
transform 1 0 42596 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_1  _1218_
timestamp 1
transform -1 0 43516 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _1219_
timestamp 1
transform 1 0 42504 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1220_
timestamp 1
transform -1 0 43148 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1221_
timestamp 1
transform 1 0 42412 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_2  _1222_
timestamp 1
transform 1 0 43332 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 1
transform -1 0 42780 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1224_
timestamp 1
transform 1 0 40480 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1225_
timestamp 1
transform -1 0 45080 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1226_
timestamp 1
transform 1 0 43240 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1227_
timestamp 1
transform 1 0 40756 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1228_
timestamp 1
transform 1 0 40388 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1229_
timestamp 1
transform 1 0 44068 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _1230_
timestamp 1
transform 1 0 44528 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1231_
timestamp 1
transform 1 0 45908 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1232_
timestamp 1
transform 1 0 17664 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1233_
timestamp 1
transform 1 0 12788 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1234_
timestamp 1
transform 1 0 11776 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1235_
timestamp 1
transform 1 0 15088 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1236_
timestamp 1
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1237_
timestamp 1
transform 1 0 15732 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1238_
timestamp 1
transform 1 0 13432 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1239_
timestamp 1
transform 1 0 11960 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _1240_
timestamp 1
transform 1 0 20148 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_1  _1241_
timestamp 1
transform -1 0 21896 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1242_
timestamp 1
transform 1 0 21068 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1243_
timestamp 1
transform 1 0 35972 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1244_
timestamp 1
transform 1 0 39284 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1245_
timestamp 1
transform 1 0 38732 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1246_
timestamp 1
transform -1 0 37076 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1247_
timestamp 1
transform 1 0 35604 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1248_
timestamp 1
transform -1 0 35972 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1249_
timestamp 1
transform 1 0 34684 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1250_
timestamp 1
transform 1 0 36156 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1251_
timestamp 1
transform 1 0 34684 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1252_
timestamp 1
transform -1 0 35880 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1253_
timestamp 1
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1254_
timestamp 1
transform -1 0 35328 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1255_
timestamp 1
transform 1 0 33672 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1256_
timestamp 1
transform 1 0 32568 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1257_
timestamp 1
transform -1 0 32568 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1258_
timestamp 1
transform -1 0 32016 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1259_
timestamp 1
transform 1 0 32936 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1260_
timestamp 1
transform -1 0 32660 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1261_
timestamp 1
transform 1 0 32108 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1262_
timestamp 1
transform -1 0 30912 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1263_
timestamp 1
transform 1 0 28152 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1264_
timestamp 1
transform -1 0 29992 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1265_
timestamp 1
transform -1 0 29164 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 1
transform -1 0 28520 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1267_
timestamp 1
transform -1 0 29256 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 1
transform 1 0 28244 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1269_
timestamp 1
transform -1 0 28060 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1270_
timestamp 1
transform -1 0 28060 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1271_
timestamp 1
transform -1 0 30084 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1272_
timestamp 1
transform -1 0 29900 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1273_
timestamp 1
transform 1 0 31096 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1274_
timestamp 1
transform 1 0 29624 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1275_
timestamp 1
transform -1 0 29624 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 1
transform 1 0 29992 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1277_
timestamp 1
transform -1 0 32384 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1278_
timestamp 1
transform 1 0 31372 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1279_
timestamp 1
transform 1 0 31372 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _1280_
timestamp 1
transform 1 0 20148 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1281_
timestamp 1
transform -1 0 23276 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp 1
transform -1 0 23460 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _1283_
timestamp 1
transform 1 0 20056 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__o22ai_2  _1284_
timestamp 1
transform -1 0 21712 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1285_
timestamp 1
transform -1 0 23184 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1286_
timestamp 1
transform -1 0 22724 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1287_
timestamp 1
transform -1 0 20792 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1288_
timestamp 1
transform 1 0 25300 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1289_
timestamp 1
transform -1 0 23000 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1290_
timestamp 1
transform -1 0 26496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1291_
timestamp 1
transform -1 0 22908 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1292_
timestamp 1
transform -1 0 28244 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1293_
timestamp 1
transform -1 0 26404 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1294_
timestamp 1
transform 1 0 27324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1295_
timestamp 1
transform 1 0 23000 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1296_
timestamp 1
transform 1 0 23460 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1297_
timestamp 1
transform 1 0 27416 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1298_
timestamp 1
transform 1 0 23920 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1
transform 1 0 23920 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1300_
timestamp 1
transform -1 0 23000 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _1301_
timestamp 1
transform 1 0 20700 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1302_
timestamp 1
transform 1 0 25208 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _1303_
timestamp 1
transform -1 0 28612 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _1304_
timestamp 1
transform 1 0 28060 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1305_
timestamp 1
transform 1 0 23460 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o311ai_4  _1306_
timestamp 1
transform 1 0 26036 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _1307_
timestamp 1
transform 1 0 29532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1308_
timestamp 1
transform -1 0 26128 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1309_
timestamp 1
transform -1 0 27508 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1310_
timestamp 1
transform 1 0 24288 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1311_
timestamp 1
transform -1 0 24840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1312_
timestamp 1
transform 1 0 23736 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1313_
timestamp 1
transform 1 0 23092 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1314_
timestamp 1
transform 1 0 23276 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1315_
timestamp 1
transform 1 0 22908 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1316_
timestamp 1
transform -1 0 26864 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1317_
timestamp 1
transform 1 0 25392 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1318_
timestamp 1
transform 1 0 25024 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1319_
timestamp 1
transform -1 0 29808 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1320_
timestamp 1
transform 1 0 21344 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1321_
timestamp 1
transform 1 0 24380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1322_
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1323_
timestamp 1
transform -1 0 28428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1324_
timestamp 1
transform -1 0 23460 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1325_
timestamp 1
transform 1 0 27232 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1326_
timestamp 1
transform -1 0 25668 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1327_
timestamp 1
transform -1 0 26404 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_2  _1328_
timestamp 1
transform -1 0 28888 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1329_
timestamp 1
transform -1 0 25760 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1330_
timestamp 1
transform -1 0 29072 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1331_
timestamp 1
transform 1 0 24380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1332_
timestamp 1
transform 1 0 25208 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1333_
timestamp 1
transform 1 0 27784 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1334_
timestamp 1
transform -1 0 28704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1335_
timestamp 1
transform 1 0 28244 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1336_
timestamp 1
transform 1 0 28428 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1337_
timestamp 1
transform -1 0 23828 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1338_
timestamp 1
transform 1 0 22172 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1339_
timestamp 1
transform 1 0 23184 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1340_
timestamp 1
transform 1 0 23644 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1341_
timestamp 1
transform 1 0 27048 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1342_
timestamp 1
transform -1 0 26496 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1343_
timestamp 1
transform 1 0 26404 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1344_
timestamp 1
transform -1 0 26496 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1345_
timestamp 1
transform 1 0 29716 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1346_
timestamp 1
transform 1 0 22540 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1347_
timestamp 1
transform 1 0 27324 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1348_
timestamp 1
transform -1 0 25852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1349_
timestamp 1
transform 1 0 27876 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1350_
timestamp 1
transform 1 0 28796 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1351_
timestamp 1
transform 1 0 27048 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1352_
timestamp 1
transform 1 0 27140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1353_
timestamp 1
transform 1 0 26404 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1354_
timestamp 1
transform -1 0 26864 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1355_
timestamp 1
transform 1 0 26588 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1356_
timestamp 1
transform -1 0 26036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1357_
timestamp 1
transform 1 0 25576 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1358_
timestamp 1
transform 1 0 24288 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1359_
timestamp 1
transform 1 0 27784 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1360_
timestamp 1
transform 1 0 27048 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1361_
timestamp 1
transform 1 0 26036 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1362_
timestamp 1
transform -1 0 27600 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1363_
timestamp 1
transform 1 0 28152 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1364_
timestamp 1
transform 1 0 28336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1365_
timestamp 1
transform -1 0 30544 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1366_
timestamp 1
transform 1 0 29900 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1367_
timestamp 1
transform -1 0 44344 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _1368_
timestamp 1
transform -1 0 43884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1369_
timestamp 1
transform 1 0 46092 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1370_
timestamp 1
transform -1 0 44712 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1371_
timestamp 1
transform 1 0 42412 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1372_
timestamp 1
transform 1 0 43424 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _1373_
timestamp 1
transform 1 0 42228 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3b_1  _1374_
timestamp 1
transform -1 0 41400 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1375_
timestamp 1
transform 1 0 47288 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1376_
timestamp 1
transform 1 0 44988 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1377_
timestamp 1
transform 1 0 43332 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1378_
timestamp 1
transform -1 0 42136 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1379_
timestamp 1
transform 1 0 42412 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1380_
timestamp 1
transform 1 0 11316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1381_
timestamp 1
transform -1 0 10028 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1382_
timestamp 1
transform -1 0 8004 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1383_
timestamp 1
transform -1 0 7820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1384_
timestamp 1
transform 1 0 7544 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1385_
timestamp 1
transform -1 0 8832 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1386_
timestamp 1
transform -1 0 7544 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1387_
timestamp 1
transform 1 0 6992 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1388_
timestamp 1
transform 1 0 7360 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _1389_
timestamp 1
transform 1 0 9292 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1390_
timestamp 1
transform -1 0 10672 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1391_
timestamp 1
transform 1 0 45172 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _1392_
timestamp 1
transform 1 0 47564 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1393_
timestamp 1
transform -1 0 42504 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1394_
timestamp 1
transform 1 0 46460 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1395_
timestamp 1
transform 1 0 45816 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1396_
timestamp 1
transform -1 0 42228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1397_
timestamp 1
transform 1 0 42412 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1398_
timestamp 1
transform -1 0 43424 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1399_
timestamp 1
transform -1 0 42964 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1400_
timestamp 1
transform 1 0 46460 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1401_
timestamp 1
transform -1 0 43240 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1402_
timestamp 1
transform 1 0 44988 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1403_
timestamp 1
transform -1 0 42596 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1404_
timestamp 1
transform 1 0 45724 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1405_
timestamp 1
transform 1 0 46644 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1406_
timestamp 1
transform -1 0 44068 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1407_
timestamp 1
transform 1 0 44068 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1408_
timestamp 1
transform -1 0 45448 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1409_
timestamp 1
transform 1 0 35696 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1410_
timestamp 1
transform 1 0 36524 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1411_
timestamp 1
transform 1 0 35880 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1412_
timestamp 1
transform -1 0 40756 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1413_
timestamp 1
transform 1 0 36156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1414_
timestamp 1
transform 1 0 37536 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1415_
timestamp 1
transform 1 0 37352 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1416_
timestamp 1
transform 1 0 38824 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1417_
timestamp 1
transform -1 0 40296 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1418_
timestamp 1
transform 1 0 38088 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1419_
timestamp 1
transform 1 0 38272 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1420_
timestamp 1
transform -1 0 44896 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1421_
timestamp 1
transform 1 0 43976 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1422_
timestamp 1
transform 1 0 42044 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1423_
timestamp 1
transform 1 0 43424 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1424_
timestamp 1
transform -1 0 44528 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1425_
timestamp 1
transform 1 0 42596 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1426_
timestamp 1
transform 1 0 44620 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1427_
timestamp 1
transform -1 0 46644 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1428_
timestamp 1
transform -1 0 43792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1429_
timestamp 1
transform -1 0 43976 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1430_
timestamp 1
transform -1 0 43792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1431_
timestamp 1
transform -1 0 51244 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1432_
timestamp 1
transform 1 0 49128 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1433_
timestamp 1
transform 1 0 49772 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1
transform 1 0 49220 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1435_
timestamp 1
transform 1 0 50324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1436_
timestamp 1
transform -1 0 50784 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1437_
timestamp 1
transform 1 0 50324 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1438_
timestamp 1
transform 1 0 50784 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1439_
timestamp 1
transform -1 0 51796 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1440_
timestamp 1
transform 1 0 51244 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1441_
timestamp 1
transform 1 0 50140 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1442_
timestamp 1
transform -1 0 51244 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1443_
timestamp 1
transform -1 0 44804 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1444_
timestamp 1
transform -1 0 49312 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1445_
timestamp 1
transform -1 0 51520 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1446_
timestamp 1
transform -1 0 49956 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1447_
timestamp 1
transform 1 0 50140 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1448_
timestamp 1
transform 1 0 50140 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1449_
timestamp 1
transform 1 0 50416 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1450_
timestamp 1
transform -1 0 51704 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1451_
timestamp 1
transform 1 0 45080 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1452_
timestamp 1
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1453_
timestamp 1
transform 1 0 48300 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1454_
timestamp 1
transform 1 0 49864 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1455_
timestamp 1
transform -1 0 56488 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 1
transform 1 0 34960 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1457_
timestamp 1
transform -1 0 37444 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1458_
timestamp 1
transform 1 0 34868 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1459_
timestamp 1
transform 1 0 35880 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1460_
timestamp 1
transform 1 0 35052 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1461_
timestamp 1
transform 1 0 35788 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1462_
timestamp 1
transform -1 0 39376 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1463_
timestamp 1
transform 1 0 36616 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1464_
timestamp 1
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1465_
timestamp 1
transform -1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1466_
timestamp 1
transform 1 0 37536 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1467_
timestamp 1
transform 1 0 35328 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1468_
timestamp 1
transform 1 0 34868 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1469_
timestamp 1
transform -1 0 39928 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1470_
timestamp 1
transform -1 0 39192 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1471_
timestamp 1
transform 1 0 39836 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1472_
timestamp 1
transform 1 0 36064 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1473_
timestamp 1
transform -1 0 37904 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1474_
timestamp 1
transform 1 0 35236 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1475_
timestamp 1
transform -1 0 36892 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1476_
timestamp 1
transform 1 0 36524 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1477_
timestamp 1
transform -1 0 40296 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1478_
timestamp 1
transform -1 0 39652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1479_
timestamp 1
transform 1 0 49956 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1480_
timestamp 1
transform 1 0 50600 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1481_
timestamp 1
transform 1 0 51060 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1482_
timestamp 1
transform 1 0 49220 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1483_
timestamp 1
transform 1 0 49680 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1484_
timestamp 1
transform 1 0 50600 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1485_
timestamp 1
transform 1 0 48392 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1486_
timestamp 1
transform 1 0 50508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1487_
timestamp 1
transform 1 0 51244 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1488_
timestamp 1
transform -1 0 56948 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1489_
timestamp 1
transform 1 0 36708 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1490_
timestamp 1
transform 1 0 36064 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1491_
timestamp 1
transform -1 0 41400 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1492_
timestamp 1
transform 1 0 37260 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1493_
timestamp 1
transform 1 0 38088 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1494_
timestamp 1
transform -1 0 42872 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1495_
timestamp 1
transform 1 0 39836 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1496_
timestamp 1
transform 1 0 40020 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1497_
timestamp 1
transform 1 0 36248 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1498_
timestamp 1
transform -1 0 37536 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o41ai_1  _1499_
timestamp 1
transform 1 0 39100 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1500_
timestamp 1
transform 1 0 39928 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1501_
timestamp 1
transform -1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1502_
timestamp 1
transform -1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1503_
timestamp 1
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1504_
timestamp 1
transform -1 0 9016 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1505_
timestamp 1
transform 1 0 56120 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1506_
timestamp 1
transform 1 0 17848 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1507_
timestamp 1
transform 1 0 17112 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1508_
timestamp 1
transform 1 0 36156 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1509_
timestamp 1
transform 1 0 43976 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1510_
timestamp 1
transform 1 0 47104 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1511_
timestamp 1
transform 1 0 45724 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1512_
timestamp 1
transform 1 0 33580 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1513_
timestamp 1
transform 1 0 29532 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1514_
timestamp 1
transform 1 0 48116 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1515_
timestamp 1
transform 1 0 31280 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1516_
timestamp 1
transform 1 0 38548 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1517_
timestamp 1
transform 1 0 41768 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1518_
timestamp 1
transform 1 0 47564 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1519_
timestamp 1
transform 1 0 47840 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1520_
timestamp 1
transform 1 0 30912 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1521_
timestamp 1
transform 1 0 27968 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1522_
timestamp 1
transform 1 0 50508 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1523_
timestamp 1
transform 1 0 33212 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1524_
timestamp 1
transform 1 0 41032 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1525_
timestamp 1
transform 1 0 39928 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1526_
timestamp 1
transform 1 0 48208 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1527_
timestamp 1
transform 1 0 49864 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1528_
timestamp 1
transform 1 0 32752 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1529_
timestamp 1
transform 1 0 32016 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1530_
timestamp 1
transform 1 0 52716 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1531_
timestamp 1
transform 1 0 35236 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1532_
timestamp 1
transform 1 0 42780 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1533_
timestamp 1
transform 1 0 39836 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1534_
timestamp 1
transform 1 0 49404 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1535_
timestamp 1
transform 1 0 51796 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1536_
timestamp 1
transform 1 0 28888 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1537_
timestamp 1
transform 1 0 30084 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1538_
timestamp 1
transform -1 0 57132 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1539_
timestamp 1
transform 1 0 37536 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1540_
timestamp 1
transform -1 0 42320 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1541_
timestamp 1
transform 1 0 42964 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1542_
timestamp 1
transform -1 0 51980 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1543_
timestamp 1
transform 1 0 53636 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1544_
timestamp 1
transform 1 0 29808 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1545_
timestamp 1
transform 1 0 28428 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1546_
timestamp 1
transform -1 0 57040 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1547_
timestamp 1
transform 1 0 39836 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1548_
timestamp 1
transform 1 0 39836 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1549_
timestamp 1
transform -1 0 41952 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1550_
timestamp 1
transform 1 0 51520 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1551_
timestamp 1
transform 1 0 54832 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1552_
timestamp 1
transform 1 0 30360 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1553_
timestamp 1
transform 1 0 29716 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1554_
timestamp 1
transform 1 0 52716 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1555_
timestamp 1
transform 1 0 41860 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1556_
timestamp 1
transform -1 0 40112 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1557_
timestamp 1
transform 1 0 39836 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1558_
timestamp 1
transform 1 0 53360 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1559_
timestamp 1
transform 1 0 51980 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1560_
timestamp 1
transform 1 0 34776 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1561_
timestamp 1
transform 1 0 32108 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1562_
timestamp 1
transform -1 0 57132 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1563_
timestamp 1
transform 1 0 43792 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1564_
timestamp 1
transform -1 0 37812 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1565_
timestamp 1
transform 1 0 41124 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1566_
timestamp 1
transform 1 0 55016 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1567_
timestamp 1
transform 1 0 54372 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1568_
timestamp 1
transform -1 0 34408 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1569_
timestamp 1
transform 1 0 32752 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1570_
timestamp 1
transform 1 0 55292 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1571_
timestamp 1
transform 1 0 45080 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1572_
timestamp 1
transform 1 0 33856 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1573_
timestamp 1
transform 1 0 42780 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1574_
timestamp 1
transform 1 0 53084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1575_
timestamp 1
transform -1 0 56488 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1576_
timestamp 1
transform 1 0 32016 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1577_
timestamp 1
transform 1 0 33396 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1578_
timestamp 1
transform 1 0 52992 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1579_
timestamp 1
transform 1 0 42688 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1580_
timestamp 1
transform 1 0 32108 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1581_
timestamp 1
transform 1 0 44988 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1582_
timestamp 1
transform 1 0 51152 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1583_
timestamp 1
transform -1 0 54372 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1584_
timestamp 1
transform -1 0 36156 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1585_
timestamp 1
transform 1 0 32844 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1586_
timestamp 1
transform 1 0 50784 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1587_
timestamp 1
transform 1 0 40388 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1588_
timestamp 1
transform 1 0 33580 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1589_
timestamp 1
transform -1 0 49404 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1590_
timestamp 1
transform 1 0 52624 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1591_
timestamp 1
transform 1 0 50232 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1592_
timestamp 1
transform 1 0 35328 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1593_
timestamp 1
transform 1 0 34776 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1594_
timestamp 1
transform -1 0 54556 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1595_
timestamp 1
transform 1 0 37904 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1596_
timestamp 1
transform 1 0 33856 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1597_
timestamp 1
transform -1 0 46828 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1598_
timestamp 1
transform 1 0 55292 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1599_
timestamp 1
transform 1 0 48024 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1600_
timestamp 1
transform 1 0 36892 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1601_
timestamp 1
transform 1 0 36340 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1602_
timestamp 1
transform 1 0 50324 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1603_
timestamp 1
transform 1 0 35696 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1604_
timestamp 1
transform 1 0 31556 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1605_
timestamp 1
transform -1 0 49404 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1606_
timestamp 1
transform 1 0 54188 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1607_
timestamp 1
transform 1 0 45264 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1608_
timestamp 1
transform 1 0 37812 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1609_
timestamp 1
transform 1 0 37812 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1610_
timestamp 1
transform 1 0 48484 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1611_
timestamp 1
transform 1 0 34408 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1612_
timestamp 1
transform 1 0 31096 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1613_
timestamp 1
transform 1 0 45264 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1614_
timestamp 1
transform 1 0 52440 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1615_
timestamp 1
transform 1 0 43056 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1616_
timestamp 1
transform 1 0 37628 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1617_
timestamp 1
transform 1 0 37812 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1618_
timestamp 1
transform 1 0 47656 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1619_
timestamp 1
transform -1 0 34316 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1620_
timestamp 1
transform 1 0 30176 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1621_
timestamp 1
transform -1 0 47472 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1622_
timestamp 1
transform 1 0 50324 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1623_
timestamp 1
transform 1 0 46828 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1624_
timestamp 1
transform -1 0 39100 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1625_
timestamp 1
transform 1 0 35696 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1626_
timestamp 1
transform 1 0 47288 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1627_
timestamp 1
transform 1 0 31096 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1628_
timestamp 1
transform 1 0 15180 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1629_
timestamp 1
transform -1 0 21528 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1630_
timestamp 1
transform 1 0 14260 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1631_
timestamp 1
transform 1 0 20608 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1
transform 1 0 17572 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _1633_
timestamp 1
transform -1 0 49588 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1634_
timestamp 1
transform -1 0 48852 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1635_
timestamp 1
transform 1 0 42228 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1636_
timestamp 1
transform 1 0 39836 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1637_
timestamp 1
transform 1 0 39652 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1638_
timestamp 1
transform 1 0 45448 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1639_
timestamp 1
transform 1 0 30176 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1640_
timestamp 1
transform 1 0 17020 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1641_
timestamp 1
transform 1 0 12144 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1642_
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1643_
timestamp 1
transform 1 0 14444 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1644_
timestamp 1
transform 1 0 13616 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1645_
timestamp 1
transform 1 0 14904 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1646_
timestamp 1
transform 1 0 12696 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1647_
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1648_
timestamp 1
transform 1 0 22080 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1649_
timestamp 1
transform 1 0 36340 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1650_
timestamp 1
transform 1 0 38180 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1651_
timestamp 1
transform 1 0 36156 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1652_
timestamp 1
transform 1 0 33856 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1653_
timestamp 1
transform 1 0 33488 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1654_
timestamp 1
transform 1 0 34316 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1655_
timestamp 1
transform -1 0 34316 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1656_
timestamp 1
transform 1 0 31188 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1657_
timestamp 1
transform -1 0 33856 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1658_
timestamp 1
transform 1 0 30176 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1659_
timestamp 1
transform 1 0 28428 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1660_
timestamp 1
transform 1 0 26956 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1661_
timestamp 1
transform 1 0 26956 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1662_
timestamp 1
transform 1 0 27324 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1663_
timestamp 1
transform -1 0 31740 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1664_
timestamp 1
transform 1 0 29532 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1665_
timestamp 1
transform -1 0 33948 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1666_
timestamp 1
transform -1 0 34316 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1667_
timestamp 1
transform -1 0 56120 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1668_
timestamp 1
transform 1 0 24564 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1669_
timestamp 1
transform 1 0 28060 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1670_
timestamp 1
transform 1 0 29440 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1671_
timestamp 1
transform 1 0 29716 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1672_
timestamp 1
transform 1 0 26496 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1673_
timestamp 1
transform 1 0 26588 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1674_
timestamp 1
transform 1 0 28060 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1675_
timestamp 1
transform 1 0 29532 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1676_
timestamp 1
transform 1 0 15640 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1677_
timestamp 1
transform 1 0 10396 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1678_
timestamp 1
transform 1 0 9476 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1679_
timestamp 1
transform 1 0 12696 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1680_
timestamp 1
transform 1 0 8556 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1681_
timestamp 1
transform 1 0 7912 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1682_
timestamp 1
transform 1 0 9016 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1683_
timestamp 1
transform 1 0 9476 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1684_
timestamp 1
transform 1 0 12236 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1685_
timestamp 1
transform -1 0 14260 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1686_
timestamp 1
transform -1 0 15456 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1687_
timestamp 1
transform 1 0 14444 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1688_
timestamp 1
transform 1 0 11592 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1689_
timestamp 1
transform -1 0 12052 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1690_
timestamp 1
transform 1 0 8740 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1691_
timestamp 1
transform 1 0 7728 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1692_
timestamp 1
transform -1 0 14812 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1693_
timestamp 1
transform 1 0 13064 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1694_
timestamp 1
transform 1 0 9936 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1695_
timestamp 1
transform -1 0 10212 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1696_
timestamp 1
transform 1 0 8924 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1697_
timestamp 1
transform 1 0 9568 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1698_
timestamp 1
transform 1 0 12052 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1699_
timestamp 1
transform 1 0 12880 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1700_
timestamp 1
transform 1 0 16652 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1701_
timestamp 1
transform 1 0 15824 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1702_
timestamp 1
transform 1 0 14720 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1703_
timestamp 1
transform 1 0 17112 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1704_
timestamp 1
transform 1 0 17664 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1705_
timestamp 1
transform -1 0 20792 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1706_
timestamp 1
transform 1 0 20516 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1707_
timestamp 1
transform -1 0 22540 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1708_
timestamp 1
transform 1 0 18216 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1709_
timestamp 1
transform -1 0 23644 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1710_
timestamp 1
transform 1 0 19228 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1711_
timestamp 1
transform 1 0 19780 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1712_
timestamp 1
transform 1 0 17296 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1713_
timestamp 1
transform 1 0 16652 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1714_
timestamp 1
transform 1 0 15548 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1715_
timestamp 1
transform 1 0 34224 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1716_
timestamp 1
transform 1 0 35972 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1717_
timestamp 1
transform -1 0 39100 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1718_
timestamp 1
transform -1 0 41032 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1719_
timestamp 1
transform -1 0 42320 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1720_
timestamp 1
transform -1 0 42688 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1721_
timestamp 1
transform 1 0 39008 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1722_
timestamp 1
transform 1 0 37444 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1723_
timestamp 1
transform 1 0 44988 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1724_
timestamp 1
transform 1 0 46920 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1725_
timestamp 1
transform 1 0 48024 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1726_
timestamp 1
transform 1 0 47748 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1727_
timestamp 1
transform 1 0 45540 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1728_
timestamp 1
transform 1 0 43148 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1729_
timestamp 1
transform 1 0 42412 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1730_
timestamp 1
transform -1 0 43424 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1731_
timestamp 1
transform 1 0 7544 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1732_
timestamp 1
transform 1 0 7820 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1733_
timestamp 1
transform 1 0 6992 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1734_
timestamp 1
transform 1 0 10120 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1
transform 1 0 37996 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1
transform -1 0 44896 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1737_
timestamp 1
transform -1 0 51152 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1
transform 1 0 56488 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1
transform 1 0 37904 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1
transform 1 0 39652 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1
transform 1 0 57132 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1
transform 1 0 39928 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1743_
timestamp 1
transform 1 0 55660 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _1744__239
timestamp 1
transform 1 0 2484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1744_
timestamp 1
transform -1 0 2116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1745__240
timestamp 1
transform 1 0 2116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1745_
timestamp 1
transform -1 0 2116 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1746__241
timestamp 1
transform 1 0 2116 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1746_
timestamp 1
transform 1 0 2116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1747__242
timestamp 1
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1747_
timestamp 1
transform -1 0 2116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1748_
timestamp 1
transform -1 0 2116 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1748__243
timestamp 1
transform 1 0 2116 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1749__244
timestamp 1
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1749_
timestamp 1
transform -1 0 2116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1750_
timestamp 1
transform -1 0 2116 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1750__245
timestamp 1
transform 1 0 2116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1751__246
timestamp 1
transform 1 0 2116 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1751_
timestamp 1
transform -1 0 2116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1752__247
timestamp 1
transform -1 0 2116 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1752_
timestamp 1
transform -1 0 2116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1753__248
timestamp 1
transform 1 0 2116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1753_
timestamp 1
transform -1 0 2116 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1754__249
timestamp 1
transform 1 0 2116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1754_
timestamp 1
transform -1 0 2116 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1755__250
timestamp 1
transform -1 0 2116 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1755_
timestamp 1
transform -1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1756__251
timestamp 1
transform 1 0 2116 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1756_
timestamp 1
transform -1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1757_
timestamp 1
transform -1 0 2116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1757__252
timestamp 1
transform -1 0 2116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1758__253
timestamp 1
transform -1 0 2116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1758_
timestamp 1
transform -1 0 2116 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1759__254
timestamp 1
transform 1 0 2116 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1759_
timestamp 1
transform -1 0 2116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1760_
timestamp 1
transform -1 0 2116 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1760__255
timestamp 1
transform -1 0 2116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1761__256
timestamp 1
transform 1 0 2116 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1761_
timestamp 1
transform -1 0 2116 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1762__189
timestamp 1
transform 1 0 40296 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1762_
timestamp 1
transform -1 0 40572 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1763__190
timestamp 1
transform -1 0 73876 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1763_
timestamp 1
transform -1 0 73140 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1764__191
timestamp 1
transform -1 0 55752 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1764_
timestamp 1
transform -1 0 55476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1765__192
timestamp 1
transform -1 0 51980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1765_
timestamp 1
transform -1 0 51704 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1766__193
timestamp 1
transform -1 0 41676 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1766_
timestamp 1
transform -1 0 41400 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1767_
timestamp 1
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1767__194
timestamp 1
transform 1 0 68080 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1768__195
timestamp 1
transform -1 0 59064 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1768_
timestamp 1
transform -1 0 58788 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1769_
timestamp 1
transform 1 0 48760 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1769__196
timestamp 1
transform -1 0 49036 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1770__197
timestamp 1
transform -1 0 59708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1770_
timestamp 1
transform -1 0 59432 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1771__198
timestamp 1
transform -1 0 60996 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1771_
timestamp 1
transform -1 0 60168 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1772__199
timestamp 1
transform -1 0 46460 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1772_
timestamp 1
transform -1 0 45908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1773__200
timestamp 1
transform -1 0 56396 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1773_
timestamp 1
transform -1 0 56120 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1774__201
timestamp 1
transform -1 0 54464 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1774_
timestamp 1
transform -1 0 54188 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1775__202
timestamp 1
transform -1 0 57132 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1775_
timestamp 1
transform -1 0 56856 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1776_
timestamp 1
transform -1 0 60720 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1776__203
timestamp 1
transform 1 0 60444 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1777__204
timestamp 1
transform -1 0 51336 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1777_
timestamp 1
transform -1 0 51060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1778__257
timestamp 1
transform 1 0 2484 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1778_
timestamp 1
transform -1 0 2116 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1779__258
timestamp 1
transform 1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1779_
timestamp 1
transform -1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1780_
timestamp 1
transform -1 0 2116 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1780__259
timestamp 1
transform 1 0 2116 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1781__260
timestamp 1
transform -1 0 2116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1781_
timestamp 1
transform 1 0 2116 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1782_
timestamp 1
transform -1 0 43148 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1782__205
timestamp 1
transform 1 0 42872 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1783__206
timestamp 1
transform -1 0 42320 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1783_
timestamp 1
transform -1 0 42044 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1784__207
timestamp 1
transform -1 0 71300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1784_
timestamp 1
transform -1 0 71024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1785__208
timestamp 1
transform -1 0 47472 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1785_
timestamp 1
transform -1 0 47196 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1786__209
timestamp 1
transform -1 0 67436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1786_
timestamp 1
transform -1 0 67160 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1787_
timestamp 1
transform -1 0 53084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1787__210
timestamp 1
transform 1 0 52716 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1788_
timestamp 1
transform -1 0 72312 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1788__211
timestamp 1
transform 1 0 72036 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1789__212
timestamp 1
transform -1 0 64860 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1789_
timestamp 1
transform -1 0 64584 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1790__213
timestamp 1
transform 1 0 40572 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1790_
timestamp 1
transform -1 0 40940 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1791__214
timestamp 1
transform -1 0 71944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1791_
timestamp 1
transform -1 0 71668 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1792_
timestamp 1
transform 1 0 60996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1792__215
timestamp 1
transform -1 0 61272 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1793_
timestamp 1
transform 1 0 42412 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1793__216
timestamp 1
transform 1 0 42320 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1794_
timestamp 1
transform 1 0 44988 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1794__217
timestamp 1
transform 1 0 44436 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1795__218
timestamp 1
transform -1 0 52624 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1795_
timestamp 1
transform -1 0 52348 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1796__219
timestamp 1
transform -1 0 70012 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1796_
timestamp 1
transform -1 0 69736 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1797__220
timestamp 1
transform -1 0 62192 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1797_
timestamp 1
transform -1 0 61916 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1798__221
timestamp 1
transform -1 0 62928 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1798_
timestamp 1
transform -1 0 62652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1799_
timestamp 1
transform 1 0 63020 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1799__222
timestamp 1
transform 1 0 62928 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1800_
timestamp 1
transform -1 0 44436 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1801__223
timestamp 1
transform -1 0 64216 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1801_
timestamp 1
transform -1 0 63940 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1802_
timestamp 1
transform -1 0 46184 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1803_
timestamp 1
transform -1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1804__224
timestamp 1
transform -1 0 49956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1804_
timestamp 1
transform -1 0 49680 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1805__225
timestamp 1
transform -1 0 68080 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1805_
timestamp 1
transform -1 0 67804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1806_
timestamp 1
transform 1 0 53268 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1806__226
timestamp 1
transform -1 0 53544 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1807_
timestamp 1
transform -1 0 58236 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1807__227
timestamp 1
transform 1 0 57868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1808_
timestamp 1
transform -1 0 47932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1808__228
timestamp 1
transform 1 0 47564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1809__229
timestamp 1
transform -1 0 48760 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1809_
timestamp 1
transform -1 0 48484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1810__230
timestamp 1
transform -1 0 65504 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1810_
timestamp 1
transform -1 0 65228 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1811_
timestamp 1
transform -1 0 49036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1812_
timestamp 1
transform -1 0 46460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1813_
timestamp 1
transform -1 0 78016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1814__231
timestamp 1
transform -1 0 66792 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1814_
timestamp 1
transform -1 0 66516 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1815_
timestamp 1
transform -1 0 78108 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1816_
timestamp 1
transform -1 0 78108 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1817_
timestamp 1
transform -1 0 77832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1818__232
timestamp 1
transform -1 0 73600 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1818_
timestamp 1
transform -1 0 72772 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1819_
timestamp 1
transform -1 0 78108 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1820_
timestamp 1
transform -1 0 47104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1821_
timestamp 1
transform -1 0 72956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1822_
timestamp 1
transform 1 0 51152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1823_
timestamp 1
transform -1 0 61824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1824__233
timestamp 1
transform -1 0 70656 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1824_
timestamp 1
transform -1 0 70380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1825_
timestamp 1
transform -1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1826_
timestamp 1
transform 1 0 68540 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1827__234
timestamp 1
transform -1 0 55108 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1827_
timestamp 1
transform -1 0 54832 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1828_
timestamp 1
transform -1 0 63756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1829_
timestamp 1
transform -1 0 45816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1830__235
timestamp 1
transform -1 0 50692 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1830_
timestamp 1
transform -1 0 50416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1831_
timestamp 1
transform -1 0 49680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1832__236
timestamp 1
transform -1 0 57776 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1832_
timestamp 1
transform -1 0 57500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1833_
timestamp 1
transform -1 0 63296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1834__237
timestamp 1
transform -1 0 69368 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1834_
timestamp 1
transform -1 0 69092 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1835_
timestamp 1
transform -1 0 64400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1836_
timestamp 1
transform -1 0 76636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1837_
timestamp 1
transform -1 0 78108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1838_
timestamp 1
transform -1 0 62468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1839__238
timestamp 1
transform -1 0 66148 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1839_
timestamp 1
transform -1 0 65872 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1840_
timestamp 1
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__D
timestamp 1
transform 1 0 65964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A
timestamp 1
transform 1 0 59248 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__C
timestamp 1
transform 1 0 59432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1
transform 1 0 28428 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B
timestamp 1
transform -1 0 54096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__C
timestamp 1
transform -1 0 57776 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A
timestamp 1
transform 1 0 29808 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1
transform 1 0 29072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A1
timestamp 1
transform 1 0 44528 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A1
timestamp 1
transform 1 0 48944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A1
timestamp 1
transform 1 0 48300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A1
timestamp 1
transform -1 0 47840 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A1
timestamp 1
transform -1 0 47196 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A1
timestamp 1
transform -1 0 30360 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A1
timestamp 1
transform 1 0 48576 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A1
timestamp 1
transform 1 0 49220 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__B1
timestamp 1
transform 1 0 48392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A1
timestamp 1
transform -1 0 42320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A1
timestamp 1
transform -1 0 50048 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1
transform -1 0 47748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1
transform 1 0 50140 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A2
timestamp 1
transform 1 0 43608 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__B1
timestamp 1
transform 1 0 42964 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B1
timestamp 1
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__B1
timestamp 1
transform -1 0 42964 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__C1
timestamp 1
transform 1 0 49312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__C1
timestamp 1
transform 1 0 54188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B1
timestamp 1
transform 1 0 39468 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B1
timestamp 1
transform 1 0 42504 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__B1
timestamp 1
transform 1 0 54648 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__C1
timestamp 1
transform 1 0 53636 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__B1
timestamp 1
transform 1 0 54924 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__C1
timestamp 1
transform -1 0 44068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__C1
timestamp 1
transform 1 0 53268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__B1
timestamp 1
transform -1 0 53176 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__C1
timestamp 1
transform 1 0 51980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A2
timestamp 1
transform 1 0 35328 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__C1
timestamp 1
transform 1 0 51796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A2
timestamp 1
transform 1 0 35052 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A2
timestamp 1
transform -1 0 53544 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__C1
timestamp 1
transform 1 0 44252 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A2
timestamp 1
transform 1 0 47564 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A2
timestamp 1
transform 1 0 35972 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__B1
timestamp 1
transform 1 0 36156 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A2
timestamp 1
transform 1 0 36432 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__C1
timestamp 1
transform 1 0 36248 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__C1
timestamp 1
transform 1 0 46184 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A2
timestamp 1
transform 1 0 46368 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__B1
timestamp 1
transform 1 0 45632 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A2
timestamp 1
transform -1 0 47472 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__B1
timestamp 1
transform 1 0 44804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__B1
timestamp 1
transform 1 0 48208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__B
timestamp 1
transform -1 0 46460 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__B1
timestamp 1
transform 1 0 46000 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A2
timestamp 1
transform -1 0 37996 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__B1
timestamp 1
transform 1 0 47840 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__S
timestamp 1
transform 1 0 47288 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__S
timestamp 1
transform 1 0 47288 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__S
timestamp 1
transform 1 0 43424 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__S
timestamp 1
transform 1 0 41308 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__S
timestamp 1
transform 1 0 41216 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__S
timestamp 1
transform 1 0 45724 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A1
timestamp 1
transform -1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__A1
timestamp 1
transform -1 0 24012 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__A0
timestamp 1
transform 1 0 30544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__A1
timestamp 1
transform 1 0 28060 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__A1
timestamp 1
transform -1 0 29716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__A1
timestamp 1
transform -1 0 27048 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__A1
timestamp 1
transform -1 0 29532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__B1
timestamp 1
transform -1 0 29992 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__A2
timestamp 1
transform 1 0 37812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__B1
timestamp 1
transform 1 0 36432 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A2
timestamp 1
transform 1 0 37168 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__B1
timestamp 1
transform 1 0 37352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__A2
timestamp 1
transform 1 0 36524 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__B1
timestamp 1
transform 1 0 36708 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A2
timestamp 1
transform 1 0 40756 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__B1
timestamp 1
transform 1 0 41492 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__A2
timestamp 1
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__B1
timestamp 1
transform 1 0 36984 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__A2
timestamp 1
transform 1 0 38272 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__B1
timestamp 1
transform 1 0 38456 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A2
timestamp 1
transform 1 0 38088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__B1
timestamp 1
transform 1 0 38640 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A2
timestamp 1
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__B1
timestamp 1
transform 1 0 40296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__A2
timestamp 1
transform 1 0 39008 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__A2
timestamp 1
transform -1 0 45540 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__B1
timestamp 1
transform -1 0 45172 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__A2
timestamp 1
transform 1 0 42688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__B1
timestamp 1
transform 1 0 42872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__A2
timestamp 1
transform 1 0 43240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__B1
timestamp 1
transform 1 0 44068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__A2
timestamp 1
transform 1 0 43608 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__B1
timestamp 1
transform 1 0 43424 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__A2
timestamp 1
transform -1 0 43516 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__B1
timestamp 1
transform 1 0 42412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__A2
timestamp 1
transform -1 0 44620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__B1
timestamp 1
transform 1 0 45356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__A1
timestamp 1
transform 1 0 45356 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__A2
timestamp 1
transform 1 0 45724 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__B1
timestamp 1
transform 1 0 45540 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__A2
timestamp 1
transform -1 0 43056 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__B1
timestamp 1
transform 1 0 43792 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__A2
timestamp 1
transform 1 0 43240 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__A2
timestamp 1
transform -1 0 51244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__B1
timestamp 1
transform 1 0 49588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__A1
timestamp 1
transform 1 0 48576 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__A2
timestamp 1
transform 1 0 48944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__B1
timestamp 1
transform 1 0 48760 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__A1
timestamp 1
transform -1 0 50048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__A2
timestamp 1
transform -1 0 49864 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__B1
timestamp 1
transform 1 0 50140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__A2
timestamp 1
transform 1 0 50140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__B1
timestamp 1
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A2
timestamp 1
transform 1 0 50140 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__B1
timestamp 1
transform 1 0 49772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__A2
timestamp 1
transform 1 0 50324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__B1
timestamp 1
transform 1 0 50140 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__A2
timestamp 1
transform -1 0 51796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__B1
timestamp 1
transform -1 0 50600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__A2
timestamp 1
transform 1 0 51428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__B1
timestamp 1
transform 1 0 50692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__B
timestamp 1
transform 1 0 49496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__A2
timestamp 1
transform 1 0 48484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__B1
timestamp 1
transform 1 0 48300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__A2
timestamp 1
transform -1 0 51704 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__B1
timestamp 1
transform 1 0 50508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__A2
timestamp 1
transform 1 0 49128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__B1
timestamp 1
transform 1 0 48944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__A2
timestamp 1
transform 1 0 49956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__B1
timestamp 1
transform 1 0 49772 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__A2
timestamp 1
transform -1 0 50968 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__B1
timestamp 1
transform 1 0 49772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__B2
timestamp 1
transform -1 0 49772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__A2
timestamp 1
transform 1 0 49496 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__B1
timestamp 1
transform 1 0 49680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__A2
timestamp 1
transform -1 0 51888 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__A1
timestamp 1
transform 1 0 46736 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__A2
timestamp 1
transform 1 0 47104 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__B1
timestamp 1
transform 1 0 44896 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__C1
timestamp 1
transform 1 0 44712 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__B1
timestamp 1
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__A2
timestamp 1
transform 1 0 55568 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__A2
timestamp 1
transform 1 0 35604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__B1
timestamp 1
transform 1 0 35788 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__A2
timestamp 1
transform 1 0 37444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__B1
timestamp 1
transform 1 0 37628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__A2
timestamp 1
transform 1 0 35512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__B1
timestamp 1
transform 1 0 36156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__A2
timestamp 1
transform 1 0 36616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__B1
timestamp 1
transform -1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__A2
timestamp 1
transform 1 0 35788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__B1
timestamp 1
transform -1 0 36156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A2
timestamp 1
transform -1 0 36708 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__B1
timestamp 1
transform -1 0 37168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A2
timestamp 1
transform 1 0 39376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__B1
timestamp 1
transform 1 0 39376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__C1
timestamp 1
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A2
timestamp 1
transform 1 0 37352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__B1
timestamp 1
transform 1 0 37536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__A2
timestamp 1
transform 1 0 38732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__A2
timestamp 1
transform 1 0 38180 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__B1
timestamp 1
transform 1 0 38180 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__A2
timestamp 1
transform -1 0 36156 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__B1
timestamp 1
transform -1 0 36340 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__A2
timestamp 1
transform 1 0 35512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__B1
timestamp 1
transform 1 0 35696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__B1
timestamp 1
transform 1 0 39928 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__A2
timestamp 1
transform 1 0 39192 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__B1
timestamp 1
transform 1 0 40112 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__B1
timestamp 1
transform -1 0 40756 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__A2
timestamp 1
transform 1 0 36800 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__B1
timestamp 1
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__A2
timestamp 1
transform 1 0 37904 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__B1
timestamp 1
transform 1 0 38088 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__A2
timestamp 1
transform -1 0 36064 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__B1
timestamp 1
transform -1 0 36248 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__A2
timestamp 1
transform 1 0 36892 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__B
timestamp 1
transform 1 0 40296 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__A2
timestamp 1
transform 1 0 49772 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__B1
timestamp 1
transform 1 0 49588 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__A2
timestamp 1
transform 1 0 50416 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__B1
timestamp 1
transform 1 0 50232 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__A2
timestamp 1
transform 1 0 50876 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__B1
timestamp 1
transform 1 0 50692 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__A2
timestamp 1
transform 1 0 49036 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__B1
timestamp 1
transform 1 0 48852 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__A2
timestamp 1
transform 1 0 49588 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__B1
timestamp 1
transform 1 0 49496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__B2
timestamp 1
transform 1 0 49128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__A2
timestamp 1
transform 1 0 50416 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__B1
timestamp 1
transform 1 0 50232 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__A1
timestamp 1
transform 1 0 49312 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__A2
timestamp 1
transform 1 0 48208 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__B1
timestamp 1
transform 1 0 48024 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__A2
timestamp 1
transform 1 0 50324 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__B1
timestamp 1
transform 1 0 50140 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__A2
timestamp 1
transform -1 0 56212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__B
timestamp 1
transform -1 0 36708 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__A2
timestamp 1
transform 1 0 36708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__B1
timestamp 1
transform 1 0 36892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__B
timestamp 1
transform 1 0 41400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__A2
timestamp 1
transform 1 0 37904 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__B1
timestamp 1
transform 1 0 38088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__A2
timestamp 1
transform 1 0 38824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__B1
timestamp 1
transform 1 0 38916 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__A2
timestamp 1
transform 1 0 42872 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__B1
timestamp 1
transform 1 0 43056 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__A2
timestamp 1
transform 1 0 40480 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__B1
timestamp 1
transform 1 0 40664 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__A2
timestamp 1
transform 1 0 40848 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__A2
timestamp 1
transform 1 0 36892 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__B1
timestamp 1
transform 1 0 37076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__A2
timestamp 1
transform 1 0 37536 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__A2
timestamp 1
transform 1 0 40664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__RESET_B
timestamp 1
transform 1 0 19688 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__RESET_B
timestamp 1
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__RESET_B
timestamp 1
transform 1 0 37996 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1509__RESET_B
timestamp 1
transform 1 0 46644 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__SET_B
timestamp 1
transform 1 0 31464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__RESET_B
timestamp 1
transform -1 0 33304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1520__RESET_B
timestamp 1
transform 1 0 32752 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__SET_B
timestamp 1
transform 1 0 30544 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1523__RESET_B
timestamp 1
transform 1 0 35052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1526__RESET_B
timestamp 1
transform 1 0 50324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1531__RESET_B
timestamp 1
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1536__RESET_B
timestamp 1
transform 1 0 31556 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1537__SET_B
timestamp 1
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1540__RESET_B
timestamp 1
transform -1 0 42596 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1544__RESET_B
timestamp 1
transform 1 0 31648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1545__SET_B
timestamp 1
transform 1 0 31004 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1550__RESET_B
timestamp 1
transform 1 0 54188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__RESET_B
timestamp 1
transform 1 0 32200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1553__SET_B
timestamp 1
transform 1 0 31648 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__RESET_B
timestamp 1
transform 1 0 56028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1561__SET_B
timestamp 1
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1566__RESET_B
timestamp 1
transform 1 0 56856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__RESET_B
timestamp 1
transform 1 0 54924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1575__RESET_B
timestamp 1
transform -1 0 56672 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__RESET_B
timestamp 1
transform 1 0 52992 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1588__RESET_B
timestamp 1
transform 1 0 35420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1590__RESET_B
timestamp 1
transform 1 0 54832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1591__RESET_B
timestamp 1
transform -1 0 52256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1596__RESET_B
timestamp 1
transform 1 0 35696 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1598__RESET_B
timestamp 1
transform -1 0 57316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__RESET_B
timestamp 1
transform 1 0 33396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1611__RESET_B
timestamp 1
transform 1 0 36248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1619__RESET_B
timestamp 1
transform -1 0 34500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1628__SET_B
timestamp 1
transform 1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__RESET_B
timestamp 1
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1631__RESET_B
timestamp 1
transform 1 0 22448 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1633__RESET_B
timestamp 1
transform 1 0 49588 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1639__D
timestamp 1
transform -1 0 30176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1639__RESET_B
timestamp 1
transform 1 0 32568 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1653__RESET_B
timestamp 1
transform 1 0 35328 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1657__RESET_B
timestamp 1
transform 1 0 33856 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1669__RESET_B
timestamp 1
transform 1 0 29900 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1672__RESET_B
timestamp 1
transform 1 0 28336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1673__SET_B
timestamp 1
transform 1 0 28520 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1686__RESET_B
timestamp 1
transform -1 0 15640 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1687__RESET_B
timestamp 1
transform 1 0 16284 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1688__RESET_B
timestamp 1
transform 1 0 13708 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1691__RESET_B
timestamp 1
transform 1 0 10304 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1693__RESET_B
timestamp 1
transform 1 0 14904 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1696__RESET_B
timestamp 1
transform 1 0 11500 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1697__RESET_B
timestamp 1
transform 1 0 12236 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1698__RESET_B
timestamp 1
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1699__RESET_B
timestamp 1
transform 1 0 14720 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1700__RESET_B
timestamp 1
transform 1 0 18492 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1701__RESET_B
timestamp 1
transform 1 0 17664 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1702__RESET_B
timestamp 1
transform 1 0 17388 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1703__RESET_B
timestamp 1
transform 1 0 18952 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1704__RESET_B
timestamp 1
transform 1 0 20240 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1705__RESET_B
timestamp 1
transform 1 0 20792 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1707__RESET_B
timestamp 1
transform -1 0 22724 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1708__RESET_B
timestamp 1
transform 1 0 18032 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1709__RESET_B
timestamp 1
transform 1 0 23644 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1710__RESET_B
timestamp 1
transform -1 0 21252 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1711__RESET_B
timestamp 1
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1712__RESET_B
timestamp 1
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1713__RESET_B
timestamp 1
transform 1 0 18492 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1714__RESET_B
timestamp 1
transform 1 0 17756 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1722__RESET_B
timestamp 1
transform 1 0 39836 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1723__RESET_B
timestamp 1
transform 1 0 46828 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1724__RESET_B
timestamp 1
transform 1 0 48760 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1725__RESET_B
timestamp 1
transform 1 0 49864 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1726__RESET_B
timestamp 1
transform 1 0 49588 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1727__RESET_B
timestamp 1
transform 1 0 47564 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1728__RESET_B
timestamp 1
transform -1 0 45540 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1813__A
timestamp 1
transform 1 0 77556 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1815__A
timestamp 1
transform -1 0 77372 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1816__A
timestamp 1
transform 1 0 77648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1817__A
timestamp 1
transform -1 0 77556 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1819__A
timestamp 1
transform -1 0 77832 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1821__A
timestamp 1
transform 1 0 72956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1823__A
timestamp 1
transform -1 0 62008 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1826__A
timestamp 1
transform -1 0 69000 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1828__A
timestamp 1
transform -1 0 63940 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1833__A
timestamp 1
transform -1 0 63480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1835__A
timestamp 1
transform -1 0 64584 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1836__A
timestamp 1
transform -1 0 76360 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1837__A
timestamp 1
transform -1 0 77832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1838__A
timestamp 1
transform -1 0 62652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1
transform 1 0 33948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_wb_clk_i_A
timestamp 1
transform 1 0 23644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_wb_clk_i_A
timestamp 1
transform 1 0 41032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1
transform 1 0 11592 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1
transform 1 0 27692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1
transform 1 0 18584 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1
transform 1 0 13524 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1
transform 1 0 21620 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1
transform 1 0 29348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1
transform 1 0 26864 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1
transform 1 0 34316 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1
transform 1 0 38824 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1
transform -1 0 36708 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1
transform 1 0 44988 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1
transform 1 0 51704 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_wb_clk_i_A
timestamp 1
transform 1 0 53176 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_wb_clk_i_A
timestamp 1
transform 1 0 43240 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_wb_clk_i_A
timestamp 1
transform 1 0 41584 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_wb_clk_i_A
timestamp 1
transform 1 0 45540 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_wb_clk_i_A
timestamp 1
transform 1 0 53176 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_wb_clk_i_A
timestamp 1
transform 1 0 50876 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_wb_clk_i_A
timestamp 1
transform 1 0 53084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_wb_clk_i_A
timestamp 1
transform 1 0 44988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_wb_clk_i_A
timestamp 1
transform -1 0 37076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_wb_clk_i_A
timestamp 1
transform 1 0 38824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_wb_clk_i_A
timestamp 1
transform 1 0 34224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_wb_clk_i_A
timestamp 1
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_wb_clk_i_A
timestamp 1
transform -1 0 30268 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_27_wb_clk_i_A
timestamp 1
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout82_A
timestamp 1
transform 1 0 32660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout83_A
timestamp 1
transform -1 0 31280 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout84_A
timestamp 1
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout85_A
timestamp 1
transform 1 0 46368 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout86_A
timestamp 1
transform -1 0 50876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout87_A
timestamp 1
transform 1 0 51336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout88_A
timestamp 1
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout95_A
timestamp 1
transform 1 0 30636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout96_A
timestamp 1
transform 1 0 30728 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout97_A
timestamp 1
transform 1 0 38180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout98_A
timestamp 1
transform 1 0 44620 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout99_A
timestamp 1
transform 1 0 43332 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout101_A
timestamp 1
transform 1 0 35880 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout102_A
timestamp 1
transform 1 0 34040 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_A
timestamp 1
transform -1 0 40756 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp 1
transform 1 0 38640 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_A
timestamp 1
transform 1 0 33948 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_A
timestamp 1
transform -1 0 29716 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout107_A
timestamp 1
transform 1 0 37444 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout119_A
timestamp 1
transform 1 0 32384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout120_A
timestamp 1
transform 1 0 33120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_A
timestamp 1
transform -1 0 36064 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_A
timestamp 1
transform -1 0 42596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout124_A
timestamp 1
transform 1 0 33672 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout125_A
timestamp 1
transform 1 0 35512 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout127_A
timestamp 1
transform 1 0 44068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout128_A
timestamp 1
transform 1 0 44068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout129_A
timestamp 1
transform 1 0 49496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout130_A
timestamp 1
transform 1 0 52440 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout133_A
timestamp 1
transform -1 0 43976 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout135_A
timestamp 1
transform 1 0 43700 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout139_A
timestamp 1
transform 1 0 32936 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout140_A
timestamp 1
transform 1 0 28152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout141_A
timestamp 1
transform 1 0 31280 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout142_A
timestamp 1
transform -1 0 37812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout143_A
timestamp 1
transform 1 0 29164 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout145_A
timestamp 1
transform 1 0 41032 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout146_A
timestamp 1
transform -1 0 49312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout147_A
timestamp 1
transform 1 0 50232 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout148_A
timestamp 1
transform 1 0 49956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout149_A
timestamp 1
transform 1 0 51336 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout150_A
timestamp 1
transform 1 0 42872 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout153_A
timestamp 1
transform 1 0 58512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout154_A
timestamp 1
transform -1 0 69184 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout157_A
timestamp 1
transform -1 0 18216 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout158_A
timestamp 1
transform -1 0 32016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout159_A
timestamp 1
transform 1 0 32108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout160_A
timestamp 1
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout161_A
timestamp 1
transform 1 0 14628 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout162_A
timestamp 1
transform -1 0 19964 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout163_A
timestamp 1
transform 1 0 18400 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout164_A
timestamp 1
transform 1 0 31096 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout165_A
timestamp 1
transform 1 0 30636 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout166_A
timestamp 1
transform 1 0 31464 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout169_A
timestamp 1
transform 1 0 44620 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout170_A
timestamp 1
transform 1 0 44344 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout171_A
timestamp 1
transform 1 0 44620 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout172_A
timestamp 1
transform 1 0 51244 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout173_A
timestamp 1
transform 1 0 55844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout175_A
timestamp 1
transform 1 0 55292 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout176_A
timestamp 1
transform -1 0 55200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout177_A
timestamp 1
transform 1 0 37720 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout178_A
timestamp 1
transform 1 0 41768 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout179_A
timestamp 1
transform -1 0 37996 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout180_A
timestamp 1
transform -1 0 44804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout181_A
timestamp 1
transform 1 0 44804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout183_A
timestamp 1
transform -1 0 56856 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout184_A
timestamp 1
transform 1 0 55568 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout185_A
timestamp 1
transform 1 0 55108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold122_A
timestamp 1
transform -1 0 58788 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold134_A
timestamp 1
transform -1 0 58052 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1
transform -1 0 1840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1
transform -1 0 1840 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1
transform -1 0 1840 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1
transform -1 0 1840 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1
transform -1 0 51520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1
transform -1 0 52900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1
transform -1 0 59340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1
transform -1 0 54280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1
transform -1 0 56856 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1
transform -1 0 56580 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1
transform -1 0 59984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1
transform -1 0 60628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1
transform -1 0 78568 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1
transform -1 0 70932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1
transform -1 0 74152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1
transform -1 0 77372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1
transform -1 0 61272 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1
transform -1 0 76084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1
transform -1 0 65136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1
transform -1 0 65780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1
transform -1 0 75440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1
transform -1 0 67068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1
transform -1 0 73508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1
transform -1 0 74796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1
transform -1 0 73968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1
transform -1 0 71576 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1
transform -1 0 67712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1
transform -1 0 58696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1
transform -1 0 78200 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1
transform -1 0 69000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1
transform -1 0 52256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1
transform -1 0 69644 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1
transform -1 0 70288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1
transform -1 0 47012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1
transform -1 0 66424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1
transform -1 0 53544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1
transform -1 0 45816 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1
transform -1 0 57500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1
transform -1 0 59156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1
transform -1 0 78292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1
transform -1 0 78108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output45_A
timestamp 1
transform 1 0 77832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output48_A
timestamp 1
transform 1 0 77832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1
transform -1 0 33304 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1
transform -1 0 23644 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1
transform 1 0 41216 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_0_wb_clk_i
timestamp 1
transform 1 0 10580 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_1_wb_clk_i
timestamp 1
transform 1 0 17480 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_2_wb_clk_i
timestamp 1
transform 1 0 27876 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_3_wb_clk_i
timestamp 1
transform 1 0 16376 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_4_wb_clk_i
timestamp 1
transform -1 0 10580 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_5_wb_clk_i
timestamp 1
transform 1 0 12512 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_6_wb_clk_i
timestamp 1
transform 1 0 20608 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_7_wb_clk_i
timestamp 1
transform 1 0 29532 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_8_wb_clk_i
timestamp 1
transform 1 0 27048 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_9_wb_clk_i
timestamp 1
transform 1 0 33304 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_10_wb_clk_i
timestamp 1
transform 1 0 37812 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_11_wb_clk_i
timestamp 1
transform 1 0 35512 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_12_wb_clk_i
timestamp 1
transform 1 0 45080 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_13_wb_clk_i
timestamp 1
transform 1 0 51612 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_14_wb_clk_i
timestamp 1
transform 1 0 53360 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_15_wb_clk_i
timestamp 1
transform 1 0 42228 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_16_wb_clk_i
timestamp 1
transform 1 0 40572 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_17_wb_clk_i
timestamp 1
transform 1 0 45724 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_18_wb_clk_i
timestamp 1
transform 1 0 53360 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_19_wb_clk_i
timestamp 1
transform 1 0 51060 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_20_wb_clk_i
timestamp 1
transform 1 0 53268 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_21_wb_clk_i
timestamp 1
transform 1 0 45172 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_22_wb_clk_i
timestamp 1
transform 1 0 35880 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_23_wb_clk_i
timestamp 1
transform 1 0 37812 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_24_wb_clk_i
timestamp 1
transform -1 0 33580 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_25_wb_clk_i
timestamp 1
transform 1 0 25576 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_26_wb_clk_i
timestamp 1
transform 1 0 30268 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_27_wb_clk_i
timestamp 1
transform 1 0 17112 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout82
timestamp 1
transform -1 0 32660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout83
timestamp 1
transform 1 0 31280 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout84
timestamp 1
transform -1 0 32016 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout85
timestamp 1
transform -1 0 46920 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout86
timestamp 1
transform -1 0 51244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout87
timestamp 1
transform 1 0 50968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout88
timestamp 1
transform 1 0 42412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout89
timestamp 1
transform 1 0 32936 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout90
timestamp 1
transform 1 0 28428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout91
timestamp 1
transform -1 0 29808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout92
timestamp 1
transform 1 0 34224 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 1
transform 1 0 44988 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout94
timestamp 1
transform -1 0 42228 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout95
timestamp 1
transform -1 0 31188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout96
timestamp 1
transform -1 0 30728 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout97
timestamp 1
transform -1 0 39284 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout98
timestamp 1
transform 1 0 44068 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout99
timestamp 1
transform 1 0 43516 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout100
timestamp 1
transform -1 0 30820 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout101
timestamp 1
transform -1 0 36524 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout102
timestamp 1
transform 1 0 32292 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout103
timestamp 1
transform -1 0 40572 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout104
timestamp 1
transform 1 0 38272 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout105
timestamp 1
transform 1 0 33028 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout106
timestamp 1
transform 1 0 29716 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout107
timestamp 1
transform 1 0 37076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout108
timestamp 1
transform 1 0 33580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout109
timestamp 1
transform -1 0 49496 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 1
transform -1 0 45356 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout111
timestamp 1
transform 1 0 55936 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout112
timestamp 1
transform -1 0 51152 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout113
timestamp 1
transform 1 0 50968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout114
timestamp 1
transform 1 0 53544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 1
transform -1 0 43792 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout116
timestamp 1
transform 1 0 43516 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout117
timestamp 1
transform 1 0 37260 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout118
timestamp 1
transform -1 0 43792 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout119
timestamp 1
transform 1 0 32016 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout120
timestamp 1
transform 1 0 33304 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout121
timestamp 1
transform -1 0 37076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout122
timestamp 1
transform 1 0 42412 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout123
timestamp 1
transform -1 0 29440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout124
timestamp 1
transform 1 0 33304 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout125
timestamp 1
transform 1 0 36616 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout126
timestamp 1
transform 1 0 31648 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout127
timestamp 1
transform 1 0 43332 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout128
timestamp 1
transform 1 0 43700 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout129
timestamp 1
transform 1 0 49680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout130
timestamp 1
transform 1 0 52716 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout131
timestamp 1
transform 1 0 52164 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout132
timestamp 1
transform -1 0 50048 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout133
timestamp 1
transform -1 0 43424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout134
timestamp 1
transform 1 0 43516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout135
timestamp 1
transform -1 0 43700 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout136
timestamp 1
transform -1 0 35052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout137
timestamp 1
transform 1 0 37260 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout138
timestamp 1
transform 1 0 37260 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout139
timestamp 1
transform 1 0 33120 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout140
timestamp 1
transform -1 0 28152 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout141
timestamp 1
transform 1 0 30728 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout142
timestamp 1
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout143
timestamp 1
transform -1 0 29164 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout144
timestamp 1
transform 1 0 42044 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout145
timestamp 1
transform 1 0 41952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout146
timestamp 1
transform 1 0 49312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout147
timestamp 1
transform 1 0 50416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout148
timestamp 1
transform 1 0 49588 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout149
timestamp 1
transform 1 0 51520 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout150
timestamp 1
transform 1 0 43056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout151
timestamp 1
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout152
timestamp 1
transform 1 0 23644 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout153
timestamp 1
transform -1 0 58512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout154
timestamp 1
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout155
timestamp 1
transform 1 0 73324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout156
timestamp 1
transform -1 0 14628 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout157
timestamp 1
transform 1 0 17480 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout158
timestamp 1
transform 1 0 32016 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout159
timestamp 1
transform 1 0 32292 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout160
timestamp 1
transform 1 0 31464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout161
timestamp 1
transform -1 0 14628 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout162
timestamp 1
transform 1 0 19228 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout163
timestamp 1
transform -1 0 18400 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout164
timestamp 1
transform 1 0 30176 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout165
timestamp 1
transform 1 0 30084 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout166
timestamp 1
transform -1 0 31464 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout167
timestamp 1
transform -1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout168
timestamp 1
transform 1 0 44896 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout169
timestamp 1
transform -1 0 44620 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout170
timestamp 1
transform 1 0 44528 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout171
timestamp 1
transform -1 0 43884 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout172
timestamp 1
transform -1 0 50784 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout173
timestamp 1
transform 1 0 55292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout174
timestamp 1
transform 1 0 56028 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout175
timestamp 1
transform 1 0 55476 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout176
timestamp 1
transform 1 0 54648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout177
timestamp 1
transform -1 0 37720 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout178
timestamp 1
transform -1 0 41768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout179
timestamp 1
transform 1 0 37260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout180
timestamp 1
transform -1 0 44252 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout181
timestamp 1
transform -1 0 44620 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout182
timestamp 1
transform 1 0 56672 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout183
timestamp 1
transform -1 0 56672 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout184
timestamp 1
transform 1 0 55752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout185
timestamp 1
transform 1 0 54740 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout186
timestamp 1
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout187
timestamp 1
transform -1 0 24196 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout188
timestamp 1
transform 1 0 27876 0 -1 11968
box -38 -48 958 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636968456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636968456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1636968456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1636968456
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_337
timestamp 1
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_345
timestamp 1
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_350
timestamp 1636968456
transform 1 0 33304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_362
timestamp 1
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1636968456
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1636968456
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_393
timestamp 1
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_419
timestamp 1
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_421
timestamp 1
transform 1 0 39836 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_432
timestamp 1636968456
transform 1 0 40848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_444
timestamp 1
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_449
timestamp 1
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_455
timestamp 1
transform 1 0 42964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_499
timestamp 1
transform 1 0 47012 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_505
timestamp 1
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_511
timestamp 1
transform 1 0 48116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_518
timestamp 1
transform 1 0 48760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_525
timestamp 1
transform 1 0 49404 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_541
timestamp 1
transform 1 0 50876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_548
timestamp 1
transform 1 0 51520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_553
timestamp 1
transform 1 0 51980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_559
timestamp 1
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_566
timestamp 1
transform 1 0 53176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_580
timestamp 1
transform 1 0 54464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_587
timestamp 1
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_592
timestamp 1
transform 1 0 55568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_636
timestamp 1
transform 1 0 59616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_643
timestamp 1
transform 1 0 60260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_650
timestamp 1
transform 1 0 60904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_657
timestamp 1
transform 1 0 61548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_665
timestamp 1
transform 1 0 62284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_673
timestamp 1
transform 1 0 63020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_679
timestamp 1
transform 1 0 63572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_686
timestamp 1
transform 1 0 64216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_693
timestamp 1
transform 1 0 64860 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_699
timestamp 1
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_706
timestamp 1
transform 1 0 66056 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_713
timestamp 1
transform 1 0 66700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_720
timestamp 1
transform 1 0 67344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_727
timestamp 1
transform 1 0 67988 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_729
timestamp 1
transform 1 0 68172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_735
timestamp 1
transform 1 0 68724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_741
timestamp 1
transform 1 0 69276 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_748
timestamp 1
transform 1 0 69920 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_755
timestamp 1
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_762
timestamp 1
transform 1 0 71208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_769
timestamp 1
transform 1 0 71852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_779
timestamp 1
transform 1 0 72772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_797
timestamp 1
transform 1 0 74428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_804
timestamp 1
transform 1 0 75072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_811
timestamp 1
transform 1 0 75716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_818
timestamp 1
transform 1 0 76360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_826
timestamp 1
transform 1 0 77096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_832
timestamp 1
transform 1 0 77648 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_841
timestamp 1
transform 1 0 78476 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636968456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1636968456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1636968456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1636968456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_329
timestamp 1
transform 1 0 31372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_333
timestamp 1
transform 1 0 31740 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_337
timestamp 1
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_342
timestamp 1636968456
transform 1 0 32568 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_354
timestamp 1636968456
transform 1 0 33672 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_366
timestamp 1
transform 1 0 34776 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_393
timestamp 1
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_399
timestamp 1
transform 1 0 37812 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_420
timestamp 1
transform 1 0 39744 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_446
timestamp 1
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_449
timestamp 1
transform 1 0 42412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_457
timestamp 1
transform 1 0 43148 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_482
timestamp 1
transform 1 0 45448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_486
timestamp 1
transform 1 0 45816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_493
timestamp 1
transform 1 0 46460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_500
timestamp 1
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_508
timestamp 1
transform 1 0 47840 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_516
timestamp 1
transform 1 0 48576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_521
timestamp 1
transform 1 0 49036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_550
timestamp 1
transform 1 0 51704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_558
timestamp 1
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_561
timestamp 1
transform 1 0 52716 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_606
timestamp 1
transform 1 0 56856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_610
timestamp 1
transform 1 0 57224 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_613
timestamp 1
transform 1 0 57500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_632
timestamp 1
transform 1 0 59248 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_645
timestamp 1636968456
transform 1 0 60444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_662
timestamp 1
transform 1 0 62008 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_669
timestamp 1
transform 1 0 62652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_683
timestamp 1
transform 1 0 63940 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_690
timestamp 1636968456
transform 1 0 64584 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_702
timestamp 1
transform 1 0 65688 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_713
timestamp 1636968456
transform 1 0 66700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_725
timestamp 1
transform 1 0 67804 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_740
timestamp 1636968456
transform 1 0 69184 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_752
timestamp 1
transform 1 0 70288 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_758
timestamp 1
transform 1 0 70840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_762
timestamp 1
transform 1 0 71208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_770
timestamp 1
transform 1 0 71944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_783
timestamp 1
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_789
timestamp 1
transform 1 0 73692 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_799
timestamp 1636968456
transform 1 0 74612 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_811
timestamp 1
transform 1 0 75716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_815
timestamp 1
transform 1 0 76084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_821
timestamp 1
transform 1 0 76636 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_829
timestamp 1
transform 1 0 77372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_841
timestamp 1
transform 1 0 78476 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1636968456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_309
timestamp 1
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_313
timestamp 1
transform 1 0 29900 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_344
timestamp 1636968456
transform 1 0 32752 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_356
timestamp 1
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1636968456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1636968456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1636968456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_401
timestamp 1
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1636968456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_433
timestamp 1
transform 1 0 40940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_455
timestamp 1
transform 1 0 42964 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_465
timestamp 1
transform 1 0 43884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 1
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_497
timestamp 1636968456
transform 1 0 46828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_509
timestamp 1636968456
transform 1 0 47932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_521
timestamp 1
transform 1 0 49036 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_529
timestamp 1
transform 1 0 49772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_533
timestamp 1
transform 1 0 50140 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_547
timestamp 1636968456
transform 1 0 51428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_559
timestamp 1636968456
transform 1 0 52532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_571
timestamp 1636968456
transform 1 0 53636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_583
timestamp 1
transform 1 0 54740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_587
timestamp 1
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_606
timestamp 1
transform 1 0 56856 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_636
timestamp 1
transform 1 0 59616 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_645
timestamp 1636968456
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_657
timestamp 1636968456
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_669
timestamp 1636968456
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_681
timestamp 1636968456
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_693
timestamp 1
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_699
timestamp 1
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_701
timestamp 1636968456
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_713
timestamp 1636968456
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_725
timestamp 1636968456
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_737
timestamp 1636968456
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_749
timestamp 1
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_755
timestamp 1
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_757
timestamp 1636968456
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_769
timestamp 1
transform 1 0 71852 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_783
timestamp 1636968456
transform 1 0 73140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_795
timestamp 1636968456
transform 1 0 74244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_807
timestamp 1
transform 1 0 75348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_811
timestamp 1
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_813
timestamp 1636968456
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_825
timestamp 1
transform 1 0 77004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_833
timestamp 1
transform 1 0 77740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_838
timestamp 1
transform 1 0 78200 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1636968456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1636968456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1636968456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1636968456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1636968456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1636968456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_329
timestamp 1
transform 1 0 31372 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1636968456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1636968456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_388
timestamp 1
transform 1 0 36800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_401
timestamp 1636968456
transform 1 0 37996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_413
timestamp 1636968456
transform 1 0 39100 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_425
timestamp 1
transform 1 0 40204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_449
timestamp 1
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_465
timestamp 1
transform 1 0 43884 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_475
timestamp 1
transform 1 0 44804 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_485
timestamp 1636968456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_497
timestamp 1
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 1
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_525
timestamp 1636968456
transform 1 0 49404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_537
timestamp 1636968456
transform 1 0 50508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_549
timestamp 1
transform 1 0 51612 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_557
timestamp 1
transform 1 0 52348 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_561
timestamp 1636968456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_573
timestamp 1636968456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_585
timestamp 1636968456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_597
timestamp 1
transform 1 0 56028 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_603
timestamp 1636968456
transform 1 0 56580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_617
timestamp 1
transform 1 0 57868 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_626
timestamp 1636968456
transform 1 0 58696 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_638
timestamp 1636968456
transform 1 0 59800 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_650
timestamp 1636968456
transform 1 0 60904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_662
timestamp 1
transform 1 0 62008 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_670
timestamp 1
transform 1 0 62744 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_673
timestamp 1636968456
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_685
timestamp 1636968456
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_697
timestamp 1636968456
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_709
timestamp 1636968456
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_721
timestamp 1
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_727
timestamp 1
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_729
timestamp 1636968456
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_741
timestamp 1636968456
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_753
timestamp 1636968456
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_765
timestamp 1636968456
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_777
timestamp 1
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_783
timestamp 1
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_785
timestamp 1636968456
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_797
timestamp 1636968456
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_809
timestamp 1636968456
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_821
timestamp 1636968456
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_833
timestamp 1
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_839
timestamp 1
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_841
timestamp 1
transform 1 0 78476 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1636968456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1636968456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1636968456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1636968456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1636968456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1636968456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1636968456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_309
timestamp 1
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_317
timestamp 1636968456
transform 1 0 30268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_329
timestamp 1
transform 1 0 31372 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_335
timestamp 1
transform 1 0 31924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_356
timestamp 1
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_365
timestamp 1
transform 1 0 34684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_409
timestamp 1
transform 1 0 38732 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_417
timestamp 1
transform 1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_449
timestamp 1
transform 1 0 42412 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_473
timestamp 1
transform 1 0 44620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_484
timestamp 1
transform 1 0 45632 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_492
timestamp 1
transform 1 0 46368 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_509
timestamp 1636968456
transform 1 0 47932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_521
timestamp 1
transform 1 0 49036 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_529
timestamp 1
transform 1 0 49772 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_553
timestamp 1636968456
transform 1 0 51980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_565
timestamp 1
transform 1 0 53084 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_575
timestamp 1636968456
transform 1 0 54004 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 1
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 1636968456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 1636968456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 1636968456
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_625
timestamp 1636968456
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_637
timestamp 1
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_643
timestamp 1
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_645
timestamp 1636968456
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_657
timestamp 1636968456
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_669
timestamp 1636968456
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_681
timestamp 1636968456
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_693
timestamp 1
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_699
timestamp 1
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_701
timestamp 1636968456
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_713
timestamp 1636968456
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_725
timestamp 1636968456
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_737
timestamp 1636968456
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_749
timestamp 1
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_755
timestamp 1
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_757
timestamp 1636968456
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_769
timestamp 1636968456
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_781
timestamp 1636968456
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_793
timestamp 1636968456
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_805
timestamp 1
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_811
timestamp 1
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_813
timestamp 1636968456
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_825
timestamp 1636968456
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636968456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636968456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1636968456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1636968456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1636968456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1636968456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1636968456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1636968456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1636968456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1636968456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1636968456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1636968456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1636968456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1636968456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_317
timestamp 1
transform 1 0 30268 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_323
timestamp 1
transform 1 0 30820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_331
timestamp 1
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_337
timestamp 1
transform 1 0 32108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_345
timestamp 1
transform 1 0 32844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_352
timestamp 1
transform 1 0 33488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_362
timestamp 1
transform 1 0 34408 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_372
timestamp 1
transform 1 0 35328 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_399
timestamp 1
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_403
timestamp 1
transform 1 0 38180 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_412
timestamp 1636968456
transform 1 0 39008 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_424
timestamp 1636968456
transform 1 0 40112 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_436
timestamp 1636968456
transform 1 0 41216 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_449
timestamp 1
transform 1 0 42412 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_469
timestamp 1636968456
transform 1 0 44252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_481
timestamp 1636968456
transform 1 0 45356 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_493
timestamp 1
transform 1 0 46460 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_501
timestamp 1
transform 1 0 47196 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_505
timestamp 1636968456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_517
timestamp 1
transform 1 0 48668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_525
timestamp 1
transform 1 0 49404 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_540
timestamp 1
transform 1 0 50784 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_548
timestamp 1
transform 1 0 51520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_557
timestamp 1
transform 1 0 52348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_561
timestamp 1
transform 1 0 52716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_578
timestamp 1
transform 1 0 54280 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_588
timestamp 1636968456
transform 1 0 55200 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_600
timestamp 1636968456
transform 1 0 56304 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_612
timestamp 1
transform 1 0 57408 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_617
timestamp 1636968456
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_629
timestamp 1636968456
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_641
timestamp 1636968456
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_653
timestamp 1636968456
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_665
timestamp 1
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_671
timestamp 1
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_673
timestamp 1636968456
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_685
timestamp 1636968456
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_697
timestamp 1636968456
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_709
timestamp 1636968456
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_721
timestamp 1
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_727
timestamp 1
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_729
timestamp 1636968456
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_741
timestamp 1636968456
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_753
timestamp 1636968456
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_765
timestamp 1636968456
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_777
timestamp 1
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_783
timestamp 1
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_785
timestamp 1636968456
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_797
timestamp 1636968456
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_809
timestamp 1636968456
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_821
timestamp 1636968456
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_833
timestamp 1
transform 1 0 77740 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_841
timestamp 1
transform 1 0 78476 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1636968456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1636968456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1636968456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1636968456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1636968456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1636968456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1636968456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1636968456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1636968456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1636968456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1636968456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_309
timestamp 1
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_317
timestamp 1
transform 1 0 30268 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_340
timestamp 1636968456
transform 1 0 32384 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_360
timestamp 1
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_373
timestamp 1636968456
transform 1 0 35420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_385
timestamp 1
transform 1 0 36524 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_394
timestamp 1
transform 1 0 37352 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_398
timestamp 1
transform 1 0 37720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1636968456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_433
timestamp 1
transform 1 0 40940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_437
timestamp 1
transform 1 0 41308 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_446
timestamp 1636968456
transform 1 0 42136 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_458
timestamp 1636968456
transform 1 0 43240 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_470
timestamp 1
transform 1 0 44344 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_497
timestamp 1636968456
transform 1 0 46828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_509
timestamp 1636968456
transform 1 0 47932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_521
timestamp 1
transform 1 0 49036 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_599
timestamp 1636968456
transform 1 0 56212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_611
timestamp 1636968456
transform 1 0 57316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_623
timestamp 1636968456
transform 1 0 58420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_635
timestamp 1
transform 1 0 59524 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_643
timestamp 1
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_645
timestamp 1636968456
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_657
timestamp 1636968456
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_669
timestamp 1636968456
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_681
timestamp 1636968456
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_693
timestamp 1
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_699
timestamp 1
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_701
timestamp 1636968456
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_713
timestamp 1636968456
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_725
timestamp 1636968456
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_737
timestamp 1636968456
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_749
timestamp 1
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_755
timestamp 1
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_757
timestamp 1636968456
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_769
timestamp 1636968456
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_781
timestamp 1636968456
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_793
timestamp 1636968456
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_805
timestamp 1
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_811
timestamp 1
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_813
timestamp 1636968456
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_825
timestamp 1
transform 1 0 77004 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_831
timestamp 1
transform 1 0 77556 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_837
timestamp 1
transform 1 0 78108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1636968456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1636968456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1636968456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1636968456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1636968456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1636968456
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1636968456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1636968456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1636968456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1636968456
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1636968456
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1636968456
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1636968456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1636968456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1636968456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1636968456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1636968456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1636968456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_305
timestamp 1
transform 1 0 29164 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_313
timestamp 1
transform 1 0 29900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_337
timestamp 1
transform 1 0 32108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_345
timestamp 1
transform 1 0 32844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_355
timestamp 1
transform 1 0 33764 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_363
timestamp 1
transform 1 0 34500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_386
timestamp 1
transform 1 0 36616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_393
timestamp 1
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_401
timestamp 1
transform 1 0 37996 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_410
timestamp 1
transform 1 0 38824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_422
timestamp 1
transform 1 0 39928 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_444
timestamp 1
transform 1 0 41952 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_449
timestamp 1
transform 1 0 42412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_462
timestamp 1
transform 1 0 43608 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_468
timestamp 1
transform 1 0 44160 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_496
timestamp 1
transform 1 0 46736 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_545
timestamp 1636968456
transform 1 0 51244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_557
timestamp 1
transform 1 0 52348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_561
timestamp 1
transform 1 0 52716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_579
timestamp 1
transform 1 0 54372 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_589
timestamp 1636968456
transform 1 0 55292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_601
timestamp 1636968456
transform 1 0 56396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_613
timestamp 1
transform 1 0 57500 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_617
timestamp 1636968456
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_629
timestamp 1636968456
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_641
timestamp 1636968456
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_653
timestamp 1636968456
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_665
timestamp 1
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_671
timestamp 1
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_673
timestamp 1636968456
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_685
timestamp 1636968456
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_697
timestamp 1636968456
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_709
timestamp 1636968456
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_721
timestamp 1
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_727
timestamp 1
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_729
timestamp 1636968456
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_741
timestamp 1636968456
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_753
timestamp 1636968456
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_765
timestamp 1636968456
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_777
timestamp 1
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_783
timestamp 1
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_785
timestamp 1636968456
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_797
timestamp 1636968456
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_809
timestamp 1636968456
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_821
timestamp 1636968456
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_833
timestamp 1
transform 1 0 77740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_841
timestamp 1
transform 1 0 78476 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1636968456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1636968456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1636968456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1636968456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1636968456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1636968456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1636968456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1636968456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1636968456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1636968456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1636968456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1636968456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1636968456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1636968456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1636968456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1636968456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1636968456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1636968456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_309
timestamp 1
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_362
timestamp 1
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_365
timestamp 1
transform 1 0 34684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_375
timestamp 1
transform 1 0 35604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_379
timestamp 1
transform 1 0 35972 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_399
timestamp 1
transform 1 0 37812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_410
timestamp 1
transform 1 0 38824 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_418
timestamp 1
transform 1 0 39560 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_421
timestamp 1
transform 1 0 39836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_427
timestamp 1
transform 1 0 40388 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_452
timestamp 1
transform 1 0 42688 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_479
timestamp 1
transform 1 0 45172 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_487
timestamp 1
transform 1 0 45908 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_506
timestamp 1636968456
transform 1 0 47656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_518
timestamp 1
transform 1 0 48760 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_531
timestamp 1
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_533
timestamp 1636968456
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_545
timestamp 1636968456
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_557
timestamp 1
transform 1 0 52348 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_565
timestamp 1
transform 1 0 53084 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_569
timestamp 1636968456
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_581
timestamp 1
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_587
timestamp 1
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_589
timestamp 1636968456
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_601
timestamp 1636968456
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_613
timestamp 1636968456
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_625
timestamp 1636968456
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_637
timestamp 1
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_643
timestamp 1
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_645
timestamp 1636968456
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_657
timestamp 1636968456
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_669
timestamp 1636968456
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_681
timestamp 1636968456
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_693
timestamp 1
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_699
timestamp 1
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_701
timestamp 1636968456
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_713
timestamp 1636968456
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_725
timestamp 1636968456
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_737
timestamp 1636968456
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_749
timestamp 1
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_755
timestamp 1
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_757
timestamp 1636968456
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_769
timestamp 1636968456
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_781
timestamp 1636968456
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_793
timestamp 1636968456
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_805
timestamp 1
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_811
timestamp 1
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_813
timestamp 1636968456
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_825
timestamp 1
transform 1 0 77004 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_831
timestamp 1
transform 1 0 77556 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_837
timestamp 1
transform 1 0 78108 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_841
timestamp 1
transform 1 0 78476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1636968456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1636968456
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1636968456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1636968456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1636968456
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1636968456
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1636968456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1636968456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1636968456
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1636968456
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1636968456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1636968456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1636968456
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1636968456
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1636968456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1636968456
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1636968456
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1636968456
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1636968456
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1636968456
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1636968456
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_317
timestamp 1
transform 1 0 30268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_321
timestamp 1
transform 1 0 30636 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_329
timestamp 1
transform 1 0 31372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_334
timestamp 1
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_359
timestamp 1636968456
transform 1 0 34132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_371
timestamp 1636968456
transform 1 0 35236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_383
timestamp 1
transform 1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_413
timestamp 1636968456
transform 1 0 39100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_425
timestamp 1636968456
transform 1 0 40204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_437
timestamp 1
transform 1 0 41308 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_445
timestamp 1
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_456
timestamp 1
transform 1 0 43056 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_469
timestamp 1636968456
transform 1 0 44252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_481
timestamp 1636968456
transform 1 0 45356 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_493
timestamp 1
transform 1 0 46460 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_501
timestamp 1
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_505
timestamp 1636968456
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_517
timestamp 1
transform 1 0 48668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_525
timestamp 1
transform 1 0 49404 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_535
timestamp 1636968456
transform 1 0 50324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_547
timestamp 1
transform 1 0 51428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_554
timestamp 1
transform 1 0 52072 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_577
timestamp 1
transform 1 0 54188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_608
timestamp 1
transform 1 0 57040 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_617
timestamp 1636968456
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_629
timestamp 1636968456
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_641
timestamp 1636968456
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_653
timestamp 1636968456
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_665
timestamp 1
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_671
timestamp 1
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_673
timestamp 1636968456
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_685
timestamp 1636968456
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_697
timestamp 1636968456
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_709
timestamp 1636968456
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_721
timestamp 1
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_727
timestamp 1
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_729
timestamp 1636968456
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_741
timestamp 1636968456
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_753
timestamp 1636968456
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_765
timestamp 1636968456
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_777
timestamp 1
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_783
timestamp 1
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_785
timestamp 1636968456
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_797
timestamp 1636968456
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_809
timestamp 1636968456
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_821
timestamp 1
transform 1 0 76636 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_829
timestamp 1
transform 1 0 77372 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_841
timestamp 1
transform 1 0 78476 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636968456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1636968456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1636968456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1636968456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1636968456
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1636968456
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1636968456
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1636968456
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1636968456
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1636968456
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1636968456
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1636968456
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1636968456
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1636968456
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1636968456
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1636968456
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1636968456
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1636968456
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1636968456
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1636968456
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1636968456
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_309
timestamp 1
transform 1 0 29532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_315
timestamp 1
transform 1 0 30084 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_337
timestamp 1636968456
transform 1 0 32108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_349
timestamp 1636968456
transform 1 0 33212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_361
timestamp 1
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_365
timestamp 1
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_376
timestamp 1
transform 1 0 35696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_383
timestamp 1
transform 1 0 36340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_387
timestamp 1
transform 1 0 36708 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_395
timestamp 1
transform 1 0 37444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_417
timestamp 1
transform 1 0 39468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_441
timestamp 1
transform 1 0 41676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_456
timestamp 1
transform 1 0 43056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_461
timestamp 1
transform 1 0 43516 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_469
timestamp 1
transform 1 0 44252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_473
timestamp 1
transform 1 0 44620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_479
timestamp 1
transform 1 0 45172 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_508
timestamp 1
transform 1 0 47840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_537
timestamp 1
transform 1 0 50508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_543
timestamp 1
transform 1 0 51060 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_564
timestamp 1
transform 1 0 52992 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 1
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_596
timestamp 1636968456
transform 1 0 55936 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_608
timestamp 1636968456
transform 1 0 57040 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_620
timestamp 1636968456
transform 1 0 58144 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_632
timestamp 1636968456
transform 1 0 59248 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_645
timestamp 1636968456
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_657
timestamp 1636968456
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_669
timestamp 1636968456
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_681
timestamp 1636968456
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_693
timestamp 1
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_699
timestamp 1
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_701
timestamp 1636968456
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_713
timestamp 1636968456
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_725
timestamp 1636968456
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_737
timestamp 1636968456
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_749
timestamp 1
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_755
timestamp 1
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_757
timestamp 1636968456
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_769
timestamp 1636968456
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_781
timestamp 1636968456
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_793
timestamp 1636968456
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_805
timestamp 1
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_811
timestamp 1
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_813
timestamp 1636968456
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_825
timestamp 1
transform 1 0 77004 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_837
timestamp 1
transform 1 0 78108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1636968456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1636968456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1636968456
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1636968456
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1636968456
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1636968456
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1636968456
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1636968456
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1636968456
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1636968456
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1636968456
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1636968456
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1636968456
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1636968456
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1636968456
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1636968456
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1636968456
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1636968456
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_293
timestamp 1
transform 1 0 28060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_301
timestamp 1
transform 1 0 28796 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_322
timestamp 1
transform 1 0 30728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_333
timestamp 1
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_337
timestamp 1
transform 1 0 32108 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_351
timestamp 1636968456
transform 1 0 33396 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_363
timestamp 1
transform 1 0 34500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_385
timestamp 1
transform 1 0 36524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_399
timestamp 1
transform 1 0 37812 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_410
timestamp 1636968456
transform 1 0 38824 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_422
timestamp 1
transform 1 0 39928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_426
timestamp 1
transform 1 0 40296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_459
timestamp 1
transform 1 0 43332 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_483
timestamp 1
transform 1 0 45540 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_505
timestamp 1
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_513
timestamp 1
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_523
timestamp 1
transform 1 0 49220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_555
timestamp 1
transform 1 0 52164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_559
timestamp 1
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_561
timestamp 1
transform 1 0 52716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_566
timestamp 1
transform 1 0 53176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_573
timestamp 1
transform 1 0 53820 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_587
timestamp 1636968456
transform 1 0 55108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_599
timestamp 1636968456
transform 1 0 56212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_611
timestamp 1
transform 1 0 57316 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 1
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_617
timestamp 1636968456
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_629
timestamp 1636968456
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_641
timestamp 1636968456
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_653
timestamp 1636968456
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_665
timestamp 1
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_671
timestamp 1
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_673
timestamp 1636968456
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_685
timestamp 1636968456
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_697
timestamp 1636968456
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_709
timestamp 1636968456
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_721
timestamp 1
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_727
timestamp 1
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_729
timestamp 1636968456
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_741
timestamp 1636968456
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_753
timestamp 1636968456
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_765
timestamp 1636968456
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_777
timestamp 1
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_783
timestamp 1
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_785
timestamp 1636968456
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_797
timestamp 1636968456
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_809
timestamp 1636968456
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_821
timestamp 1636968456
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_833
timestamp 1
transform 1 0 77740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_841
timestamp 1
transform 1 0 78476 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1636968456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1636968456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1636968456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1636968456
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1636968456
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1636968456
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1636968456
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1636968456
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1636968456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1636968456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1636968456
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1636968456
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1636968456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1636968456
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1636968456
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1636968456
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1636968456
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_265
timestamp 1
transform 1 0 25484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_273
timestamp 1
transform 1 0 26220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_298
timestamp 1
transform 1 0 28520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_306
timestamp 1
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1636968456
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_327
timestamp 1
transform 1 0 31188 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_335
timestamp 1
transform 1 0 31924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_373
timestamp 1
transform 1 0 35420 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_377
timestamp 1
transform 1 0 35788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_398
timestamp 1
transform 1 0 37720 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_402
timestamp 1
transform 1 0 38088 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_410
timestamp 1
transform 1 0 38824 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_418
timestamp 1
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1636968456
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_433
timestamp 1
transform 1 0 40940 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_449
timestamp 1
transform 1 0 42412 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_453
timestamp 1
transform 1 0 42780 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_456
timestamp 1
transform 1 0 43056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_472
timestamp 1
transform 1 0 44528 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_477
timestamp 1
transform 1 0 44988 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_483
timestamp 1636968456
transform 1 0 45540 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_495
timestamp 1636968456
transform 1 0 46644 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_507
timestamp 1636968456
transform 1 0 47748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_519
timestamp 1
transform 1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_524
timestamp 1
transform 1 0 49312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 1
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_535
timestamp 1
transform 1 0 50324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_551
timestamp 1636968456
transform 1 0 51796 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_563
timestamp 1636968456
transform 1 0 52900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_575
timestamp 1636968456
transform 1 0 54004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 1
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_589
timestamp 1636968456
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_601
timestamp 1636968456
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_613
timestamp 1636968456
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_625
timestamp 1636968456
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_637
timestamp 1
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_643
timestamp 1
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_645
timestamp 1636968456
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_657
timestamp 1636968456
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_669
timestamp 1636968456
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_681
timestamp 1636968456
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_693
timestamp 1
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_699
timestamp 1
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_701
timestamp 1636968456
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_713
timestamp 1636968456
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_725
timestamp 1636968456
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_737
timestamp 1636968456
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_749
timestamp 1
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_755
timestamp 1
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_757
timestamp 1636968456
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_769
timestamp 1636968456
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_781
timestamp 1636968456
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_793
timestamp 1636968456
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_805
timestamp 1
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_811
timestamp 1
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_813
timestamp 1636968456
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_825
timestamp 1636968456
transform 1 0 77004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_837
timestamp 1
transform 1 0 78108 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_841
timestamp 1
transform 1 0 78476 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1636968456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1636968456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1636968456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1636968456
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1636968456
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1636968456
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1636968456
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1636968456
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1636968456
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1636968456
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1636968456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1636968456
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1636968456
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1636968456
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1636968456
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1636968456
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1636968456
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1636968456
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_281
timestamp 1
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_315
timestamp 1636968456
transform 1 0 30084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_327
timestamp 1
transform 1 0 31188 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_337
timestamp 1
transform 1 0 32108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_351
timestamp 1
transform 1 0 33396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_362
timestamp 1
transform 1 0 34408 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_379
timestamp 1636968456
transform 1 0 35972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_393
timestamp 1
transform 1 0 37260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_438
timestamp 1
transform 1 0 41400 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_466
timestamp 1636968456
transform 1 0 43976 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_478
timestamp 1
transform 1 0 45080 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_491
timestamp 1636968456
transform 1 0 46276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 1
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_505
timestamp 1636968456
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_532
timestamp 1
transform 1 0 50048 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_553
timestamp 1
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_559
timestamp 1
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_561
timestamp 1
transform 1 0 52716 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_568
timestamp 1636968456
transform 1 0 53360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_594
timestamp 1
transform 1 0 55752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_605
timestamp 1
transform 1 0 56764 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_613
timestamp 1
transform 1 0 57500 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_617
timestamp 1636968456
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_629
timestamp 1636968456
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_641
timestamp 1636968456
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_653
timestamp 1636968456
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_665
timestamp 1
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_671
timestamp 1
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_673
timestamp 1636968456
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_685
timestamp 1636968456
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_697
timestamp 1636968456
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_709
timestamp 1636968456
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_721
timestamp 1
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_727
timestamp 1
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_729
timestamp 1636968456
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_741
timestamp 1636968456
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_753
timestamp 1636968456
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_765
timestamp 1636968456
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_777
timestamp 1
transform 1 0 72588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_783
timestamp 1
transform 1 0 73140 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_785
timestamp 1636968456
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_797
timestamp 1636968456
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_809
timestamp 1636968456
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_821
timestamp 1636968456
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_833
timestamp 1
transform 1 0 77740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_839
timestamp 1
transform 1 0 78292 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_841
timestamp 1
transform 1 0 78476 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1636968456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1636968456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1636968456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1636968456
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1636968456
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1636968456
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1636968456
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1636968456
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1636968456
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1636968456
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1636968456
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1636968456
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_201
timestamp 1
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_204
timestamp 1636968456
transform 1 0 19872 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_216
timestamp 1636968456
transform 1 0 20976 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_228
timestamp 1636968456
transform 1 0 22080 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_240
timestamp 1636968456
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_253
timestamp 1
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_261
timestamp 1
transform 1 0 25116 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_284
timestamp 1636968456
transform 1 0 27232 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_296
timestamp 1636968456
transform 1 0 28336 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1636968456
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_321
timestamp 1
transform 1 0 30636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_354
timestamp 1
transform 1 0 33672 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_373
timestamp 1636968456
transform 1 0 35420 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_385
timestamp 1636968456
transform 1 0 36524 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_397
timestamp 1
transform 1 0 37628 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_405
timestamp 1
transform 1 0 38364 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_421
timestamp 1
transform 1 0 39836 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_462
timestamp 1
transform 1 0 43608 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_469
timestamp 1
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_475
timestamp 1
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_477
timestamp 1
transform 1 0 44988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_508
timestamp 1
transform 1 0 47840 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_551
timestamp 1
transform 1 0 51796 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_611
timestamp 1636968456
transform 1 0 57316 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_623
timestamp 1636968456
transform 1 0 58420 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_635
timestamp 1
transform 1 0 59524 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_643
timestamp 1
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_645
timestamp 1636968456
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_657
timestamp 1636968456
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_669
timestamp 1636968456
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_681
timestamp 1636968456
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_693
timestamp 1
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_699
timestamp 1
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_701
timestamp 1636968456
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_713
timestamp 1636968456
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_725
timestamp 1636968456
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_737
timestamp 1636968456
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_749
timestamp 1
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_755
timestamp 1
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_757
timestamp 1636968456
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_769
timestamp 1636968456
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_781
timestamp 1636968456
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_793
timestamp 1636968456
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_805
timestamp 1
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_811
timestamp 1
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_813
timestamp 1636968456
transform 1 0 75900 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_825
timestamp 1636968456
transform 1 0 77004 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_837
timestamp 1
transform 1 0 78108 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_841
timestamp 1
transform 1 0 78476 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1636968456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1636968456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1636968456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1636968456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1636968456
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1636968456
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1636968456
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1636968456
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1636968456
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1636968456
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1636968456
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1636968456
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_181
timestamp 1
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1636968456
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1636968456
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1636968456
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_261
timestamp 1
transform 1 0 25116 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_269
timestamp 1
transform 1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1636968456
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_293
timestamp 1
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_304
timestamp 1
transform 1 0 29072 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_312
timestamp 1636968456
transform 1 0 29808 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_324
timestamp 1636968456
transform 1 0 30912 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_345
timestamp 1
transform 1 0 32844 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_374
timestamp 1
transform 1 0 35512 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_388
timestamp 1
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_393
timestamp 1
transform 1 0 37260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_412
timestamp 1
transform 1 0 39008 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_418
timestamp 1636968456
transform 1 0 39560 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_430
timestamp 1
transform 1 0 40664 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_497
timestamp 1
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_503
timestamp 1
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_537
timestamp 1
transform 1 0 50508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_554
timestamp 1
transform 1 0 52072 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_561
timestamp 1636968456
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_573
timestamp 1
transform 1 0 53820 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_586
timestamp 1636968456
transform 1 0 55016 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_598
timestamp 1636968456
transform 1 0 56120 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_610
timestamp 1
transform 1 0 57224 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_617
timestamp 1636968456
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_629
timestamp 1636968456
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_641
timestamp 1636968456
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_653
timestamp 1636968456
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_665
timestamp 1
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_671
timestamp 1
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_673
timestamp 1636968456
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_685
timestamp 1636968456
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_697
timestamp 1636968456
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_709
timestamp 1636968456
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_721
timestamp 1
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_727
timestamp 1
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_729
timestamp 1636968456
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_741
timestamp 1636968456
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_753
timestamp 1636968456
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_765
timestamp 1636968456
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_777
timestamp 1
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_783
timestamp 1
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_785
timestamp 1636968456
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_797
timestamp 1636968456
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_809
timestamp 1636968456
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_821
timestamp 1636968456
transform 1 0 76636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_833
timestamp 1
transform 1 0 77740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_839
timestamp 1
transform 1 0 78292 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_841
timestamp 1
transform 1 0 78476 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1636968456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1636968456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1636968456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1636968456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1636968456
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1636968456
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1636968456
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1636968456
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1636968456
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1636968456
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1636968456
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_165
timestamp 1
transform 1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_173
timestamp 1
transform 1 0 17020 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1636968456
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_209
timestamp 1
transform 1 0 20332 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_234
timestamp 1
transform 1 0 22632 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_238
timestamp 1
transform 1 0 23000 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_244
timestamp 1
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_253
timestamp 1
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_261
timestamp 1
transform 1 0 25116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_280
timestamp 1
transform 1 0 26864 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_288
timestamp 1
transform 1 0 27600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_300
timestamp 1
transform 1 0 28704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_309
timestamp 1
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_322
timestamp 1636968456
transform 1 0 30728 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_334
timestamp 1636968456
transform 1 0 31832 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_346
timestamp 1636968456
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_358
timestamp 1
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_365
timestamp 1
transform 1 0 34684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_373
timestamp 1
transform 1 0 35420 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_396
timestamp 1
transform 1 0 37536 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 1636968456
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_433
timestamp 1
transform 1 0 40940 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_441
timestamp 1
transform 1 0 41676 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_451
timestamp 1
transform 1 0 42596 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_463
timestamp 1
transform 1 0 43700 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_474
timestamp 1
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_477
timestamp 1
transform 1 0 44988 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_487
timestamp 1636968456
transform 1 0 45908 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_499
timestamp 1636968456
transform 1 0 47012 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_511
timestamp 1
transform 1 0 48116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_515
timestamp 1
transform 1 0 48484 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_522
timestamp 1
transform 1 0 49128 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_530
timestamp 1
transform 1 0 49864 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_533
timestamp 1636968456
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_545
timestamp 1
transform 1 0 51244 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_551
timestamp 1
transform 1 0 51796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_567
timestamp 1
transform 1 0 53268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_579
timestamp 1
transform 1 0 54372 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_587
timestamp 1
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_589
timestamp 1636968456
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_601
timestamp 1636968456
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_613
timestamp 1636968456
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_625
timestamp 1636968456
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_637
timestamp 1
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_643
timestamp 1
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_645
timestamp 1636968456
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_657
timestamp 1636968456
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_669
timestamp 1636968456
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_681
timestamp 1636968456
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_693
timestamp 1
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_699
timestamp 1
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_701
timestamp 1636968456
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_713
timestamp 1636968456
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_725
timestamp 1636968456
transform 1 0 67804 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_737
timestamp 1636968456
transform 1 0 68908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_749
timestamp 1
transform 1 0 70012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_755
timestamp 1
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_757
timestamp 1636968456
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_769
timestamp 1636968456
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_781
timestamp 1636968456
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_793
timestamp 1636968456
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_805
timestamp 1
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_811
timestamp 1
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_813
timestamp 1636968456
transform 1 0 75900 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_825
timestamp 1636968456
transform 1 0 77004 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_837
timestamp 1
transform 1 0 78108 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_841
timestamp 1
transform 1 0 78476 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1636968456
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1636968456
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1636968456
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1636968456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1636968456
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1636968456
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1636968456
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1636968456
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_125
timestamp 1
transform 1 0 12604 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_146
timestamp 1636968456
transform 1 0 14536 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_158
timestamp 1
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_169
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_183
timestamp 1636968456
transform 1 0 17940 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_195
timestamp 1636968456
transform 1 0 19044 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_207
timestamp 1636968456
transform 1 0 20148 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_219
timestamp 1
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_225
timestamp 1
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_233
timestamp 1
transform 1 0 22540 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_255
timestamp 1
transform 1 0 24564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_261
timestamp 1
transform 1 0 25116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_276
timestamp 1
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_281
timestamp 1
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_301
timestamp 1
transform 1 0 28796 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_307
timestamp 1
transform 1 0 29348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_328
timestamp 1
transform 1 0 31280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_337
timestamp 1
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_363
timestamp 1636968456
transform 1 0 34500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_375
timestamp 1
transform 1 0 35604 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_381
timestamp 1
transform 1 0 36156 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_401
timestamp 1
transform 1 0 37996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_409
timestamp 1
transform 1 0 38732 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_428
timestamp 1636968456
transform 1 0 40480 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_440
timestamp 1
transform 1 0 41584 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_449
timestamp 1636968456
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_461
timestamp 1636968456
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_473
timestamp 1636968456
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_485
timestamp 1636968456
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_497
timestamp 1
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_503
timestamp 1
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_505
timestamp 1
transform 1 0 47564 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_535
timestamp 1
transform 1 0 50324 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_546
timestamp 1
transform 1 0 51336 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_571
timestamp 1
transform 1 0 53636 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_597
timestamp 1636968456
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_609
timestamp 1
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_615
timestamp 1
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_617
timestamp 1636968456
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_629
timestamp 1636968456
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_641
timestamp 1636968456
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_653
timestamp 1636968456
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_665
timestamp 1
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_671
timestamp 1
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_673
timestamp 1636968456
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_685
timestamp 1636968456
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_697
timestamp 1636968456
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_709
timestamp 1636968456
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_721
timestamp 1
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_727
timestamp 1
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_729
timestamp 1636968456
transform 1 0 68172 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_741
timestamp 1636968456
transform 1 0 69276 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_753
timestamp 1636968456
transform 1 0 70380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_765
timestamp 1636968456
transform 1 0 71484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_777
timestamp 1
transform 1 0 72588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_783
timestamp 1
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_785
timestamp 1636968456
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_797
timestamp 1636968456
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_809
timestamp 1636968456
transform 1 0 75532 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_821
timestamp 1636968456
transform 1 0 76636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_833
timestamp 1
transform 1 0 77740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_839
timestamp 1
transform 1 0 78292 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_841
timestamp 1
transform 1 0 78476 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636968456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1636968456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1636968456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1636968456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1636968456
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1636968456
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1636968456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1636968456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1636968456
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1636968456
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_147
timestamp 1
transform 1 0 14628 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_190
timestamp 1
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_205
timestamp 1
transform 1 0 19964 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_213
timestamp 1
transform 1 0 20700 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_219
timestamp 1636968456
transform 1 0 21252 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_231
timestamp 1
transform 1 0 22356 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_239
timestamp 1
transform 1 0 23092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_256
timestamp 1
transform 1 0 24656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_268
timestamp 1
transform 1 0 25760 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_276
timestamp 1
transform 1 0 26496 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_306
timestamp 1
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1636968456
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_321
timestamp 1
transform 1 0 30636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_325
timestamp 1
transform 1 0 31004 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_346
timestamp 1
transform 1 0 32936 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_361
timestamp 1
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_365
timestamp 1
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_376
timestamp 1636968456
transform 1 0 35696 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_388
timestamp 1
transform 1 0 36800 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_392
timestamp 1
transform 1 0 37168 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_397
timestamp 1
transform 1 0 37628 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_406
timestamp 1636968456
transform 1 0 38456 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_418
timestamp 1
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_421
timestamp 1
transform 1 0 39836 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_455
timestamp 1636968456
transform 1 0 42964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_467
timestamp 1
transform 1 0 44068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_472
timestamp 1
transform 1 0 44528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_477
timestamp 1
transform 1 0 44988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_486
timestamp 1
transform 1 0 45816 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_521
timestamp 1
transform 1 0 49036 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_529
timestamp 1
transform 1 0 49772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_533
timestamp 1
transform 1 0 50140 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_555
timestamp 1
transform 1 0 52164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_578
timestamp 1
transform 1 0 54280 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_586
timestamp 1
transform 1 0 55016 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_603
timestamp 1636968456
transform 1 0 56580 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_615
timestamp 1636968456
transform 1 0 57684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_627
timestamp 1636968456
transform 1 0 58788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_639
timestamp 1
transform 1 0 59892 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_643
timestamp 1
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_645
timestamp 1636968456
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_657
timestamp 1636968456
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_669
timestamp 1636968456
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_681
timestamp 1636968456
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_693
timestamp 1
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_699
timestamp 1
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_701
timestamp 1636968456
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_713
timestamp 1636968456
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_725
timestamp 1636968456
transform 1 0 67804 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_737
timestamp 1636968456
transform 1 0 68908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_749
timestamp 1
transform 1 0 70012 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_755
timestamp 1
transform 1 0 70564 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_757
timestamp 1636968456
transform 1 0 70748 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_769
timestamp 1636968456
transform 1 0 71852 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_781
timestamp 1636968456
transform 1 0 72956 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_793
timestamp 1636968456
transform 1 0 74060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_805
timestamp 1
transform 1 0 75164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_811
timestamp 1
transform 1 0 75716 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_813
timestamp 1636968456
transform 1 0 75900 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_825
timestamp 1636968456
transform 1 0 77004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_837
timestamp 1
transform 1 0 78108 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_841
timestamp 1
transform 1 0 78476 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1636968456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1636968456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1636968456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1636968456
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1636968456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1636968456
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1636968456
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1636968456
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1636968456
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_125
timestamp 1
transform 1 0 12604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_133
timestamp 1
transform 1 0 13340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_158
timestamp 1
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_169
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_209
timestamp 1
transform 1 0 20332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_213
timestamp 1
transform 1 0 20700 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_233
timestamp 1636968456
transform 1 0 22540 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_245
timestamp 1636968456
transform 1 0 23644 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_257
timestamp 1
transform 1 0 24748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_261
timestamp 1
transform 1 0 25116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_269
timestamp 1
transform 1 0 25852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_277
timestamp 1
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1636968456
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1636968456
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1636968456
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_317
timestamp 1
transform 1 0 30268 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_337
timestamp 1
transform 1 0 32108 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_360
timestamp 1
transform 1 0 34224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_384
timestamp 1
transform 1 0 36432 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_404
timestamp 1
transform 1 0 38272 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_412
timestamp 1636968456
transform 1 0 39008 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_424
timestamp 1
transform 1 0 40112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_433
timestamp 1
transform 1 0 40940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_445
timestamp 1
transform 1 0 42044 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_449
timestamp 1
transform 1 0 42412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_498
timestamp 1
transform 1 0 46920 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_505
timestamp 1636968456
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_517
timestamp 1636968456
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_529
timestamp 1
transform 1 0 49772 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_537
timestamp 1
transform 1 0 50508 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_545
timestamp 1636968456
transform 1 0 51244 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_557
timestamp 1
transform 1 0 52348 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_561
timestamp 1636968456
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_573
timestamp 1636968456
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_585
timestamp 1636968456
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_597
timestamp 1636968456
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_609
timestamp 1
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_615
timestamp 1
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_617
timestamp 1636968456
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_629
timestamp 1636968456
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_641
timestamp 1636968456
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_653
timestamp 1636968456
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_665
timestamp 1
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_671
timestamp 1
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_673
timestamp 1636968456
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_685
timestamp 1636968456
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_697
timestamp 1636968456
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_709
timestamp 1636968456
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_721
timestamp 1
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_727
timestamp 1
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_729
timestamp 1636968456
transform 1 0 68172 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_741
timestamp 1636968456
transform 1 0 69276 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_753
timestamp 1636968456
transform 1 0 70380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_765
timestamp 1636968456
transform 1 0 71484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_777
timestamp 1
transform 1 0 72588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_783
timestamp 1
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_785
timestamp 1636968456
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_797
timestamp 1636968456
transform 1 0 74428 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_809
timestamp 1636968456
transform 1 0 75532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_821
timestamp 1636968456
transform 1 0 76636 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_833
timestamp 1
transform 1 0 77740 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_839
timestamp 1
transform 1 0 78292 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_841
timestamp 1
transform 1 0 78476 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1636968456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1636968456
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1636968456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1636968456
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1636968456
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_77
timestamp 1
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_107
timestamp 1636968456
transform 1 0 10948 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_119
timestamp 1636968456
transform 1 0 12052 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_131
timestamp 1
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1636968456
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1636968456
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_165
timestamp 1
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp 1
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_205
timestamp 1636968456
transform 1 0 19964 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_217
timestamp 1
transform 1 0 21068 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_225
timestamp 1636968456
transform 1 0 21804 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_237
timestamp 1
transform 1 0 22908 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 1
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1636968456
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_265
timestamp 1
transform 1 0 25484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_273
timestamp 1
transform 1 0 26220 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_282
timestamp 1
transform 1 0 27048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_288
timestamp 1
transform 1 0 27600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_309
timestamp 1
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_320
timestamp 1636968456
transform 1 0 30544 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_332
timestamp 1
transform 1 0 31648 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_336
timestamp 1
transform 1 0 32016 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1636968456
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 1
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_365
timestamp 1
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_373
timestamp 1
transform 1 0 35420 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_385
timestamp 1
transform 1 0 36524 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_398
timestamp 1
transform 1 0 37720 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_410
timestamp 1
transform 1 0 38824 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_432
timestamp 1
transform 1 0 40848 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_440
timestamp 1636968456
transform 1 0 41584 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_452
timestamp 1
transform 1 0 42688 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_475
timestamp 1
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_485
timestamp 1636968456
transform 1 0 45724 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_497
timestamp 1636968456
transform 1 0 46828 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_509
timestamp 1636968456
transform 1 0 47932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_521
timestamp 1
transform 1 0 49036 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_529
timestamp 1
transform 1 0 49772 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_540
timestamp 1636968456
transform 1 0 50784 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_552
timestamp 1636968456
transform 1 0 51888 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_564
timestamp 1
transform 1 0 52992 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_572
timestamp 1
transform 1 0 53728 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_579
timestamp 1
transform 1 0 54372 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_587
timestamp 1
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_589
timestamp 1636968456
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_601
timestamp 1636968456
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_613
timestamp 1636968456
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_625
timestamp 1636968456
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_637
timestamp 1
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_643
timestamp 1
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_645
timestamp 1636968456
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_657
timestamp 1636968456
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_669
timestamp 1636968456
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_681
timestamp 1636968456
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_693
timestamp 1
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_699
timestamp 1
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_701
timestamp 1636968456
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_713
timestamp 1636968456
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_725
timestamp 1636968456
transform 1 0 67804 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_737
timestamp 1636968456
transform 1 0 68908 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_749
timestamp 1
transform 1 0 70012 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_755
timestamp 1
transform 1 0 70564 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_757
timestamp 1636968456
transform 1 0 70748 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_769
timestamp 1636968456
transform 1 0 71852 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_781
timestamp 1636968456
transform 1 0 72956 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_793
timestamp 1636968456
transform 1 0 74060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_805
timestamp 1
transform 1 0 75164 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_811
timestamp 1
transform 1 0 75716 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_813
timestamp 1636968456
transform 1 0 75900 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_825
timestamp 1636968456
transform 1 0 77004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_837
timestamp 1
transform 1 0 78108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_841
timestamp 1
transform 1 0 78476 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_8
timestamp 1636968456
transform 1 0 1840 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_20
timestamp 1636968456
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_32
timestamp 1636968456
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_44
timestamp 1636968456
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1636968456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_69
timestamp 1
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_73
timestamp 1
transform 1 0 7820 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_95
timestamp 1636968456
transform 1 0 9844 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_133
timestamp 1636968456
transform 1 0 13340 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_145
timestamp 1636968456
transform 1 0 14444 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_157
timestamp 1
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1636968456
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_190
timestamp 1636968456
transform 1 0 18584 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_202
timestamp 1636968456
transform 1 0 19688 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_214
timestamp 1
transform 1 0 20792 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_225
timestamp 1
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_243
timestamp 1
transform 1 0 23460 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_275
timestamp 1
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_281
timestamp 1
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_297
timestamp 1636968456
transform 1 0 28428 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_329
timestamp 1
transform 1 0 31372 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_337
timestamp 1
transform 1 0 32108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_350
timestamp 1
transform 1 0 33304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_354
timestamp 1
transform 1 0 33672 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_363
timestamp 1636968456
transform 1 0 34500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_375
timestamp 1
transform 1 0 35604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_379
timestamp 1
transform 1 0 35972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1636968456
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_405
timestamp 1636968456
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_417
timestamp 1
transform 1 0 39468 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_434
timestamp 1636968456
transform 1 0 41032 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_446
timestamp 1
transform 1 0 42136 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_449
timestamp 1636968456
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_461
timestamp 1
transform 1 0 43516 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_484
timestamp 1
transform 1 0 45632 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_501
timestamp 1
transform 1 0 47196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_507
timestamp 1
transform 1 0 47748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_528
timestamp 1
transform 1 0 49680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_550
timestamp 1
transform 1 0 51704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_559
timestamp 1
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_561
timestamp 1
transform 1 0 52716 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_569
timestamp 1
transform 1 0 53452 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_591
timestamp 1636968456
transform 1 0 55476 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_603
timestamp 1636968456
transform 1 0 56580 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_615
timestamp 1
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_617
timestamp 1636968456
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_629
timestamp 1636968456
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_641
timestamp 1636968456
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_653
timestamp 1636968456
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_665
timestamp 1
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_671
timestamp 1
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_673
timestamp 1636968456
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_685
timestamp 1636968456
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_697
timestamp 1636968456
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_709
timestamp 1636968456
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_721
timestamp 1
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_727
timestamp 1
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_729
timestamp 1636968456
transform 1 0 68172 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_741
timestamp 1636968456
transform 1 0 69276 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_753
timestamp 1636968456
transform 1 0 70380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_765
timestamp 1636968456
transform 1 0 71484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_777
timestamp 1
transform 1 0 72588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_783
timestamp 1
transform 1 0 73140 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_785
timestamp 1636968456
transform 1 0 73324 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_797
timestamp 1636968456
transform 1 0 74428 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_809
timestamp 1636968456
transform 1 0 75532 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_821
timestamp 1636968456
transform 1 0 76636 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_833
timestamp 1
transform 1 0 77740 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_839
timestamp 1
transform 1 0 78292 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_841
timestamp 1
transform 1 0 78476 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_8
timestamp 1636968456
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_20
timestamp 1
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1636968456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1636968456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_65
timestamp 1
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_74
timestamp 1
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1636968456
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1636968456
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_109
timestamp 1
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_117
timestamp 1
transform 1 0 11868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_127
timestamp 1
transform 1 0 12788 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_136
timestamp 1
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_149
timestamp 1
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_186
timestamp 1
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_215
timestamp 1636968456
transform 1 0 20884 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_227
timestamp 1
transform 1 0 21988 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_239
timestamp 1
transform 1 0 23092 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1636968456
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1636968456
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_277
timestamp 1
transform 1 0 26588 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_295
timestamp 1636968456
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_309
timestamp 1
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_320
timestamp 1
transform 1 0 30544 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_360
timestamp 1
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_369
timestamp 1
transform 1 0 35052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_373
timestamp 1
transform 1 0 35420 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_401
timestamp 1636968456
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_413
timestamp 1
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 1
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 1636968456
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_433
timestamp 1
transform 1 0 40940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_437
timestamp 1
transform 1 0 41308 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_446
timestamp 1
transform 1 0 42136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_458
timestamp 1
transform 1 0 43240 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_475
timestamp 1
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_481
timestamp 1
transform 1 0 45356 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_520
timestamp 1
transform 1 0 48944 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_540
timestamp 1
transform 1 0 50784 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_587
timestamp 1
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_589
timestamp 1636968456
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_601
timestamp 1636968456
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_613
timestamp 1636968456
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_625
timestamp 1636968456
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_637
timestamp 1
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_643
timestamp 1
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_645
timestamp 1636968456
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_657
timestamp 1636968456
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_669
timestamp 1636968456
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_681
timestamp 1636968456
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_693
timestamp 1
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_699
timestamp 1
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_701
timestamp 1636968456
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_713
timestamp 1636968456
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_725
timestamp 1636968456
transform 1 0 67804 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_737
timestamp 1636968456
transform 1 0 68908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_749
timestamp 1
transform 1 0 70012 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_755
timestamp 1
transform 1 0 70564 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_757
timestamp 1636968456
transform 1 0 70748 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_769
timestamp 1636968456
transform 1 0 71852 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_781
timestamp 1636968456
transform 1 0 72956 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_793
timestamp 1636968456
transform 1 0 74060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_805
timestamp 1
transform 1 0 75164 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_811
timestamp 1
transform 1 0 75716 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_813
timestamp 1636968456
transform 1 0 75900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_825
timestamp 1636968456
transform 1 0 77004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_837
timestamp 1
transform 1 0 78108 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_841
timestamp 1
transform 1 0 78476 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1636968456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1636968456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1636968456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1636968456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_79
timestamp 1
transform 1 0 8372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_86
timestamp 1
transform 1 0 9016 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_90
timestamp 1
transform 1 0 9384 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1636968456
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_125
timestamp 1
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_134
timestamp 1636968456
transform 1 0 13432 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_146
timestamp 1636968456
transform 1 0 14536 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_158
timestamp 1
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_176
timestamp 1636968456
transform 1 0 17296 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_188
timestamp 1
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_212
timestamp 1636968456
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_225
timestamp 1
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_231
timestamp 1
transform 1 0 22356 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_235
timestamp 1
transform 1 0 22724 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_243
timestamp 1
transform 1 0 23460 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_247
timestamp 1
transform 1 0 23828 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_253
timestamp 1
transform 1 0 24380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_261
timestamp 1
transform 1 0 25116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_268
timestamp 1
transform 1 0 25760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_272
timestamp 1
transform 1 0 26128 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_276
timestamp 1
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_281
timestamp 1
transform 1 0 26956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_290
timestamp 1
transform 1 0 27784 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_296
timestamp 1
transform 1 0 28336 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1636968456
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1636968456
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_337
timestamp 1
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 1
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_395
timestamp 1
transform 1 0 37444 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_416
timestamp 1
transform 1 0 39376 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_431
timestamp 1
transform 1 0 40756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_455
timestamp 1
transform 1 0 42964 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_473
timestamp 1
transform 1 0 44620 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_477
timestamp 1
transform 1 0 44988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_486
timestamp 1
transform 1 0 45816 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_498
timestamp 1
transform 1 0 46920 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_505
timestamp 1
transform 1 0 47564 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_515
timestamp 1
transform 1 0 48484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_519
timestamp 1
transform 1 0 48852 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_526
timestamp 1
transform 1 0 49496 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_544
timestamp 1636968456
transform 1 0 51152 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_556
timestamp 1
transform 1 0 52256 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_561
timestamp 1636968456
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_573
timestamp 1
transform 1 0 53820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_579
timestamp 1
transform 1 0 54372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_583
timestamp 1
transform 1 0 54740 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_604
timestamp 1636968456
transform 1 0 56672 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_617
timestamp 1636968456
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_629
timestamp 1636968456
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_641
timestamp 1636968456
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_653
timestamp 1636968456
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_665
timestamp 1
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_671
timestamp 1
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_673
timestamp 1636968456
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_685
timestamp 1636968456
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_697
timestamp 1636968456
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_709
timestamp 1636968456
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_721
timestamp 1
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_727
timestamp 1
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_729
timestamp 1636968456
transform 1 0 68172 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_741
timestamp 1636968456
transform 1 0 69276 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_753
timestamp 1636968456
transform 1 0 70380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_765
timestamp 1636968456
transform 1 0 71484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_777
timestamp 1
transform 1 0 72588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_783
timestamp 1
transform 1 0 73140 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_785
timestamp 1636968456
transform 1 0 73324 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_797
timestamp 1636968456
transform 1 0 74428 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_809
timestamp 1636968456
transform 1 0 75532 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_821
timestamp 1636968456
transform 1 0 76636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_833
timestamp 1
transform 1 0 77740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_839
timestamp 1
transform 1 0 78292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_841
timestamp 1
transform 1 0 78476 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_8
timestamp 1636968456
transform 1 0 1840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_20
timestamp 1
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1636968456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1636968456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1636968456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_65
timestamp 1
transform 1 0 7084 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_73
timestamp 1
transform 1 0 7820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 1
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1636968456
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1636968456
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_109
timestamp 1
transform 1 0 11132 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_115
timestamp 1
transform 1 0 11684 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_125
timestamp 1
transform 1 0 12604 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_135
timestamp 1
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 1
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_152
timestamp 1
transform 1 0 15088 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1636968456
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1636968456
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_208
timestamp 1
transform 1 0 20240 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_224
timestamp 1
transform 1 0 21712 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_232
timestamp 1
transform 1 0 22448 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_241
timestamp 1
transform 1 0 23276 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_249
timestamp 1
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_253
timestamp 1
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_261
timestamp 1
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_269
timestamp 1
transform 1 0 25852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_292
timestamp 1
transform 1 0 27968 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_300
timestamp 1
transform 1 0 28704 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_331
timestamp 1
transform 1 0 31556 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_339
timestamp 1
transform 1 0 32292 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_353
timestamp 1
transform 1 0 33580 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_362
timestamp 1
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_397
timestamp 1
transform 1 0 37628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_418
timestamp 1
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_441
timestamp 1
transform 1 0 41676 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_471
timestamp 1
transform 1 0 44436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_475
timestamp 1
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_477
timestamp 1
transform 1 0 44988 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_498
timestamp 1636968456
transform 1 0 46920 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_510
timestamp 1636968456
transform 1 0 48024 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_522
timestamp 1
transform 1 0 49128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_526
timestamp 1
transform 1 0 49496 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_531
timestamp 1
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_542
timestamp 1636968456
transform 1 0 50968 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_554
timestamp 1636968456
transform 1 0 52072 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_568
timestamp 1
transform 1 0 53360 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_576
timestamp 1
transform 1 0 54096 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_585
timestamp 1
transform 1 0 54924 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_600
timestamp 1636968456
transform 1 0 56304 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_612
timestamp 1636968456
transform 1 0 57408 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_624
timestamp 1636968456
transform 1 0 58512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_636
timestamp 1
transform 1 0 59616 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_645
timestamp 1636968456
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_657
timestamp 1636968456
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_669
timestamp 1636968456
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_681
timestamp 1636968456
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_693
timestamp 1
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_699
timestamp 1
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_701
timestamp 1636968456
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_713
timestamp 1636968456
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_725
timestamp 1636968456
transform 1 0 67804 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_737
timestamp 1636968456
transform 1 0 68908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_749
timestamp 1
transform 1 0 70012 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_755
timestamp 1
transform 1 0 70564 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_757
timestamp 1636968456
transform 1 0 70748 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_769
timestamp 1636968456
transform 1 0 71852 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_781
timestamp 1636968456
transform 1 0 72956 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_793
timestamp 1636968456
transform 1 0 74060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_805
timestamp 1
transform 1 0 75164 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_811
timestamp 1
transform 1 0 75716 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_813
timestamp 1636968456
transform 1 0 75900 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_825
timestamp 1636968456
transform 1 0 77004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_837
timestamp 1
transform 1 0 78108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_841
timestamp 1
transform 1 0 78476 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_8
timestamp 1636968456
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_20
timestamp 1636968456
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_32
timestamp 1636968456
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_44
timestamp 1636968456
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1636968456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1636968456
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_102
timestamp 1
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_133
timestamp 1
transform 1 0 13340 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_164
timestamp 1
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_169
timestamp 1
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_186
timestamp 1636968456
transform 1 0 18216 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_198
timestamp 1
transform 1 0 19320 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_206
timestamp 1
transform 1 0 20056 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_212
timestamp 1
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_218
timestamp 1
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1636968456
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_237
timestamp 1
transform 1 0 22908 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_258
timestamp 1
transform 1 0 24840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_272
timestamp 1
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_281
timestamp 1
transform 1 0 26956 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_287
timestamp 1
transform 1 0 27508 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_291
timestamp 1
transform 1 0 27876 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_295
timestamp 1
transform 1 0 28244 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_301
timestamp 1636968456
transform 1 0 28796 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_313
timestamp 1636968456
transform 1 0 29900 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_325
timestamp 1
transform 1 0 31004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_333
timestamp 1
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_344
timestamp 1636968456
transform 1 0 32752 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_380
timestamp 1636968456
transform 1 0 36064 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1636968456
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 1636968456
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 1636968456
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_429
timestamp 1636968456
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_441
timestamp 1
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_447
timestamp 1
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_449
timestamp 1636968456
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_461
timestamp 1636968456
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_473
timestamp 1
transform 1 0 44620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_519
timestamp 1
transform 1 0 48852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_524
timestamp 1
transform 1 0 49312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_567
timestamp 1
transform 1 0 53268 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_599
timestamp 1
transform 1 0 56212 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_607
timestamp 1
transform 1 0 56948 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_619
timestamp 1636968456
transform 1 0 58052 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_631
timestamp 1636968456
transform 1 0 59156 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_643
timestamp 1636968456
transform 1 0 60260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_655
timestamp 1636968456
transform 1 0 61364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_667
timestamp 1
transform 1 0 62468 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_671
timestamp 1
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_673
timestamp 1636968456
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_685
timestamp 1636968456
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_697
timestamp 1636968456
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_709
timestamp 1636968456
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_721
timestamp 1
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_727
timestamp 1
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_729
timestamp 1636968456
transform 1 0 68172 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_741
timestamp 1636968456
transform 1 0 69276 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_753
timestamp 1636968456
transform 1 0 70380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_765
timestamp 1636968456
transform 1 0 71484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_777
timestamp 1
transform 1 0 72588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_783
timestamp 1
transform 1 0 73140 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_785
timestamp 1636968456
transform 1 0 73324 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_797
timestamp 1636968456
transform 1 0 74428 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_809
timestamp 1636968456
transform 1 0 75532 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_821
timestamp 1636968456
transform 1 0 76636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_833
timestamp 1
transform 1 0 77740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_839
timestamp 1
transform 1 0 78292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_841
timestamp 1
transform 1 0 78476 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1636968456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1636968456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1636968456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1636968456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1636968456
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1636968456
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_97
timestamp 1
transform 1 0 10028 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_116
timestamp 1
transform 1 0 11776 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_129
timestamp 1
transform 1 0 12972 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1636968456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1636968456
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1636968456
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_177
timestamp 1
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_197
timestamp 1
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_205
timestamp 1
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_217
timestamp 1636968456
transform 1 0 21068 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_229
timestamp 1
transform 1 0 22172 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_253
timestamp 1
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_261
timestamp 1
transform 1 0 25116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_280
timestamp 1
transform 1 0 26864 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_291
timestamp 1
transform 1 0 27876 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_300
timestamp 1
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1636968456
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1
transform 1 0 30636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_329
timestamp 1
transform 1 0 31372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_353
timestamp 1
transform 1 0 33580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_361
timestamp 1
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1636968456
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_377
timestamp 1
transform 1 0 35788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_403
timestamp 1
transform 1 0 38180 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_413
timestamp 1
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_419
timestamp 1
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_421
timestamp 1636968456
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_433
timestamp 1
transform 1 0 40940 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_454
timestamp 1
transform 1 0 42872 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_477
timestamp 1
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_487
timestamp 1
transform 1 0 45908 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_531
timestamp 1
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_550
timestamp 1
transform 1 0 51704 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_587
timestamp 1
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_589
timestamp 1
transform 1 0 55292 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_618
timestamp 1636968456
transform 1 0 57960 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_630
timestamp 1636968456
transform 1 0 59064 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_642
timestamp 1
transform 1 0 60168 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_645
timestamp 1636968456
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_657
timestamp 1636968456
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_669
timestamp 1636968456
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_681
timestamp 1636968456
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_693
timestamp 1
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_699
timestamp 1
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_701
timestamp 1636968456
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_713
timestamp 1636968456
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_725
timestamp 1636968456
transform 1 0 67804 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_737
timestamp 1636968456
transform 1 0 68908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_749
timestamp 1
transform 1 0 70012 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_755
timestamp 1
transform 1 0 70564 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_757
timestamp 1636968456
transform 1 0 70748 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_769
timestamp 1636968456
transform 1 0 71852 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_781
timestamp 1636968456
transform 1 0 72956 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_793
timestamp 1636968456
transform 1 0 74060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_805
timestamp 1
transform 1 0 75164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_811
timestamp 1
transform 1 0 75716 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_813
timestamp 1636968456
transform 1 0 75900 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_825
timestamp 1636968456
transform 1 0 77004 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_837
timestamp 1
transform 1 0 78108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_841
timestamp 1
transform 1 0 78476 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1636968456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1636968456
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1636968456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1636968456
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_81
timestamp 1
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_89
timestamp 1
transform 1 0 9292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 1
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_119
timestamp 1
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_147
timestamp 1
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_151
timestamp 1
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_169
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_201
timestamp 1
transform 1 0 19596 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_218
timestamp 1
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1636968456
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_237
timestamp 1
transform 1 0 22908 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_247
timestamp 1636968456
transform 1 0 23828 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_259
timestamp 1636968456
transform 1 0 24932 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_271
timestamp 1
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_281
timestamp 1
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_299
timestamp 1
transform 1 0 28612 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_303
timestamp 1
transform 1 0 28980 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_339
timestamp 1
transform 1 0 32292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_359
timestamp 1
transform 1 0 34132 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_367
timestamp 1636968456
transform 1 0 34868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_379
timestamp 1
transform 1 0 35972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_383
timestamp 1
transform 1 0 36340 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_393
timestamp 1
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_427
timestamp 1
transform 1 0 40388 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_433
timestamp 1
transform 1 0 40940 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_442
timestamp 1
transform 1 0 41768 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_451
timestamp 1
transform 1 0 42596 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_464
timestamp 1
transform 1 0 43792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_472
timestamp 1
transform 1 0 44528 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_484
timestamp 1
transform 1 0 45632 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_494
timestamp 1
transform 1 0 46552 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_502
timestamp 1
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_505
timestamp 1
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_517
timestamp 1636968456
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_533
timestamp 1
transform 1 0 50140 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_539
timestamp 1636968456
transform 1 0 50692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_551
timestamp 1
transform 1 0 51796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_559
timestamp 1
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_561
timestamp 1
transform 1 0 52716 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_569
timestamp 1
transform 1 0 53452 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_581
timestamp 1636968456
transform 1 0 54556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_593
timestamp 1636968456
transform 1 0 55660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_605
timestamp 1
transform 1 0 56764 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_613
timestamp 1
transform 1 0 57500 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_617
timestamp 1636968456
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_629
timestamp 1636968456
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_641
timestamp 1636968456
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_653
timestamp 1636968456
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_665
timestamp 1
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_671
timestamp 1
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_673
timestamp 1636968456
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_685
timestamp 1636968456
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_697
timestamp 1636968456
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_709
timestamp 1636968456
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_721
timestamp 1
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_727
timestamp 1
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_729
timestamp 1636968456
transform 1 0 68172 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_741
timestamp 1636968456
transform 1 0 69276 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_753
timestamp 1636968456
transform 1 0 70380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_765
timestamp 1636968456
transform 1 0 71484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_777
timestamp 1
transform 1 0 72588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_783
timestamp 1
transform 1 0 73140 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_785
timestamp 1636968456
transform 1 0 73324 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_797
timestamp 1636968456
transform 1 0 74428 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_809
timestamp 1636968456
transform 1 0 75532 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_821
timestamp 1636968456
transform 1 0 76636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_833
timestamp 1
transform 1 0 77740 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_841
timestamp 1
transform 1 0 78476 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1636968456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1636968456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1636968456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1636968456
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1636968456
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1636968456
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_97
timestamp 1
transform 1 0 10028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_122
timestamp 1
transform 1 0 12328 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_126
timestamp 1
transform 1 0 12696 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_136
timestamp 1
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_141
timestamp 1
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_173
timestamp 1
transform 1 0 17020 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_177
timestamp 1
transform 1 0 17388 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_199
timestamp 1
transform 1 0 19412 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_218
timestamp 1
transform 1 0 21160 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_226
timestamp 1636968456
transform 1 0 21896 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_238
timestamp 1636968456
transform 1 0 23000 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1636968456
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_265
timestamp 1
transform 1 0 25484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_272
timestamp 1
transform 1 0 26128 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_289
timestamp 1
transform 1 0 27692 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_297
timestamp 1
transform 1 0 28428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_305
timestamp 1
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_309
timestamp 1
transform 1 0 29532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_318
timestamp 1
transform 1 0 30360 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_323
timestamp 1
transform 1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_356
timestamp 1
transform 1 0 33856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_372
timestamp 1
transform 1 0 35328 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_375
timestamp 1
transform 1 0 35604 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_383
timestamp 1
transform 1 0 36340 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_397
timestamp 1
transform 1 0 37628 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_415
timestamp 1
transform 1 0 39284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 1
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_464
timestamp 1
transform 1 0 43792 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_477
timestamp 1
transform 1 0 44988 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_483
timestamp 1
transform 1 0 45540 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_493
timestamp 1
transform 1 0 46460 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_504
timestamp 1
transform 1 0 47472 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_515
timestamp 1636968456
transform 1 0 48484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_527
timestamp 1
transform 1 0 49588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_531
timestamp 1
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_533
timestamp 1636968456
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_545
timestamp 1
transform 1 0 51244 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_552
timestamp 1
transform 1 0 51888 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_560
timestamp 1
transform 1 0 52624 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_569
timestamp 1
transform 1 0 53452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_573
timestamp 1
transform 1 0 53820 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_582
timestamp 1
transform 1 0 54648 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_589
timestamp 1636968456
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_601
timestamp 1636968456
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_613
timestamp 1636968456
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_625
timestamp 1636968456
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_637
timestamp 1
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_643
timestamp 1
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_645
timestamp 1636968456
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_657
timestamp 1636968456
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_669
timestamp 1636968456
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_681
timestamp 1636968456
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_693
timestamp 1
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_699
timestamp 1
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_701
timestamp 1636968456
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_713
timestamp 1636968456
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_725
timestamp 1636968456
transform 1 0 67804 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_737
timestamp 1636968456
transform 1 0 68908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_749
timestamp 1
transform 1 0 70012 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_755
timestamp 1
transform 1 0 70564 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_757
timestamp 1636968456
transform 1 0 70748 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_769
timestamp 1636968456
transform 1 0 71852 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_781
timestamp 1636968456
transform 1 0 72956 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_793
timestamp 1636968456
transform 1 0 74060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_805
timestamp 1
transform 1 0 75164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_811
timestamp 1
transform 1 0 75716 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_813
timestamp 1636968456
transform 1 0 75900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_825
timestamp 1636968456
transform 1 0 77004 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_837
timestamp 1
transform 1 0 78108 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_841
timestamp 1
transform 1 0 78476 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1636968456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1636968456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1636968456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1636968456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1636968456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1636968456
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1636968456
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_96
timestamp 1636968456
transform 1 0 9936 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_108
timestamp 1
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1636968456
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_125
timestamp 1
transform 1 0 12604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_133
timestamp 1
transform 1 0 13340 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_144
timestamp 1636968456
transform 1 0 14352 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_156
timestamp 1636968456
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1636968456
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_181
timestamp 1
transform 1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_189
timestamp 1
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_195
timestamp 1
transform 1 0 19044 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_203
timestamp 1
transform 1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_213
timestamp 1
transform 1 0 20700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_225
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_248
timestamp 1
transform 1 0 23920 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_255
timestamp 1
transform 1 0 24564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_259
timestamp 1
transform 1 0 24932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_281
timestamp 1
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_289
timestamp 1
transform 1 0 27692 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_309
timestamp 1
transform 1 0 29532 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_317
timestamp 1
transform 1 0 30268 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_324
timestamp 1636968456
transform 1 0 30912 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_344
timestamp 1
transform 1 0 32752 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_352
timestamp 1
transform 1 0 33488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_373
timestamp 1
transform 1 0 35420 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_383
timestamp 1
transform 1 0 36340 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_401
timestamp 1
transform 1 0 37996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_404
timestamp 1
transform 1 0 38272 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_412
timestamp 1
transform 1 0 39008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_422
timestamp 1
transform 1 0 39928 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_473
timestamp 1
transform 1 0 44620 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_479
timestamp 1
transform 1 0 45172 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_500
timestamp 1
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_505
timestamp 1
transform 1 0 47564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_509
timestamp 1
transform 1 0 47932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_530
timestamp 1
transform 1 0 49864 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_548
timestamp 1
transform 1 0 51520 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_559
timestamp 1
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_561
timestamp 1
transform 1 0 52716 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_578
timestamp 1
transform 1 0 54280 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_604
timestamp 1636968456
transform 1 0 56672 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_617
timestamp 1636968456
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_629
timestamp 1636968456
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_641
timestamp 1636968456
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_653
timestamp 1636968456
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_665
timestamp 1
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_671
timestamp 1
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_673
timestamp 1636968456
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_685
timestamp 1636968456
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_697
timestamp 1636968456
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_709
timestamp 1636968456
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_721
timestamp 1
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_727
timestamp 1
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_729
timestamp 1636968456
transform 1 0 68172 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_741
timestamp 1636968456
transform 1 0 69276 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_753
timestamp 1636968456
transform 1 0 70380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_765
timestamp 1636968456
transform 1 0 71484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_777
timestamp 1
transform 1 0 72588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_783
timestamp 1
transform 1 0 73140 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_785
timestamp 1636968456
transform 1 0 73324 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_797
timestamp 1636968456
transform 1 0 74428 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_809
timestamp 1636968456
transform 1 0 75532 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_821
timestamp 1636968456
transform 1 0 76636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_833
timestamp 1
transform 1 0 77740 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_839
timestamp 1
transform 1 0 78292 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_841
timestamp 1
transform 1 0 78476 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1636968456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1636968456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1636968456
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_53
timestamp 1
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_61
timestamp 1
transform 1 0 6716 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_85
timestamp 1
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_100
timestamp 1636968456
transform 1 0 10304 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_112
timestamp 1636968456
transform 1 0 11408 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_124
timestamp 1636968456
transform 1 0 12512 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 1
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1636968456
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_153
timestamp 1
transform 1 0 15180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_157
timestamp 1
transform 1 0 15548 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_179
timestamp 1
transform 1 0 17572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_183
timestamp 1
transform 1 0 17940 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_193
timestamp 1
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_204
timestamp 1636968456
transform 1 0 19872 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_216
timestamp 1636968456
transform 1 0 20976 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_228
timestamp 1
transform 1 0 22080 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_242
timestamp 1
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1636968456
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1636968456
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1636968456
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_289
timestamp 1
transform 1 0 27692 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_293
timestamp 1
transform 1 0 28060 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_314
timestamp 1636968456
transform 1 0 29992 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_333
timestamp 1
transform 1 0 31740 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_344
timestamp 1
transform 1 0 32752 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_348
timestamp 1
transform 1 0 33120 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_365
timestamp 1
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_375
timestamp 1
transform 1 0 35604 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_389
timestamp 1
transform 1 0 36892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_428
timestamp 1
transform 1 0 40480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_433
timestamp 1
transform 1 0 40940 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_460
timestamp 1
transform 1 0 43424 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_471
timestamp 1
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_475
timestamp 1
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_477
timestamp 1636968456
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_489
timestamp 1636968456
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_501
timestamp 1
transform 1 0 47196 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_509
timestamp 1
transform 1 0 47932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_518
timestamp 1
transform 1 0 48760 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_533
timestamp 1
transform 1 0 50140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_556
timestamp 1
transform 1 0 52256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_585
timestamp 1
transform 1 0 54924 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_589
timestamp 1636968456
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_601
timestamp 1636968456
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_613
timestamp 1636968456
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_625
timestamp 1636968456
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_637
timestamp 1
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_643
timestamp 1
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_645
timestamp 1636968456
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_657
timestamp 1636968456
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_669
timestamp 1636968456
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_681
timestamp 1636968456
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_693
timestamp 1
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_699
timestamp 1
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_701
timestamp 1636968456
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_713
timestamp 1636968456
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_725
timestamp 1636968456
transform 1 0 67804 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_737
timestamp 1636968456
transform 1 0 68908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_749
timestamp 1
transform 1 0 70012 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_755
timestamp 1
transform 1 0 70564 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_757
timestamp 1636968456
transform 1 0 70748 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_769
timestamp 1636968456
transform 1 0 71852 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_781
timestamp 1636968456
transform 1 0 72956 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_793
timestamp 1636968456
transform 1 0 74060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_805
timestamp 1
transform 1 0 75164 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_811
timestamp 1
transform 1 0 75716 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_813
timestamp 1636968456
transform 1 0 75900 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_825
timestamp 1636968456
transform 1 0 77004 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_837
timestamp 1
transform 1 0 78108 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_841
timestamp 1
transform 1 0 78476 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1636968456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1636968456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1636968456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1636968456
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_57
timestamp 1
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_65
timestamp 1
transform 1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_74
timestamp 1636968456
transform 1 0 7912 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_86
timestamp 1
transform 1 0 9016 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_94
timestamp 1
transform 1 0 9752 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_106
timestamp 1
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_113
timestamp 1
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_117
timestamp 1
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_121
timestamp 1
transform 1 0 12236 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_125
timestamp 1
transform 1 0 12604 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_147
timestamp 1636968456
transform 1 0 14628 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_159
timestamp 1
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_169
timestamp 1
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_177
timestamp 1
transform 1 0 17388 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_203
timestamp 1636968456
transform 1 0 19780 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_215
timestamp 1
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1636968456
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1636968456
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_249
timestamp 1
transform 1 0 24012 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_275
timestamp 1
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_288
timestamp 1
transform 1 0 27600 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_292
timestamp 1
transform 1 0 27968 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_313
timestamp 1
transform 1 0 29900 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_350
timestamp 1636968456
transform 1 0 33304 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_362
timestamp 1636968456
transform 1 0 34408 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_374
timestamp 1
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_393
timestamp 1
transform 1 0 37260 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_408
timestamp 1
transform 1 0 38640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_416
timestamp 1
transform 1 0 39376 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_431
timestamp 1
transform 1 0 40756 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_441
timestamp 1
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_447
timestamp 1
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_451
timestamp 1
transform 1 0 42596 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_466
timestamp 1
transform 1 0 43976 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_476
timestamp 1636968456
transform 1 0 44896 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_488
timestamp 1636968456
transform 1 0 46000 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_500
timestamp 1
transform 1 0 47104 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_513
timestamp 1636968456
transform 1 0 48300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_525
timestamp 1636968456
transform 1 0 49404 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_537
timestamp 1
transform 1 0 50508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_541
timestamp 1
transform 1 0 50876 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_546
timestamp 1636968456
transform 1 0 51336 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_558
timestamp 1
transform 1 0 52440 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_561
timestamp 1636968456
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_573
timestamp 1636968456
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_585
timestamp 1636968456
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_597
timestamp 1636968456
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_609
timestamp 1
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_615
timestamp 1
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_617
timestamp 1636968456
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_629
timestamp 1636968456
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_641
timestamp 1636968456
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_653
timestamp 1636968456
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_665
timestamp 1
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_671
timestamp 1
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_673
timestamp 1636968456
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_685
timestamp 1636968456
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_697
timestamp 1636968456
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_709
timestamp 1636968456
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_721
timestamp 1
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_727
timestamp 1
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_729
timestamp 1636968456
transform 1 0 68172 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_741
timestamp 1636968456
transform 1 0 69276 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_753
timestamp 1636968456
transform 1 0 70380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_765
timestamp 1636968456
transform 1 0 71484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_777
timestamp 1
transform 1 0 72588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_783
timestamp 1
transform 1 0 73140 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_785
timestamp 1636968456
transform 1 0 73324 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_797
timestamp 1636968456
transform 1 0 74428 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_809
timestamp 1636968456
transform 1 0 75532 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_821
timestamp 1636968456
transform 1 0 76636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_833
timestamp 1
transform 1 0 77740 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_839
timestamp 1
transform 1 0 78292 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_841
timestamp 1
transform 1 0 78476 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_7
timestamp 1636968456
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_19
timestamp 1
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1636968456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1636968456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_53
timestamp 1
transform 1 0 5980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_61
timestamp 1
transform 1 0 6716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_75
timestamp 1
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_85
timestamp 1
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_118
timestamp 1
transform 1 0 11960 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_131
timestamp 1
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_163
timestamp 1636968456
transform 1 0 16100 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_175
timestamp 1
transform 1 0 17204 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_191
timestamp 1
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1636968456
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1636968456
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1636968456
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1636968456
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1636968456
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1636968456
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_300
timestamp 1
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1636968456
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1
transform 1 0 30636 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_329
timestamp 1
transform 1 0 31372 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_359
timestamp 1
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_372
timestamp 1636968456
transform 1 0 35328 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_384
timestamp 1
transform 1 0 36432 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 1636968456
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_401
timestamp 1636968456
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_413
timestamp 1
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_419
timestamp 1
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 1636968456
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_433
timestamp 1
transform 1 0 40940 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_441
timestamp 1
transform 1 0 41676 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_450
timestamp 1636968456
transform 1 0 42504 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_462
timestamp 1636968456
transform 1 0 43608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_474
timestamp 1
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_477
timestamp 1
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_485
timestamp 1
transform 1 0 45724 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_507
timestamp 1
transform 1 0 47748 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_513
timestamp 1
transform 1 0 48300 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_525
timestamp 1
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_531
timestamp 1
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_548
timestamp 1
transform 1 0 51520 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_563
timestamp 1636968456
transform 1 0 52900 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_575
timestamp 1636968456
transform 1 0 54004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_587
timestamp 1
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_609
timestamp 1636968456
transform 1 0 57132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_621
timestamp 1636968456
transform 1 0 58236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_633
timestamp 1
transform 1 0 59340 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_641
timestamp 1
transform 1 0 60076 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_645
timestamp 1636968456
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_657
timestamp 1636968456
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_669
timestamp 1636968456
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_681
timestamp 1636968456
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_693
timestamp 1
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_699
timestamp 1
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_701
timestamp 1636968456
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_713
timestamp 1636968456
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_725
timestamp 1636968456
transform 1 0 67804 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_737
timestamp 1636968456
transform 1 0 68908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_749
timestamp 1
transform 1 0 70012 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_755
timestamp 1
transform 1 0 70564 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_757
timestamp 1636968456
transform 1 0 70748 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_769
timestamp 1636968456
transform 1 0 71852 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_781
timestamp 1636968456
transform 1 0 72956 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_793
timestamp 1636968456
transform 1 0 74060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_805
timestamp 1
transform 1 0 75164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_811
timestamp 1
transform 1 0 75716 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_813
timestamp 1636968456
transform 1 0 75900 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_825
timestamp 1636968456
transform 1 0 77004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_837
timestamp 1
transform 1 0 78108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_841
timestamp 1
transform 1 0 78476 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1636968456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1636968456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1636968456
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1636968456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_69
timestamp 1
transform 1 0 7452 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_93
timestamp 1
transform 1 0 9660 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_97
timestamp 1
transform 1 0 10028 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_104
timestamp 1
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_113
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_141
timestamp 1
transform 1 0 14076 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_151
timestamp 1636968456
transform 1 0 14996 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_163
timestamp 1
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1636968456
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1636968456
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1636968456
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 1636968456
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_247
timestamp 1636968456
transform 1 0 23828 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_259
timestamp 1636968456
transform 1 0 24932 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_271
timestamp 1
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_281
timestamp 1
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_302
timestamp 1636968456
transform 1 0 28888 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_314
timestamp 1636968456
transform 1 0 29992 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_326
timestamp 1
transform 1 0 31096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_334
timestamp 1
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_372
timestamp 1636968456
transform 1 0 35328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_408
timestamp 1
transform 1 0 38640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_416
timestamp 1
transform 1 0 39376 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_426
timestamp 1
transform 1 0 40296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_444
timestamp 1
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_449
timestamp 1
transform 1 0 42412 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_457
timestamp 1
transform 1 0 43148 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_466
timestamp 1636968456
transform 1 0 43976 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_478
timestamp 1636968456
transform 1 0 45080 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_490
timestamp 1
transform 1 0 46184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_502
timestamp 1
transform 1 0 47288 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_505
timestamp 1
transform 1 0 47564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_532
timestamp 1
transform 1 0 50048 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_536
timestamp 1
transform 1 0 50416 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_557
timestamp 1
transform 1 0 52348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_581
timestamp 1
transform 1 0 54556 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_591
timestamp 1
transform 1 0 55476 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_610
timestamp 1
transform 1 0 57224 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_617
timestamp 1636968456
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_629
timestamp 1636968456
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_641
timestamp 1636968456
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_653
timestamp 1636968456
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_665
timestamp 1
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_671
timestamp 1
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_673
timestamp 1636968456
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_685
timestamp 1636968456
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_697
timestamp 1636968456
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_709
timestamp 1636968456
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_721
timestamp 1
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_727
timestamp 1
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_729
timestamp 1636968456
transform 1 0 68172 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_741
timestamp 1636968456
transform 1 0 69276 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_753
timestamp 1636968456
transform 1 0 70380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_765
timestamp 1636968456
transform 1 0 71484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_777
timestamp 1
transform 1 0 72588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_783
timestamp 1
transform 1 0 73140 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_785
timestamp 1636968456
transform 1 0 73324 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_797
timestamp 1636968456
transform 1 0 74428 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_809
timestamp 1636968456
transform 1 0 75532 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_821
timestamp 1636968456
transform 1 0 76636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_833
timestamp 1
transform 1 0 77740 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_839
timestamp 1
transform 1 0 78292 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_841
timestamp 1
transform 1 0 78476 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_7
timestamp 1636968456
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_19
timestamp 1
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1636968456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1636968456
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_53
timestamp 1
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_61
timestamp 1
transform 1 0 6716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_85
timestamp 1
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_93
timestamp 1
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_102
timestamp 1
transform 1 0 10488 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_110
timestamp 1
transform 1 0 11224 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_114
timestamp 1636968456
transform 1 0 11592 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_126
timestamp 1636968456
transform 1 0 12696 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_149
timestamp 1636968456
transform 1 0 14812 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_161
timestamp 1636968456
transform 1 0 15916 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_173
timestamp 1636968456
transform 1 0 17020 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_185
timestamp 1
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_193
timestamp 1
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1636968456
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1636968456
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1636968456
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1636968456
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 1
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1636968456
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1636968456
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1636968456
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 1636968456
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 1
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_332
timestamp 1636968456
transform 1 0 31648 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_344
timestamp 1636968456
transform 1 0 32752 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_356
timestamp 1
transform 1 0 33856 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_365
timestamp 1
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_374
timestamp 1
transform 1 0 35512 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_378
timestamp 1
transform 1 0 35880 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_399
timestamp 1
transform 1 0 37812 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_441
timestamp 1
transform 1 0 41676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_445
timestamp 1
transform 1 0 42044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_455
timestamp 1636968456
transform 1 0 42964 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_481
timestamp 1636968456
transform 1 0 45356 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_493
timestamp 1636968456
transform 1 0 46460 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_505
timestamp 1
transform 1 0 47564 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_513
timestamp 1
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_525
timestamp 1
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_531
timestamp 1
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_533
timestamp 1
transform 1 0 50140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_545
timestamp 1
transform 1 0 51244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_549
timestamp 1
transform 1 0 51612 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_558
timestamp 1
transform 1 0 52440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_568
timestamp 1
transform 1 0 53360 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_586
timestamp 1
transform 1 0 55016 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_606
timestamp 1636968456
transform 1 0 56856 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_618
timestamp 1636968456
transform 1 0 57960 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_630
timestamp 1636968456
transform 1 0 59064 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_642
timestamp 1
transform 1 0 60168 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_645
timestamp 1636968456
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_657
timestamp 1636968456
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_669
timestamp 1636968456
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_681
timestamp 1636968456
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_693
timestamp 1
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_699
timestamp 1
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_701
timestamp 1636968456
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_713
timestamp 1636968456
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_725
timestamp 1636968456
transform 1 0 67804 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_737
timestamp 1636968456
transform 1 0 68908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_749
timestamp 1
transform 1 0 70012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_755
timestamp 1
transform 1 0 70564 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_757
timestamp 1636968456
transform 1 0 70748 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_769
timestamp 1636968456
transform 1 0 71852 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_781
timestamp 1636968456
transform 1 0 72956 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_793
timestamp 1636968456
transform 1 0 74060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_805
timestamp 1
transform 1 0 75164 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_811
timestamp 1
transform 1 0 75716 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_813
timestamp 1636968456
transform 1 0 75900 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_825
timestamp 1636968456
transform 1 0 77004 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_837
timestamp 1
transform 1 0 78108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_841
timestamp 1
transform 1 0 78476 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_7
timestamp 1636968456
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_19
timestamp 1636968456
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_31
timestamp 1636968456
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_43
timestamp 1636968456
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1636968456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_69
timestamp 1
transform 1 0 7452 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_91
timestamp 1636968456
transform 1 0 9476 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_103
timestamp 1
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_113
timestamp 1
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_121
timestamp 1
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_143
timestamp 1636968456
transform 1 0 14260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_155
timestamp 1636968456
transform 1 0 15364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1636968456
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1636968456
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1636968456
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1636968456
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1636968456
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1636968456
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1636968456
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 1636968456
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 1
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1636968456
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1636968456
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_305
timestamp 1
transform 1 0 29164 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_332
timestamp 1
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1636968456
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_349
timestamp 1
transform 1 0 33212 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_355
timestamp 1
transform 1 0 33764 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_384
timestamp 1
transform 1 0 36432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_400
timestamp 1
transform 1 0 37904 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_424
timestamp 1636968456
transform 1 0 40112 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_436
timestamp 1636968456
transform 1 0 41216 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_449
timestamp 1636968456
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_461
timestamp 1636968456
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_482
timestamp 1
transform 1 0 45448 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_494
timestamp 1
transform 1 0 46552 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_502
timestamp 1
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_514
timestamp 1636968456
transform 1 0 48392 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_526
timestamp 1
transform 1 0 49496 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_546
timestamp 1636968456
transform 1 0 51336 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_558
timestamp 1
transform 1 0 52440 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_561
timestamp 1
transform 1 0 52716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_565
timestamp 1
transform 1 0 53084 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_568
timestamp 1636968456
transform 1 0 53360 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_580
timestamp 1
transform 1 0 54464 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_608
timestamp 1
transform 1 0 57040 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_617
timestamp 1636968456
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_629
timestamp 1636968456
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_641
timestamp 1636968456
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_653
timestamp 1636968456
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_665
timestamp 1
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_671
timestamp 1
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_673
timestamp 1636968456
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_685
timestamp 1636968456
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_697
timestamp 1636968456
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_709
timestamp 1636968456
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_721
timestamp 1
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_727
timestamp 1
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_729
timestamp 1636968456
transform 1 0 68172 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_741
timestamp 1636968456
transform 1 0 69276 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_753
timestamp 1636968456
transform 1 0 70380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_765
timestamp 1636968456
transform 1 0 71484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_777
timestamp 1
transform 1 0 72588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_783
timestamp 1
transform 1 0 73140 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_785
timestamp 1636968456
transform 1 0 73324 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_797
timestamp 1636968456
transform 1 0 74428 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_809
timestamp 1636968456
transform 1 0 75532 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_821
timestamp 1636968456
transform 1 0 76636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_833
timestamp 1
transform 1 0 77740 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_839
timestamp 1
transform 1 0 78292 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_841
timestamp 1
transform 1 0 78476 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_7
timestamp 1636968456
transform 1 0 1748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_19
timestamp 1
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1636968456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1636968456
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1636968456
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1636968456
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1636968456
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_97
timestamp 1
transform 1 0 10028 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_119
timestamp 1
transform 1 0 12052 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_125
timestamp 1
transform 1 0 12604 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_132
timestamp 1
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_141
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_151
timestamp 1636968456
transform 1 0 14996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_163
timestamp 1
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_167
timestamp 1
transform 1 0 16468 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_175
timestamp 1636968456
transform 1 0 17204 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_187
timestamp 1
transform 1 0 18308 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_191
timestamp 1
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1636968456
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1636968456
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1636968456
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 1636968456
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1636968456
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1636968456
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1636968456
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1636968456
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_301
timestamp 1
transform 1 0 28796 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_330
timestamp 1
transform 1 0 31464 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1636968456
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1636968456
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_389
timestamp 1
transform 1 0 36892 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_400
timestamp 1
transform 1 0 37904 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_405
timestamp 1
transform 1 0 38364 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_413
timestamp 1
transform 1 0 39100 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_416
timestamp 1
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 1636968456
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_433
timestamp 1
transform 1 0 40940 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_441
timestamp 1
transform 1 0 41676 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_460
timestamp 1636968456
transform 1 0 43424 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_472
timestamp 1
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_504
timestamp 1636968456
transform 1 0 47472 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_516
timestamp 1
transform 1 0 48576 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_530
timestamp 1
transform 1 0 49864 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_537
timestamp 1636968456
transform 1 0 50508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_549
timestamp 1636968456
transform 1 0 51612 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_579
timestamp 1
transform 1 0 54372 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_587
timestamp 1
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_589
timestamp 1636968456
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_601
timestamp 1636968456
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_613
timestamp 1636968456
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_625
timestamp 1636968456
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_637
timestamp 1
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_643
timestamp 1
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_645
timestamp 1636968456
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_657
timestamp 1636968456
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_669
timestamp 1636968456
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_681
timestamp 1636968456
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_693
timestamp 1
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_699
timestamp 1
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_701
timestamp 1636968456
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_713
timestamp 1636968456
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_725
timestamp 1636968456
transform 1 0 67804 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_737
timestamp 1636968456
transform 1 0 68908 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_749
timestamp 1
transform 1 0 70012 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_755
timestamp 1
transform 1 0 70564 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_757
timestamp 1636968456
transform 1 0 70748 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_769
timestamp 1636968456
transform 1 0 71852 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_781
timestamp 1636968456
transform 1 0 72956 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_793
timestamp 1636968456
transform 1 0 74060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_805
timestamp 1
transform 1 0 75164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_811
timestamp 1
transform 1 0 75716 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_813
timestamp 1636968456
transform 1 0 75900 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_825
timestamp 1636968456
transform 1 0 77004 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_837
timestamp 1
transform 1 0 78108 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_841
timestamp 1
transform 1 0 78476 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1636968456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1636968456
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1636968456
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1636968456
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1636968456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1636968456
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_81
timestamp 1
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_89
timestamp 1
transform 1 0 9292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_103
timestamp 1
transform 1 0 10580 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_115
timestamp 1636968456
transform 1 0 11684 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_127
timestamp 1
transform 1 0 12788 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_135
timestamp 1
transform 1 0 13524 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_158
timestamp 1
transform 1 0 15640 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 1
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1636968456
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1636968456
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1636968456
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1636968456
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 1636968456
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_281
timestamp 1
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_289
timestamp 1
transform 1 0 27692 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_322
timestamp 1636968456
transform 1 0 30728 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_334
timestamp 1
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_351
timestamp 1636968456
transform 1 0 33396 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_363
timestamp 1
transform 1 0 34500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_378
timestamp 1
transform 1 0 35880 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_384
timestamp 1
transform 1 0 36432 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_390
timestamp 1
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_393
timestamp 1
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_426
timestamp 1636968456
transform 1 0 40296 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_438
timestamp 1
transform 1 0 41400 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_446
timestamp 1
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_458
timestamp 1
transform 1 0 43240 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_466
timestamp 1636968456
transform 1 0 43976 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_478
timestamp 1636968456
transform 1 0 45080 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_490
timestamp 1636968456
transform 1 0 46184 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_502
timestamp 1
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_505
timestamp 1
transform 1 0 47564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_509
timestamp 1
transform 1 0 47932 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_536
timestamp 1
transform 1 0 50416 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_551
timestamp 1
transform 1 0 51796 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_559
timestamp 1
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_581
timestamp 1
transform 1 0 54556 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_591
timestamp 1
transform 1 0 55476 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_607
timestamp 1
transform 1 0 56948 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_615
timestamp 1
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_627
timestamp 1636968456
transform 1 0 58788 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_639
timestamp 1636968456
transform 1 0 59892 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_651
timestamp 1636968456
transform 1 0 60996 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_663
timestamp 1
transform 1 0 62100 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_671
timestamp 1
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_673
timestamp 1636968456
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_685
timestamp 1636968456
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_697
timestamp 1636968456
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_709
timestamp 1636968456
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_721
timestamp 1
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_727
timestamp 1
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_729
timestamp 1636968456
transform 1 0 68172 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_741
timestamp 1636968456
transform 1 0 69276 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_753
timestamp 1636968456
transform 1 0 70380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_765
timestamp 1636968456
transform 1 0 71484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_777
timestamp 1
transform 1 0 72588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_783
timestamp 1
transform 1 0 73140 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_785
timestamp 1636968456
transform 1 0 73324 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_797
timestamp 1636968456
transform 1 0 74428 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_809
timestamp 1636968456
transform 1 0 75532 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_821
timestamp 1636968456
transform 1 0 76636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_833
timestamp 1
transform 1 0 77740 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_839
timestamp 1
transform 1 0 78292 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_841
timestamp 1
transform 1 0 78476 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_3
timestamp 1
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_18
timestamp 1
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_26
timestamp 1
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1636968456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1636968456
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1636968456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1636968456
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1636968456
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_97
timestamp 1
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_110
timestamp 1636968456
transform 1 0 11224 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_122
timestamp 1636968456
transform 1 0 12328 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_134
timestamp 1
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_149
timestamp 1636968456
transform 1 0 14812 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_161
timestamp 1
transform 1 0 15916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_165
timestamp 1
transform 1 0 16284 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_192
timestamp 1
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_199
timestamp 1636968456
transform 1 0 19412 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_211
timestamp 1636968456
transform 1 0 20516 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_223
timestamp 1636968456
transform 1 0 21620 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_235
timestamp 1636968456
transform 1 0 22724 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_247
timestamp 1
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1636968456
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1636968456
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1636968456
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 1636968456
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 1
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_329
timestamp 1636968456
transform 1 0 31372 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_341
timestamp 1
transform 1 0 32476 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_349
timestamp 1
transform 1 0 33212 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 1
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_365
timestamp 1
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_391
timestamp 1636968456
transform 1 0 37076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_403
timestamp 1636968456
transform 1 0 38180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_415
timestamp 1
transform 1 0 39284 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_419
timestamp 1
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_431
timestamp 1
transform 1 0 40756 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_437
timestamp 1
transform 1 0 41308 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_474
timestamp 1
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_484
timestamp 1
transform 1 0 45632 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_488
timestamp 1
transform 1 0 46000 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_494
timestamp 1
transform 1 0 46552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_529
timestamp 1
transform 1 0 49772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_533
timestamp 1
transform 1 0 50140 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_551
timestamp 1636968456
transform 1 0 51796 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_574
timestamp 1
transform 1 0 53912 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_583
timestamp 1
transform 1 0 54740 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_587
timestamp 1
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_625
timestamp 1636968456
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_637
timestamp 1
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_643
timestamp 1
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_645
timestamp 1636968456
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_657
timestamp 1636968456
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_669
timestamp 1636968456
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_681
timestamp 1636968456
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_693
timestamp 1
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_699
timestamp 1
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_701
timestamp 1636968456
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_713
timestamp 1636968456
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_725
timestamp 1636968456
transform 1 0 67804 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_737
timestamp 1636968456
transform 1 0 68908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_749
timestamp 1
transform 1 0 70012 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_755
timestamp 1
transform 1 0 70564 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_757
timestamp 1636968456
transform 1 0 70748 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_769
timestamp 1636968456
transform 1 0 71852 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_781
timestamp 1636968456
transform 1 0 72956 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_793
timestamp 1636968456
transform 1 0 74060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_805
timestamp 1
transform 1 0 75164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_811
timestamp 1
transform 1 0 75716 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_813
timestamp 1636968456
transform 1 0 75900 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_825
timestamp 1636968456
transform 1 0 77004 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_837
timestamp 1
transform 1 0 78108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_841
timestamp 1
transform 1 0 78476 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_3
timestamp 1
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_14
timestamp 1636968456
transform 1 0 2392 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_26
timestamp 1636968456
transform 1 0 3496 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_38
timestamp 1636968456
transform 1 0 4600 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_50
timestamp 1
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1636968456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1636968456
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_81
timestamp 1
transform 1 0 8556 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_109
timestamp 1
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1636968456
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1636968456
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_137
timestamp 1
transform 1 0 13708 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1636968456
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_169
timestamp 1
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_227
timestamp 1636968456
transform 1 0 21988 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_239
timestamp 1636968456
transform 1 0 23092 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_251
timestamp 1636968456
transform 1 0 24196 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_263
timestamp 1636968456
transform 1 0 25300 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_275
timestamp 1
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1636968456
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1636968456
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_305
timestamp 1
transform 1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_313
timestamp 1
transform 1 0 29900 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_339
timestamp 1
transform 1 0 32292 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_343
timestamp 1
transform 1 0 32660 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_379
timestamp 1
transform 1 0 35972 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_404
timestamp 1
transform 1 0 38272 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_410
timestamp 1
transform 1 0 38824 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_435
timestamp 1636968456
transform 1 0 41124 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 1
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_460
timestamp 1
transform 1 0 43424 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_475
timestamp 1
transform 1 0 44804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_483
timestamp 1
transform 1 0 45540 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_496
timestamp 1
transform 1 0 46736 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_505
timestamp 1
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_517
timestamp 1
transform 1 0 48668 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_533
timestamp 1
transform 1 0 50140 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_545
timestamp 1636968456
transform 1 0 51244 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_557
timestamp 1
transform 1 0 52348 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_561
timestamp 1636968456
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_573
timestamp 1
transform 1 0 53820 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_577
timestamp 1
transform 1 0 54188 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_585
timestamp 1636968456
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_597
timestamp 1636968456
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_609
timestamp 1
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_615
timestamp 1
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_617
timestamp 1636968456
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_629
timestamp 1636968456
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_641
timestamp 1636968456
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_653
timestamp 1636968456
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_665
timestamp 1
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_671
timestamp 1
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_673
timestamp 1636968456
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_685
timestamp 1636968456
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_697
timestamp 1636968456
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_709
timestamp 1636968456
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_721
timestamp 1
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_727
timestamp 1
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_729
timestamp 1636968456
transform 1 0 68172 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_741
timestamp 1636968456
transform 1 0 69276 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_753
timestamp 1636968456
transform 1 0 70380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_765
timestamp 1636968456
transform 1 0 71484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_777
timestamp 1
transform 1 0 72588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_783
timestamp 1
transform 1 0 73140 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_785
timestamp 1636968456
transform 1 0 73324 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_797
timestamp 1636968456
transform 1 0 74428 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_809
timestamp 1636968456
transform 1 0 75532 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_821
timestamp 1636968456
transform 1 0 76636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_833
timestamp 1
transform 1 0 77740 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_841
timestamp 1
transform 1 0 78476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_3
timestamp 1
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_7
timestamp 1
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_11
timestamp 1636968456
transform 1 0 2116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_23
timestamp 1
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1636968456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1636968456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1636968456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1636968456
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_92
timestamp 1
transform 1 0 9568 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_109
timestamp 1
transform 1 0 11132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_113
timestamp 1
transform 1 0 11500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_141
timestamp 1
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_167
timestamp 1
transform 1 0 16468 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_175
timestamp 1
transform 1 0 17204 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_180
timestamp 1636968456
transform 1 0 17664 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_192
timestamp 1
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1636968456
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_209
timestamp 1
transform 1 0 20332 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_218
timestamp 1636968456
transform 1 0 21160 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_230
timestamp 1636968456
transform 1 0 22264 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_242
timestamp 1
transform 1 0 23368 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_250
timestamp 1
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1636968456
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1636968456
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1636968456
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1636968456
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1636968456
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_321
timestamp 1
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_325
timestamp 1
transform 1 0 31004 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1636968456
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_345
timestamp 1
transform 1 0 32844 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_349
timestamp 1
transform 1 0 33212 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1636968456
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_377
timestamp 1
transform 1 0 35788 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_383
timestamp 1636968456
transform 1 0 36340 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_395
timestamp 1636968456
transform 1 0 37444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_407
timestamp 1636968456
transform 1 0 38548 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 1
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_428
timestamp 1636968456
transform 1 0 40480 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_440
timestamp 1
transform 1 0 41584 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_453
timestamp 1
transform 1 0 42780 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_461
timestamp 1
transform 1 0 43516 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_472
timestamp 1
transform 1 0 44528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_477
timestamp 1
transform 1 0 44988 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_481
timestamp 1
transform 1 0 45356 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_505
timestamp 1
transform 1 0 47564 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_511
timestamp 1
transform 1 0 48116 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_533
timestamp 1
transform 1 0 50140 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_539
timestamp 1
transform 1 0 50692 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_560
timestamp 1
transform 1 0 52624 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_569
timestamp 1636968456
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_581
timestamp 1
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_587
timestamp 1
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_596
timestamp 1636968456
transform 1 0 55936 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_608
timestamp 1636968456
transform 1 0 57040 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_620
timestamp 1636968456
transform 1 0 58144 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_632
timestamp 1636968456
transform 1 0 59248 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_645
timestamp 1636968456
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_657
timestamp 1636968456
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_669
timestamp 1636968456
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_681
timestamp 1636968456
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_693
timestamp 1
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_699
timestamp 1
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_701
timestamp 1636968456
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_713
timestamp 1636968456
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_725
timestamp 1636968456
transform 1 0 67804 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_737
timestamp 1636968456
transform 1 0 68908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_749
timestamp 1
transform 1 0 70012 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_755
timestamp 1
transform 1 0 70564 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_757
timestamp 1636968456
transform 1 0 70748 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_769
timestamp 1636968456
transform 1 0 71852 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_781
timestamp 1636968456
transform 1 0 72956 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_793
timestamp 1636968456
transform 1 0 74060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_805
timestamp 1
transform 1 0 75164 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_811
timestamp 1
transform 1 0 75716 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_813
timestamp 1636968456
transform 1 0 75900 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_825
timestamp 1636968456
transform 1 0 77004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_837
timestamp 1
transform 1 0 78108 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_841
timestamp 1
transform 1 0 78476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_3
timestamp 1
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_14
timestamp 1636968456
transform 1 0 2392 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_26
timestamp 1636968456
transform 1 0 3496 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_38
timestamp 1636968456
transform 1 0 4600 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_50
timestamp 1
transform 1 0 5704 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1636968456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_69
timestamp 1
transform 1 0 7452 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_102
timestamp 1
transform 1 0 10488 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_113
timestamp 1
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_121
timestamp 1
transform 1 0 12236 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_125
timestamp 1
transform 1 0 12604 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_159
timestamp 1
transform 1 0 15732 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_169
timestamp 1
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_183
timestamp 1636968456
transform 1 0 17940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_195
timestamp 1
transform 1 0 19044 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_203
timestamp 1
transform 1 0 19780 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_209
timestamp 1636968456
transform 1 0 20332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_221
timestamp 1
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1636968456
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1636968456
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1636968456
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1636968456
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1636968456
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_293
timestamp 1
transform 1 0 28060 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_327
timestamp 1
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1636968456
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_349
timestamp 1
transform 1 0 33212 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_372
timestamp 1636968456
transform 1 0 35328 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_393
timestamp 1
transform 1 0 37260 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_410
timestamp 1636968456
transform 1 0 38824 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_422
timestamp 1636968456
transform 1 0 39928 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_434
timestamp 1
transform 1 0 41032 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_442
timestamp 1
transform 1 0 41768 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_447
timestamp 1
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_470
timestamp 1
transform 1 0 44344 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_480
timestamp 1636968456
transform 1 0 45264 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_492
timestamp 1636968456
transform 1 0 46368 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_505
timestamp 1
transform 1 0 47564 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_534
timestamp 1
transform 1 0 50232 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_547
timestamp 1
transform 1 0 51428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_551
timestamp 1
transform 1 0 51796 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_561
timestamp 1
transform 1 0 52716 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_584
timestamp 1
transform 1 0 54832 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_594
timestamp 1636968456
transform 1 0 55752 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_606
timestamp 1
transform 1 0 56856 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_614
timestamp 1
transform 1 0 57592 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_617
timestamp 1636968456
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_629
timestamp 1636968456
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_641
timestamp 1636968456
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_653
timestamp 1636968456
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_665
timestamp 1
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_671
timestamp 1
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_673
timestamp 1636968456
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_685
timestamp 1636968456
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_697
timestamp 1636968456
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_709
timestamp 1636968456
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_721
timestamp 1
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_727
timestamp 1
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_729
timestamp 1636968456
transform 1 0 68172 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_741
timestamp 1636968456
transform 1 0 69276 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_753
timestamp 1636968456
transform 1 0 70380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_765
timestamp 1636968456
transform 1 0 71484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_777
timestamp 1
transform 1 0 72588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_783
timestamp 1
transform 1 0 73140 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_785
timestamp 1636968456
transform 1 0 73324 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_797
timestamp 1636968456
transform 1 0 74428 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_809
timestamp 1636968456
transform 1 0 75532 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_821
timestamp 1636968456
transform 1 0 76636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_833
timestamp 1
transform 1 0 77740 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_839
timestamp 1
transform 1 0 78292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_841
timestamp 1
transform 1 0 78476 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_3
timestamp 1
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_14
timestamp 1636968456
transform 1 0 2392 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_26
timestamp 1
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1636968456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1636968456
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1636968456
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1636968456
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1636968456
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1636968456
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_121
timestamp 1
transform 1 0 12236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_125
timestamp 1
transform 1 0 12604 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_135
timestamp 1
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_150
timestamp 1
transform 1 0 14904 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_156
timestamp 1
transform 1 0 15456 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_192
timestamp 1
transform 1 0 18768 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_219
timestamp 1636968456
transform 1 0 21252 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_231
timestamp 1636968456
transform 1 0 22356 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_243
timestamp 1
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1636968456
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1636968456
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_277
timestamp 1
transform 1 0 26588 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_293
timestamp 1636968456
transform 1 0 28060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_305
timestamp 1
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1636968456
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_321
timestamp 1
transform 1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_332
timestamp 1636968456
transform 1 0 31648 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_344
timestamp 1636968456
transform 1 0 32752 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_356
timestamp 1
transform 1 0 33856 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_372
timestamp 1
transform 1 0 35328 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_397
timestamp 1
transform 1 0 37628 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_421
timestamp 1
transform 1 0 39836 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_429
timestamp 1
transform 1 0 40572 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_446
timestamp 1
transform 1 0 42136 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_464
timestamp 1636968456
transform 1 0 43792 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_477
timestamp 1636968456
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_489
timestamp 1636968456
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_501
timestamp 1636968456
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_513
timestamp 1636968456
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_525
timestamp 1
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_531
timestamp 1
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_533
timestamp 1636968456
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_545
timestamp 1
transform 1 0 51244 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_554
timestamp 1
transform 1 0 52072 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_562
timestamp 1
transform 1 0 52808 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_573
timestamp 1636968456
transform 1 0 53820 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_585
timestamp 1
transform 1 0 54924 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_609
timestamp 1636968456
transform 1 0 57132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_621
timestamp 1636968456
transform 1 0 58236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_633
timestamp 1
transform 1 0 59340 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_641
timestamp 1
transform 1 0 60076 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_645
timestamp 1636968456
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_657
timestamp 1636968456
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_669
timestamp 1636968456
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_681
timestamp 1636968456
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_693
timestamp 1
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_699
timestamp 1
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_701
timestamp 1636968456
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_713
timestamp 1636968456
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_725
timestamp 1636968456
transform 1 0 67804 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_737
timestamp 1636968456
transform 1 0 68908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_749
timestamp 1
transform 1 0 70012 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_755
timestamp 1
transform 1 0 70564 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_757
timestamp 1636968456
transform 1 0 70748 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_769
timestamp 1636968456
transform 1 0 71852 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_781
timestamp 1636968456
transform 1 0 72956 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_793
timestamp 1636968456
transform 1 0 74060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_805
timestamp 1
transform 1 0 75164 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_811
timestamp 1
transform 1 0 75716 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_813
timestamp 1636968456
transform 1 0 75900 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_825
timestamp 1636968456
transform 1 0 77004 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_837
timestamp 1
transform 1 0 78108 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_841
timestamp 1
transform 1 0 78476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_3
timestamp 1
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_14
timestamp 1636968456
transform 1 0 2392 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_26
timestamp 1636968456
transform 1 0 3496 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_38
timestamp 1636968456
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_50
timestamp 1
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1636968456
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1636968456
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1636968456
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1636968456
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1636968456
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1636968456
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_149
timestamp 1
transform 1 0 14812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_169
timestamp 1
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_183
timestamp 1636968456
transform 1 0 17940 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_195
timestamp 1
transform 1 0 19044 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_205
timestamp 1
transform 1 0 19964 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_247
timestamp 1636968456
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_259
timestamp 1636968456
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_271
timestamp 1
transform 1 0 26036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1636968456
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1636968456
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_305
timestamp 1
transform 1 0 29164 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_334
timestamp 1
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_337
timestamp 1
transform 1 0 32108 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_347
timestamp 1636968456
transform 1 0 33028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_359
timestamp 1
transform 1 0 34132 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_370
timestamp 1636968456
transform 1 0 35144 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_382
timestamp 1
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_390
timestamp 1
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_408
timestamp 1636968456
transform 1 0 38640 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_420
timestamp 1
transform 1 0 39744 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_428
timestamp 1
transform 1 0 40480 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_434
timestamp 1636968456
transform 1 0 41032 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_446
timestamp 1
transform 1 0 42136 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_449
timestamp 1
transform 1 0 42412 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_455
timestamp 1636968456
transform 1 0 42964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_467
timestamp 1
transform 1 0 44068 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_477
timestamp 1636968456
transform 1 0 44988 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_495
timestamp 1
transform 1 0 46644 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_501
timestamp 1
transform 1 0 47196 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_514
timestamp 1
transform 1 0 48392 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_522
timestamp 1
transform 1 0 49128 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_531
timestamp 1636968456
transform 1 0 49956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_552
timestamp 1
transform 1 0 51888 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_570
timestamp 1636968456
transform 1 0 53544 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_582
timestamp 1636968456
transform 1 0 54648 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_594
timestamp 1636968456
transform 1 0 55752 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_606
timestamp 1
transform 1 0 56856 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_614
timestamp 1
transform 1 0 57592 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_617
timestamp 1636968456
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_629
timestamp 1636968456
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_641
timestamp 1636968456
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_653
timestamp 1636968456
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_665
timestamp 1
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_671
timestamp 1
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_673
timestamp 1636968456
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_685
timestamp 1636968456
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_697
timestamp 1636968456
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_709
timestamp 1636968456
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_721
timestamp 1
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_727
timestamp 1
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_729
timestamp 1636968456
transform 1 0 68172 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_741
timestamp 1636968456
transform 1 0 69276 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_753
timestamp 1636968456
transform 1 0 70380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_765
timestamp 1636968456
transform 1 0 71484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_777
timestamp 1
transform 1 0 72588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_783
timestamp 1
transform 1 0 73140 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_785
timestamp 1636968456
transform 1 0 73324 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_797
timestamp 1636968456
transform 1 0 74428 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_809
timestamp 1636968456
transform 1 0 75532 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_821
timestamp 1636968456
transform 1 0 76636 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_833
timestamp 1
transform 1 0 77740 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_839
timestamp 1
transform 1 0 78292 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_841
timestamp 1
transform 1 0 78476 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_3
timestamp 1
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_11
timestamp 1636968456
transform 1 0 2116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_23
timestamp 1
transform 1 0 3220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1636968456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1636968456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1636968456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1636968456
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_85
timestamp 1
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_93
timestamp 1
transform 1 0 9660 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_124
timestamp 1636968456
transform 1 0 12512 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_136
timestamp 1
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1636968456
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1636968456
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1636968456
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1636968456
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_197
timestamp 1
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_203
timestamp 1
transform 1 0 19780 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_210
timestamp 1
transform 1 0 20424 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_218
timestamp 1
transform 1 0 21160 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_228
timestamp 1636968456
transform 1 0 22080 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_240
timestamp 1636968456
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1636968456
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1636968456
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1636968456
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1636968456
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_309
timestamp 1
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_317
timestamp 1
transform 1 0 30268 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_327
timestamp 1
transform 1 0 31188 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_335
timestamp 1
transform 1 0 31924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_344
timestamp 1636968456
transform 1 0 32752 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_356
timestamp 1
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_374
timestamp 1636968456
transform 1 0 35512 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_386
timestamp 1636968456
transform 1 0 36616 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_398
timestamp 1636968456
transform 1 0 37720 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_410
timestamp 1
transform 1 0 38824 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_418
timestamp 1
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_421
timestamp 1
transform 1 0 39836 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_438
timestamp 1636968456
transform 1 0 41400 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_450
timestamp 1636968456
transform 1 0 42504 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_462
timestamp 1
transform 1 0 43608 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_466
timestamp 1
transform 1 0 43976 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_472
timestamp 1
transform 1 0 44528 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_494
timestamp 1
transform 1 0 46552 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_519
timestamp 1
transform 1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_529
timestamp 1
transform 1 0 49772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_548
timestamp 1
transform 1 0 51520 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_560
timestamp 1
transform 1 0 52624 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_576
timestamp 1636968456
transform 1 0 54096 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_589
timestamp 1636968456
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_601
timestamp 1636968456
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_613
timestamp 1636968456
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_625
timestamp 1636968456
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_637
timestamp 1
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_643
timestamp 1
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_645
timestamp 1636968456
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_657
timestamp 1636968456
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_669
timestamp 1636968456
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_681
timestamp 1636968456
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_693
timestamp 1
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_699
timestamp 1
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_701
timestamp 1636968456
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_713
timestamp 1636968456
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_725
timestamp 1636968456
transform 1 0 67804 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_737
timestamp 1636968456
transform 1 0 68908 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_749
timestamp 1
transform 1 0 70012 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_755
timestamp 1
transform 1 0 70564 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_757
timestamp 1636968456
transform 1 0 70748 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_769
timestamp 1636968456
transform 1 0 71852 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_781
timestamp 1636968456
transform 1 0 72956 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_793
timestamp 1636968456
transform 1 0 74060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_805
timestamp 1
transform 1 0 75164 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_811
timestamp 1
transform 1 0 75716 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_813
timestamp 1636968456
transform 1 0 75900 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_825
timestamp 1636968456
transform 1 0 77004 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_837
timestamp 1
transform 1 0 78108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_841
timestamp 1
transform 1 0 78476 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_3
timestamp 1
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_7
timestamp 1
transform 1 0 1748 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_11
timestamp 1636968456
transform 1 0 2116 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_23
timestamp 1636968456
transform 1 0 3220 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_35
timestamp 1636968456
transform 1 0 4324 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_47
timestamp 1
transform 1 0 5428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1636968456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1636968456
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1636968456
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_93
timestamp 1
transform 1 0 9660 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_97
timestamp 1
transform 1 0 10028 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_106
timestamp 1
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_120
timestamp 1
transform 1 0 12144 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1636968456
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1636968456
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_181
timestamp 1
transform 1 0 17756 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_206
timestamp 1
transform 1 0 20056 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_213
timestamp 1
transform 1 0 20700 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_221
timestamp 1
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1636968456
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1636968456
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1636968456
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1636968456
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1636968456
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1636968456
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1636968456
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1636968456
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_329
timestamp 1
transform 1 0 31372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_333
timestamp 1
transform 1 0 31740 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_358
timestamp 1
transform 1 0 34040 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_366
timestamp 1
transform 1 0 34776 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_378
timestamp 1
transform 1 0 35880 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_390
timestamp 1
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_393
timestamp 1
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_401
timestamp 1
transform 1 0 37996 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_409
timestamp 1
transform 1 0 38732 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_417
timestamp 1
transform 1 0 39468 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_442
timestamp 1
transform 1 0 41768 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_453
timestamp 1
transform 1 0 42780 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_457
timestamp 1
transform 1 0 43148 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_478
timestamp 1
transform 1 0 45080 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_486
timestamp 1
transform 1 0 45816 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_490
timestamp 1636968456
transform 1 0 46184 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_502
timestamp 1
transform 1 0 47288 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_505
timestamp 1
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_513
timestamp 1
transform 1 0 48300 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_555
timestamp 1
transform 1 0 52164 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_559
timestamp 1
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_581
timestamp 1636968456
transform 1 0 54556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_593
timestamp 1636968456
transform 1 0 55660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_605
timestamp 1
transform 1 0 56764 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_613
timestamp 1
transform 1 0 57500 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_617
timestamp 1636968456
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_629
timestamp 1636968456
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_641
timestamp 1636968456
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_653
timestamp 1636968456
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_665
timestamp 1
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_671
timestamp 1
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_673
timestamp 1636968456
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_685
timestamp 1636968456
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_697
timestamp 1636968456
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_709
timestamp 1636968456
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_721
timestamp 1
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_727
timestamp 1
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_729
timestamp 1636968456
transform 1 0 68172 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_741
timestamp 1636968456
transform 1 0 69276 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_753
timestamp 1636968456
transform 1 0 70380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_765
timestamp 1636968456
transform 1 0 71484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_777
timestamp 1
transform 1 0 72588 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_783
timestamp 1
transform 1 0 73140 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_785
timestamp 1636968456
transform 1 0 73324 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_797
timestamp 1636968456
transform 1 0 74428 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_809
timestamp 1636968456
transform 1 0 75532 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_821
timestamp 1636968456
transform 1 0 76636 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_833
timestamp 1
transform 1 0 77740 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_839
timestamp 1
transform 1 0 78292 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_841
timestamp 1
transform 1 0 78476 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_3
timestamp 1
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_14
timestamp 1636968456
transform 1 0 2392 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_26
timestamp 1
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1636968456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1636968456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1636968456
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1636968456
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_97
timestamp 1
transform 1 0 10028 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_110
timestamp 1636968456
transform 1 0 11224 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_129
timestamp 1
transform 1 0 12972 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_149
timestamp 1
transform 1 0 14812 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_157
timestamp 1
transform 1 0 15548 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_182
timestamp 1636968456
transform 1 0 17848 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_194
timestamp 1
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_235
timestamp 1636968456
transform 1 0 22724 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_247
timestamp 1
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1636968456
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1636968456
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1636968456
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1636968456
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1636968456
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1636968456
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1636968456
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_345
timestamp 1
transform 1 0 32844 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_353
timestamp 1
transform 1 0 33580 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_365
timestamp 1
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_369
timestamp 1
transform 1 0 35052 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_377
timestamp 1
transform 1 0 35788 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_383
timestamp 1
transform 1 0 36340 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_393
timestamp 1
transform 1 0 37260 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 1636968456
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_433
timestamp 1636968456
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_445
timestamp 1
transform 1 0 42044 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_449
timestamp 1
transform 1 0 42412 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_467
timestamp 1
transform 1 0 44068 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_475
timestamp 1
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_477
timestamp 1
transform 1 0 44988 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_485
timestamp 1
transform 1 0 45724 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_489
timestamp 1636968456
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_501
timestamp 1636968456
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_513
timestamp 1636968456
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_525
timestamp 1
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_531
timestamp 1
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_533
timestamp 1636968456
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_545
timestamp 1636968456
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_557
timestamp 1636968456
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_569
timestamp 1636968456
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_581
timestamp 1
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_587
timestamp 1
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_589
timestamp 1636968456
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_601
timestamp 1636968456
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_613
timestamp 1636968456
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_625
timestamp 1636968456
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_637
timestamp 1
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_643
timestamp 1
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_645
timestamp 1636968456
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_657
timestamp 1636968456
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_669
timestamp 1636968456
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_681
timestamp 1636968456
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_693
timestamp 1
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_699
timestamp 1
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_701
timestamp 1636968456
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_713
timestamp 1636968456
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_725
timestamp 1636968456
transform 1 0 67804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_737
timestamp 1636968456
transform 1 0 68908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_749
timestamp 1
transform 1 0 70012 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_755
timestamp 1
transform 1 0 70564 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_757
timestamp 1636968456
transform 1 0 70748 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_769
timestamp 1636968456
transform 1 0 71852 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_781
timestamp 1636968456
transform 1 0 72956 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_793
timestamp 1636968456
transform 1 0 74060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_805
timestamp 1
transform 1 0 75164 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_811
timestamp 1
transform 1 0 75716 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_813
timestamp 1636968456
transform 1 0 75900 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_825
timestamp 1636968456
transform 1 0 77004 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_837
timestamp 1
transform 1 0 78108 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_841
timestamp 1
transform 1 0 78476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_3
timestamp 1
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_14
timestamp 1636968456
transform 1 0 2392 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_26
timestamp 1636968456
transform 1 0 3496 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_38
timestamp 1636968456
transform 1 0 4600 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_50
timestamp 1
transform 1 0 5704 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_69
timestamp 1
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_77
timestamp 1
transform 1 0 8188 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_110
timestamp 1
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1636968456
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_125
timestamp 1
transform 1 0 12604 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_129
timestamp 1
transform 1 0 12972 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_152
timestamp 1
transform 1 0 15088 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_164
timestamp 1
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_191
timestamp 1636968456
transform 1 0 18676 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_203
timestamp 1
transform 1 0 19780 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_220
timestamp 1
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1636968456
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1636968456
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1636968456
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1636968456
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1636968456
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1636968456
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1636968456
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1636968456
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_337
timestamp 1
transform 1 0 32108 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_387
timestamp 1
transform 1 0 36708 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1636968456
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_405
timestamp 1636968456
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_417
timestamp 1636968456
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_429
timestamp 1
transform 1 0 40572 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_445
timestamp 1
transform 1 0 42044 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_449
timestamp 1
transform 1 0 42412 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_461
timestamp 1
transform 1 0 43516 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_472
timestamp 1
transform 1 0 44528 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_493
timestamp 1
transform 1 0 46460 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_501
timestamp 1
transform 1 0 47196 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_514
timestamp 1636968456
transform 1 0 48392 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_526
timestamp 1636968456
transform 1 0 49496 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_538
timestamp 1636968456
transform 1 0 50600 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_550
timestamp 1
transform 1 0 51704 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_558
timestamp 1
transform 1 0 52440 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_561
timestamp 1636968456
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_573
timestamp 1636968456
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_585
timestamp 1636968456
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_597
timestamp 1636968456
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_609
timestamp 1
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_615
timestamp 1
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_617
timestamp 1636968456
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_629
timestamp 1636968456
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_641
timestamp 1636968456
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_653
timestamp 1636968456
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_665
timestamp 1
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_671
timestamp 1
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_673
timestamp 1636968456
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_685
timestamp 1636968456
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_697
timestamp 1636968456
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_709
timestamp 1636968456
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_721
timestamp 1
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_727
timestamp 1
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_729
timestamp 1636968456
transform 1 0 68172 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_741
timestamp 1636968456
transform 1 0 69276 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_753
timestamp 1636968456
transform 1 0 70380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_765
timestamp 1636968456
transform 1 0 71484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_777
timestamp 1
transform 1 0 72588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_783
timestamp 1
transform 1 0 73140 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_785
timestamp 1636968456
transform 1 0 73324 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_797
timestamp 1636968456
transform 1 0 74428 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_809
timestamp 1636968456
transform 1 0 75532 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_821
timestamp 1636968456
transform 1 0 76636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_833
timestamp 1
transform 1 0 77740 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_839
timestamp 1
transform 1 0 78292 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_841
timestamp 1
transform 1 0 78476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_3
timestamp 1
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_11
timestamp 1636968456
transform 1 0 2116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_23
timestamp 1
transform 1 0 3220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1636968456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1636968456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1636968456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1636968456
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_85
timestamp 1
transform 1 0 8924 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_99
timestamp 1
transform 1 0 10212 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_103
timestamp 1
transform 1 0 10580 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_116
timestamp 1
transform 1 0 11776 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_137
timestamp 1
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_141
timestamp 1
transform 1 0 14076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_149
timestamp 1
transform 1 0 14812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_168
timestamp 1
transform 1 0 16560 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_178
timestamp 1636968456
transform 1 0 17480 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_190
timestamp 1
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_197
timestamp 1
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_205
timestamp 1
transform 1 0 19964 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_211
timestamp 1
transform 1 0 20516 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_217
timestamp 1636968456
transform 1 0 21068 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_229
timestamp 1636968456
transform 1 0 22172 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_241
timestamp 1
transform 1 0 23276 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_249
timestamp 1
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1636968456
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1636968456
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1636968456
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1636968456
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1636968456
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1636968456
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 1636968456
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 1636968456
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1636968456
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_377
timestamp 1
transform 1 0 35788 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_414
timestamp 1
transform 1 0 39192 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_444
timestamp 1
transform 1 0 41952 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_448
timestamp 1
transform 1 0 42320 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_461
timestamp 1636968456
transform 1 0 43516 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_473
timestamp 1
transform 1 0 44620 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_477
timestamp 1
transform 1 0 44988 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_485
timestamp 1
transform 1 0 45724 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_496
timestamp 1
transform 1 0 46736 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_529
timestamp 1
transform 1 0 49772 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_533
timestamp 1636968456
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_545
timestamp 1636968456
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_557
timestamp 1636968456
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_569
timestamp 1636968456
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_581
timestamp 1
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_587
timestamp 1
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_589
timestamp 1636968456
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_601
timestamp 1636968456
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_613
timestamp 1636968456
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_625
timestamp 1636968456
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_637
timestamp 1
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_643
timestamp 1
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_645
timestamp 1636968456
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_657
timestamp 1636968456
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_669
timestamp 1636968456
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_681
timestamp 1636968456
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_693
timestamp 1
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_699
timestamp 1
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_701
timestamp 1636968456
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_713
timestamp 1636968456
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_725
timestamp 1636968456
transform 1 0 67804 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_737
timestamp 1636968456
transform 1 0 68908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_749
timestamp 1
transform 1 0 70012 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_755
timestamp 1
transform 1 0 70564 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_757
timestamp 1636968456
transform 1 0 70748 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_769
timestamp 1636968456
transform 1 0 71852 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_781
timestamp 1636968456
transform 1 0 72956 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_793
timestamp 1636968456
transform 1 0 74060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_805
timestamp 1
transform 1 0 75164 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_811
timestamp 1
transform 1 0 75716 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_813
timestamp 1636968456
transform 1 0 75900 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_825
timestamp 1636968456
transform 1 0 77004 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_837
timestamp 1
transform 1 0 78108 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_841
timestamp 1
transform 1 0 78476 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_3
timestamp 1
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_14
timestamp 1636968456
transform 1 0 2392 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_26
timestamp 1636968456
transform 1 0 3496 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_38
timestamp 1636968456
transform 1 0 4600 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_50
timestamp 1
transform 1 0 5704 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1636968456
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1636968456
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1636968456
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_93
timestamp 1
transform 1 0 9660 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_101
timestamp 1
transform 1 0 10396 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_110
timestamp 1
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_121
timestamp 1
transform 1 0 12236 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_127
timestamp 1
transform 1 0 12788 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_150
timestamp 1
transform 1 0 14904 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_154
timestamp 1
transform 1 0 15272 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_158
timestamp 1
transform 1 0 15640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_166
timestamp 1
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_172
timestamp 1636968456
transform 1 0 16928 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_184
timestamp 1
transform 1 0 18032 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_192
timestamp 1
transform 1 0 18768 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_216
timestamp 1
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_233
timestamp 1636968456
transform 1 0 22540 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_245
timestamp 1636968456
transform 1 0 23644 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_257
timestamp 1636968456
transform 1 0 24748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_269
timestamp 1
transform 1 0 25852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_277
timestamp 1
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1636968456
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1636968456
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_305
timestamp 1
transform 1 0 29164 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_313
timestamp 1
transform 1 0 29900 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1636968456
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_357
timestamp 1636968456
transform 1 0 33948 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_369
timestamp 1636968456
transform 1 0 35052 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_381
timestamp 1
transform 1 0 36156 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_389
timestamp 1
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_393
timestamp 1
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_425
timestamp 1
transform 1 0 40204 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_439
timestamp 1
transform 1 0 41492 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_447
timestamp 1
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_449
timestamp 1
transform 1 0 42412 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_462
timestamp 1
transform 1 0 43608 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_472
timestamp 1
transform 1 0 44528 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_480
timestamp 1
transform 1 0 45264 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_494
timestamp 1
transform 1 0 46552 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_502
timestamp 1
transform 1 0 47288 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_505
timestamp 1
transform 1 0 47564 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_511
timestamp 1
transform 1 0 48116 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_518
timestamp 1636968456
transform 1 0 48760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_530
timestamp 1636968456
transform 1 0 49864 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_542
timestamp 1636968456
transform 1 0 50968 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_554
timestamp 1
transform 1 0 52072 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_561
timestamp 1636968456
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_573
timestamp 1636968456
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_585
timestamp 1636968456
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_597
timestamp 1636968456
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_609
timestamp 1
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_615
timestamp 1
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_617
timestamp 1636968456
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_629
timestamp 1636968456
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_641
timestamp 1636968456
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_653
timestamp 1636968456
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_665
timestamp 1
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_671
timestamp 1
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_673
timestamp 1636968456
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_685
timestamp 1636968456
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_697
timestamp 1636968456
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_709
timestamp 1636968456
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_721
timestamp 1
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_727
timestamp 1
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_729
timestamp 1636968456
transform 1 0 68172 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_741
timestamp 1636968456
transform 1 0 69276 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_753
timestamp 1636968456
transform 1 0 70380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_765
timestamp 1636968456
transform 1 0 71484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_777
timestamp 1
transform 1 0 72588 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_783
timestamp 1
transform 1 0 73140 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_785
timestamp 1636968456
transform 1 0 73324 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_797
timestamp 1636968456
transform 1 0 74428 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_809
timestamp 1636968456
transform 1 0 75532 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_821
timestamp 1636968456
transform 1 0 76636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_833
timestamp 1
transform 1 0 77740 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_839
timestamp 1
transform 1 0 78292 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_841
timestamp 1
transform 1 0 78476 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_3
timestamp 1
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_7
timestamp 1
transform 1 0 1748 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_11
timestamp 1636968456
transform 1 0 2116 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_23
timestamp 1
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1636968456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1636968456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1636968456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1636968456
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_115
timestamp 1636968456
transform 1 0 11684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_127
timestamp 1636968456
transform 1 0 12788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_141
timestamp 1
transform 1 0 14076 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_149
timestamp 1
transform 1 0 14812 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_158
timestamp 1
transform 1 0 15640 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1636968456
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_177
timestamp 1
transform 1 0 17388 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_200
timestamp 1
transform 1 0 19504 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_231
timestamp 1636968456
transform 1 0 22356 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_243
timestamp 1
transform 1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1636968456
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1636968456
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1636968456
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1636968456
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_329
timestamp 1
transform 1 0 31372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_333
timestamp 1
transform 1 0 31740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_342
timestamp 1636968456
transform 1 0 32568 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_354
timestamp 1
transform 1 0 33672 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_362
timestamp 1
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_371
timestamp 1
transform 1 0 35236 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_412
timestamp 1
transform 1 0 39008 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_421
timestamp 1636968456
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_433
timestamp 1636968456
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_445
timestamp 1
transform 1 0 42044 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_470
timestamp 1
transform 1 0 44344 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_477
timestamp 1636968456
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_489
timestamp 1636968456
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_501
timestamp 1636968456
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_513
timestamp 1636968456
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_525
timestamp 1
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_531
timestamp 1
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_533
timestamp 1636968456
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_545
timestamp 1636968456
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_557
timestamp 1636968456
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_569
timestamp 1636968456
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_581
timestamp 1
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_587
timestamp 1
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_589
timestamp 1636968456
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_601
timestamp 1636968456
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_613
timestamp 1636968456
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_625
timestamp 1636968456
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_637
timestamp 1
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_643
timestamp 1
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_645
timestamp 1636968456
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_657
timestamp 1636968456
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_669
timestamp 1636968456
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_681
timestamp 1636968456
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_693
timestamp 1
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_699
timestamp 1
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_701
timestamp 1636968456
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_713
timestamp 1636968456
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_725
timestamp 1636968456
transform 1 0 67804 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_737
timestamp 1636968456
transform 1 0 68908 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_749
timestamp 1
transform 1 0 70012 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_755
timestamp 1
transform 1 0 70564 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_757
timestamp 1636968456
transform 1 0 70748 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_769
timestamp 1636968456
transform 1 0 71852 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_781
timestamp 1636968456
transform 1 0 72956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_793
timestamp 1636968456
transform 1 0 74060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_805
timestamp 1
transform 1 0 75164 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_811
timestamp 1
transform 1 0 75716 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_813
timestamp 1636968456
transform 1 0 75900 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_825
timestamp 1636968456
transform 1 0 77004 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_837
timestamp 1
transform 1 0 78108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_841
timestamp 1
transform 1 0 78476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_3
timestamp 1
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_14
timestamp 1636968456
transform 1 0 2392 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_26
timestamp 1636968456
transform 1 0 3496 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_38
timestamp 1636968456
transform 1 0 4600 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_50
timestamp 1
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1636968456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1636968456
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1636968456
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1636968456
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_113
timestamp 1
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_119
timestamp 1
transform 1 0 12052 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_136
timestamp 1
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_148
timestamp 1
transform 1 0 14720 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_156
timestamp 1
transform 1 0 15456 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_164
timestamp 1
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_169
timestamp 1
transform 1 0 16652 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_182
timestamp 1
transform 1 0 17848 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_191
timestamp 1
transform 1 0 18676 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_200
timestamp 1636968456
transform 1 0 19504 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_212
timestamp 1636968456
transform 1 0 20608 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1636968456
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1636968456
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1636968456
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1636968456
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1636968456
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1636968456
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_305
timestamp 1
transform 1 0 29164 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_340
timestamp 1
transform 1 0 32384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_349
timestamp 1
transform 1 0 33212 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_357
timestamp 1
transform 1 0 33948 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_388
timestamp 1
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_401
timestamp 1636968456
transform 1 0 37996 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_413
timestamp 1
transform 1 0 39100 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_434
timestamp 1636968456
transform 1 0 41032 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_446
timestamp 1
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_477
timestamp 1636968456
transform 1 0 44988 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_489
timestamp 1
transform 1 0 46092 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_499
timestamp 1
transform 1 0 47012 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_503
timestamp 1
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_505
timestamp 1636968456
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_517
timestamp 1636968456
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_529
timestamp 1636968456
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_541
timestamp 1636968456
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_553
timestamp 1
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_559
timestamp 1
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_561
timestamp 1636968456
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_573
timestamp 1636968456
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_585
timestamp 1636968456
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_597
timestamp 1636968456
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_609
timestamp 1
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_615
timestamp 1
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_617
timestamp 1636968456
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_629
timestamp 1636968456
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_641
timestamp 1636968456
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_653
timestamp 1636968456
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_665
timestamp 1
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_671
timestamp 1
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_673
timestamp 1636968456
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_685
timestamp 1636968456
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_697
timestamp 1636968456
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_709
timestamp 1636968456
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_721
timestamp 1
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_727
timestamp 1
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_729
timestamp 1636968456
transform 1 0 68172 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_741
timestamp 1636968456
transform 1 0 69276 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_753
timestamp 1636968456
transform 1 0 70380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_765
timestamp 1636968456
transform 1 0 71484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_777
timestamp 1
transform 1 0 72588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_783
timestamp 1
transform 1 0 73140 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_785
timestamp 1636968456
transform 1 0 73324 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_797
timestamp 1636968456
transform 1 0 74428 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_809
timestamp 1636968456
transform 1 0 75532 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_821
timestamp 1636968456
transform 1 0 76636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_833
timestamp 1
transform 1 0 77740 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_839
timestamp 1
transform 1 0 78292 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_841
timestamp 1
transform 1 0 78476 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_3
timestamp 1
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_14
timestamp 1636968456
transform 1 0 2392 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 1
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1636968456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1636968456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1636968456
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1636968456
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1636968456
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_97
timestamp 1
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_105
timestamp 1
transform 1 0 10764 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_113
timestamp 1
transform 1 0 11500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1636968456
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1636968456
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_157
timestamp 1636968456
transform 1 0 15548 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_169
timestamp 1
transform 1 0 16652 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_173
timestamp 1
transform 1 0 17020 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_178
timestamp 1
transform 1 0 17480 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_190
timestamp 1
transform 1 0 18584 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1636968456
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1636968456
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1636968456
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1636968456
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1636968456
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1636968456
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_277
timestamp 1
transform 1 0 26588 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_305
timestamp 1
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1636968456
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_323
timestamp 1
transform 1 0 30820 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_338
timestamp 1
transform 1 0 32200 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_361
timestamp 1
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1636968456
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_377
timestamp 1
transform 1 0 35788 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_385
timestamp 1
transform 1 0 36524 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_403
timestamp 1636968456
transform 1 0 38180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_415
timestamp 1
transform 1 0 39284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_419
timestamp 1
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_421
timestamp 1
transform 1 0 39836 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_432
timestamp 1
transform 1 0 40848 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_460
timestamp 1
transform 1 0 43424 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_465
timestamp 1
transform 1 0 43884 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_473
timestamp 1
transform 1 0 44620 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_497
timestamp 1
transform 1 0 46828 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_520
timestamp 1636968456
transform 1 0 48944 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_533
timestamp 1636968456
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_545
timestamp 1636968456
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_557
timestamp 1636968456
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_569
timestamp 1636968456
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_581
timestamp 1
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_587
timestamp 1
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_589
timestamp 1636968456
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_601
timestamp 1636968456
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_613
timestamp 1636968456
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_625
timestamp 1636968456
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_637
timestamp 1
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_643
timestamp 1
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_645
timestamp 1636968456
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_657
timestamp 1636968456
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_669
timestamp 1636968456
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_681
timestamp 1636968456
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_693
timestamp 1
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_699
timestamp 1
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_701
timestamp 1636968456
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_713
timestamp 1636968456
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_725
timestamp 1636968456
transform 1 0 67804 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_737
timestamp 1636968456
transform 1 0 68908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_749
timestamp 1
transform 1 0 70012 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_755
timestamp 1
transform 1 0 70564 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_757
timestamp 1636968456
transform 1 0 70748 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_769
timestamp 1636968456
transform 1 0 71852 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_781
timestamp 1636968456
transform 1 0 72956 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_793
timestamp 1636968456
transform 1 0 74060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_805
timestamp 1
transform 1 0 75164 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_811
timestamp 1
transform 1 0 75716 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_813
timestamp 1636968456
transform 1 0 75900 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_825
timestamp 1636968456
transform 1 0 77004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_837
timestamp 1
transform 1 0 78108 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_841
timestamp 1
transform 1 0 78476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_3
timestamp 1
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_11
timestamp 1636968456
transform 1 0 2116 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_23
timestamp 1636968456
transform 1 0 3220 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_35
timestamp 1636968456
transform 1 0 4324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_47
timestamp 1
transform 1 0 5428 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1636968456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1636968456
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_81
timestamp 1
transform 1 0 8556 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_89
timestamp 1
transform 1 0 9292 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_123
timestamp 1
transform 1 0 12420 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_143
timestamp 1
transform 1 0 14260 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_147
timestamp 1
transform 1 0 14628 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_179
timestamp 1
transform 1 0 17572 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_210
timestamp 1636968456
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_222
timestamp 1
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1636968456
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1636968456
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1636968456
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1636968456
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_281
timestamp 1
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_285
timestamp 1
transform 1 0 27324 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_293
timestamp 1
transform 1 0 28060 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_297
timestamp 1
transform 1 0 28428 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_306
timestamp 1
transform 1 0 29256 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_315
timestamp 1
transform 1 0 30084 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_331
timestamp 1
transform 1 0 31556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1636968456
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1636968456
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 1636968456
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 1636968456
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_385
timestamp 1
transform 1 0 36524 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_413
timestamp 1
transform 1 0 39100 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_419
timestamp 1
transform 1 0 39652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_436
timestamp 1
transform 1 0 41216 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_442
timestamp 1
transform 1 0 41768 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_457
timestamp 1636968456
transform 1 0 43148 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_469
timestamp 1
transform 1 0 44252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_473
timestamp 1
transform 1 0 44620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_491
timestamp 1
transform 1 0 46276 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_501
timestamp 1
transform 1 0 47196 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_505
timestamp 1636968456
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_517
timestamp 1636968456
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_529
timestamp 1636968456
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_541
timestamp 1636968456
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_553
timestamp 1
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_559
timestamp 1
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_561
timestamp 1636968456
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_573
timestamp 1636968456
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_585
timestamp 1636968456
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_597
timestamp 1636968456
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_609
timestamp 1
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_615
timestamp 1
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_617
timestamp 1636968456
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_629
timestamp 1636968456
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_641
timestamp 1636968456
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_653
timestamp 1636968456
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_665
timestamp 1
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_671
timestamp 1
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_673
timestamp 1636968456
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_685
timestamp 1636968456
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_697
timestamp 1636968456
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_709
timestamp 1636968456
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_721
timestamp 1
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_727
timestamp 1
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_729
timestamp 1636968456
transform 1 0 68172 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_741
timestamp 1636968456
transform 1 0 69276 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_753
timestamp 1636968456
transform 1 0 70380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_765
timestamp 1636968456
transform 1 0 71484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_777
timestamp 1
transform 1 0 72588 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_783
timestamp 1
transform 1 0 73140 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_785
timestamp 1636968456
transform 1 0 73324 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_797
timestamp 1636968456
transform 1 0 74428 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_809
timestamp 1636968456
transform 1 0 75532 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_821
timestamp 1636968456
transform 1 0 76636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_833
timestamp 1
transform 1 0 77740 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_839
timestamp 1
transform 1 0 78292 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_841
timestamp 1
transform 1 0 78476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_3
timestamp 1
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_14
timestamp 1636968456
transform 1 0 2392 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_26
timestamp 1
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1636968456
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1636968456
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1636968456
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1636968456
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1636968456
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1636968456
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_109
timestamp 1
transform 1 0 11132 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_117
timestamp 1
transform 1 0 11868 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_143
timestamp 1636968456
transform 1 0 14260 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_158
timestamp 1
transform 1 0 15640 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_166
timestamp 1
transform 1 0 16376 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_175
timestamp 1
transform 1 0 17204 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_181
timestamp 1
transform 1 0 17756 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_190
timestamp 1
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1636968456
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_209
timestamp 1
transform 1 0 20332 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_225
timestamp 1636968456
transform 1 0 21804 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_237
timestamp 1636968456
transform 1 0 22908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_249
timestamp 1
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1636968456
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1636968456
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1636968456
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_289
timestamp 1
transform 1 0 27692 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_293
timestamp 1636968456
transform 1 0 28060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_305
timestamp 1
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1636968456
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1636968456
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 1
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_371
timestamp 1636968456
transform 1 0 35236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_383
timestamp 1
transform 1 0 36340 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_391
timestamp 1
transform 1 0 37076 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_397
timestamp 1636968456
transform 1 0 37628 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_409
timestamp 1
transform 1 0 38732 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_417
timestamp 1
transform 1 0 39468 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 1636968456
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_433
timestamp 1636968456
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_445
timestamp 1636968456
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_457
timestamp 1
transform 1 0 43148 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_472
timestamp 1
transform 1 0 44528 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_477
timestamp 1636968456
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_494
timestamp 1636968456
transform 1 0 46552 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_506
timestamp 1636968456
transform 1 0 47656 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_518
timestamp 1636968456
transform 1 0 48760 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_530
timestamp 1
transform 1 0 49864 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_533
timestamp 1636968456
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_545
timestamp 1636968456
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_557
timestamp 1636968456
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_569
timestamp 1636968456
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_581
timestamp 1
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_587
timestamp 1
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_589
timestamp 1636968456
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_601
timestamp 1636968456
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_613
timestamp 1636968456
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_625
timestamp 1636968456
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_637
timestamp 1
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_643
timestamp 1
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_645
timestamp 1636968456
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_657
timestamp 1636968456
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_669
timestamp 1636968456
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_681
timestamp 1636968456
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_693
timestamp 1
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_699
timestamp 1
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_701
timestamp 1636968456
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_713
timestamp 1636968456
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_725
timestamp 1636968456
transform 1 0 67804 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_737
timestamp 1636968456
transform 1 0 68908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_749
timestamp 1
transform 1 0 70012 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_755
timestamp 1
transform 1 0 70564 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_757
timestamp 1636968456
transform 1 0 70748 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_769
timestamp 1636968456
transform 1 0 71852 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_781
timestamp 1636968456
transform 1 0 72956 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_793
timestamp 1636968456
transform 1 0 74060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_805
timestamp 1
transform 1 0 75164 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_811
timestamp 1
transform 1 0 75716 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_813
timestamp 1636968456
transform 1 0 75900 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_825
timestamp 1636968456
transform 1 0 77004 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_837
timestamp 1
transform 1 0 78108 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_841
timestamp 1
transform 1 0 78476 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_3
timestamp 1
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_7
timestamp 1
transform 1 0 1748 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_11
timestamp 1636968456
transform 1 0 2116 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_23
timestamp 1636968456
transform 1 0 3220 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_35
timestamp 1636968456
transform 1 0 4324 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_47
timestamp 1
transform 1 0 5428 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1636968456
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1636968456
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1636968456
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1636968456
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1636968456
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1636968456
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1636968456
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1636968456
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_169
timestamp 1
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_173
timestamp 1
transform 1 0 17020 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_196
timestamp 1636968456
transform 1 0 19136 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_208
timestamp 1636968456
transform 1 0 20240 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_220
timestamp 1
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1636968456
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1636968456
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1636968456
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1636968456
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_306
timestamp 1
transform 1 0 29256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_337
timestamp 1
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_389
timestamp 1
transform 1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1636968456
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1636968456
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 1636968456
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_429
timestamp 1636968456
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_441
timestamp 1
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_447
timestamp 1
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_449
timestamp 1
transform 1 0 42412 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_457
timestamp 1
transform 1 0 43148 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_477
timestamp 1
transform 1 0 44988 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_484
timestamp 1
transform 1 0 45632 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_491
timestamp 1636968456
transform 1 0 46276 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_503
timestamp 1
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_514
timestamp 1636968456
transform 1 0 48392 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_526
timestamp 1636968456
transform 1 0 49496 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_538
timestamp 1636968456
transform 1 0 50600 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_550
timestamp 1
transform 1 0 51704 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_558
timestamp 1
transform 1 0 52440 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_561
timestamp 1636968456
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_573
timestamp 1636968456
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_585
timestamp 1636968456
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_597
timestamp 1636968456
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_609
timestamp 1
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_615
timestamp 1
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_617
timestamp 1636968456
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_629
timestamp 1636968456
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_641
timestamp 1636968456
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_653
timestamp 1636968456
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_665
timestamp 1
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_671
timestamp 1
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_673
timestamp 1636968456
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_685
timestamp 1636968456
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_697
timestamp 1636968456
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_709
timestamp 1636968456
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_721
timestamp 1
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_727
timestamp 1
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_729
timestamp 1636968456
transform 1 0 68172 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_741
timestamp 1636968456
transform 1 0 69276 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_753
timestamp 1636968456
transform 1 0 70380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_765
timestamp 1636968456
transform 1 0 71484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_777
timestamp 1
transform 1 0 72588 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_783
timestamp 1
transform 1 0 73140 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_785
timestamp 1636968456
transform 1 0 73324 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_797
timestamp 1636968456
transform 1 0 74428 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_809
timestamp 1636968456
transform 1 0 75532 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_821
timestamp 1636968456
transform 1 0 76636 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_833
timestamp 1
transform 1 0 77740 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_839
timestamp 1
transform 1 0 78292 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_841
timestamp 1
transform 1 0 78476 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_3
timestamp 1
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_14
timestamp 1636968456
transform 1 0 2392 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_26
timestamp 1
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1636968456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1636968456
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1636968456
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1636968456
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1636968456
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1636968456
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1636968456
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1636968456
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1636968456
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1636968456
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1636968456
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1636968456
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1636968456
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1636968456
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1636968456
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1636968456
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1636968456
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1636968456
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1636968456
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_289
timestamp 1
transform 1 0 27692 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_298
timestamp 1
transform 1 0 28520 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_320
timestamp 1636968456
transform 1 0 30544 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_332
timestamp 1
transform 1 0 31648 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_341
timestamp 1
transform 1 0 32476 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_345
timestamp 1
transform 1 0 32844 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_361
timestamp 1
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_365
timestamp 1
transform 1 0 34684 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_378
timestamp 1636968456
transform 1 0 35880 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_423
timestamp 1
transform 1 0 40020 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_431
timestamp 1
transform 1 0 40756 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_452
timestamp 1
transform 1 0 42688 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_460
timestamp 1
transform 1 0 43424 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_474
timestamp 1
transform 1 0 44712 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_497
timestamp 1
transform 1 0 46828 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_533
timestamp 1636968456
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_545
timestamp 1636968456
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_557
timestamp 1636968456
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_569
timestamp 1636968456
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_581
timestamp 1
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_587
timestamp 1
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_589
timestamp 1636968456
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_601
timestamp 1636968456
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_613
timestamp 1636968456
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_625
timestamp 1636968456
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_637
timestamp 1
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_643
timestamp 1
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_645
timestamp 1636968456
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_657
timestamp 1636968456
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_669
timestamp 1636968456
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_681
timestamp 1636968456
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_693
timestamp 1
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_699
timestamp 1
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_701
timestamp 1636968456
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_713
timestamp 1636968456
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_725
timestamp 1636968456
transform 1 0 67804 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_737
timestamp 1636968456
transform 1 0 68908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_749
timestamp 1
transform 1 0 70012 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_755
timestamp 1
transform 1 0 70564 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_757
timestamp 1636968456
transform 1 0 70748 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_769
timestamp 1636968456
transform 1 0 71852 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_781
timestamp 1636968456
transform 1 0 72956 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_793
timestamp 1636968456
transform 1 0 74060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_805
timestamp 1
transform 1 0 75164 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_811
timestamp 1
transform 1 0 75716 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_813
timestamp 1636968456
transform 1 0 75900 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_825
timestamp 1636968456
transform 1 0 77004 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_837
timestamp 1
transform 1 0 78108 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_841
timestamp 1
transform 1 0 78476 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_3
timestamp 1
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_14
timestamp 1636968456
transform 1 0 2392 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_26
timestamp 1636968456
transform 1 0 3496 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_38
timestamp 1636968456
transform 1 0 4600 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_50
timestamp 1
transform 1 0 5704 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1636968456
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1636968456
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1636968456
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1636968456
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1636968456
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1636968456
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1636968456
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1636968456
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1636968456
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1636968456
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1636968456
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1636968456
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1636968456
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1636968456
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1636968456
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1636968456
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1636968456
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_293
timestamp 1
transform 1 0 28060 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_298
timestamp 1
transform 1 0 28520 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_314
timestamp 1
transform 1 0 29992 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_324
timestamp 1636968456
transform 1 0 30912 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_345
timestamp 1636968456
transform 1 0 32844 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_357
timestamp 1636968456
transform 1 0 33948 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_369
timestamp 1
transform 1 0 35052 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_376
timestamp 1
transform 1 0 35696 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_382
timestamp 1
transform 1 0 36248 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_386
timestamp 1
transform 1 0 36616 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_393
timestamp 1
transform 1 0 37260 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_399
timestamp 1
transform 1 0 37812 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_408
timestamp 1
transform 1 0 38640 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_424
timestamp 1
transform 1 0 40112 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_438
timestamp 1
transform 1 0 41400 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_447
timestamp 1
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_455
timestamp 1636968456
transform 1 0 42964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_467
timestamp 1
transform 1 0 44068 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_477
timestamp 1
transform 1 0 44988 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_496
timestamp 1
transform 1 0 46736 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_501
timestamp 1
transform 1 0 47196 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_505
timestamp 1
transform 1 0 47564 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_529
timestamp 1636968456
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_541
timestamp 1636968456
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_553
timestamp 1
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_559
timestamp 1
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_561
timestamp 1636968456
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_573
timestamp 1636968456
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_585
timestamp 1636968456
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_597
timestamp 1636968456
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_609
timestamp 1
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_615
timestamp 1
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_617
timestamp 1636968456
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_629
timestamp 1636968456
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_641
timestamp 1636968456
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_653
timestamp 1636968456
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_665
timestamp 1
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_671
timestamp 1
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_673
timestamp 1636968456
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_685
timestamp 1636968456
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_697
timestamp 1636968456
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_709
timestamp 1636968456
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_721
timestamp 1
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_727
timestamp 1
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_729
timestamp 1636968456
transform 1 0 68172 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_741
timestamp 1636968456
transform 1 0 69276 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_753
timestamp 1636968456
transform 1 0 70380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_765
timestamp 1636968456
transform 1 0 71484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_777
timestamp 1
transform 1 0 72588 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_783
timestamp 1
transform 1 0 73140 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_785
timestamp 1636968456
transform 1 0 73324 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_797
timestamp 1636968456
transform 1 0 74428 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_809
timestamp 1636968456
transform 1 0 75532 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_821
timestamp 1636968456
transform 1 0 76636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_833
timestamp 1
transform 1 0 77740 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_839
timestamp 1
transform 1 0 78292 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_841
timestamp 1
transform 1 0 78476 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_3
timestamp 1
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_11
timestamp 1636968456
transform 1 0 2116 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_23
timestamp 1
transform 1 0 3220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1636968456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1636968456
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1636968456
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1636968456
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1636968456
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1636968456
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1636968456
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1636968456
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1636968456
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1636968456
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1636968456
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1636968456
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1636968456
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1636968456
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1636968456
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1636968456
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1636968456
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1636968456
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_277
timestamp 1
transform 1 0 26588 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_305
timestamp 1
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_309
timestamp 1
transform 1 0 29532 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_315
timestamp 1
transform 1 0 30084 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_343
timestamp 1636968456
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_355
timestamp 1
transform 1 0 33764 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_377
timestamp 1
transform 1 0 35788 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_403
timestamp 1
transform 1 0 38180 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_418
timestamp 1
transform 1 0 39560 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_426
timestamp 1
transform 1 0 40296 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_438
timestamp 1636968456
transform 1 0 41400 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_450
timestamp 1
transform 1 0 42504 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_456
timestamp 1
transform 1 0 43056 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_463
timestamp 1636968456
transform 1 0 43700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_475
timestamp 1
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_479
timestamp 1636968456
transform 1 0 45172 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_491
timestamp 1636968456
transform 1 0 46276 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_503
timestamp 1636968456
transform 1 0 47380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_515
timestamp 1636968456
transform 1 0 48484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_527
timestamp 1
transform 1 0 49588 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_531
timestamp 1
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_533
timestamp 1636968456
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_545
timestamp 1636968456
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_557
timestamp 1636968456
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_569
timestamp 1636968456
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_581
timestamp 1
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_587
timestamp 1
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_589
timestamp 1636968456
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_601
timestamp 1636968456
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_613
timestamp 1636968456
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_625
timestamp 1636968456
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_637
timestamp 1
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_643
timestamp 1
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_645
timestamp 1636968456
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_657
timestamp 1636968456
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_669
timestamp 1636968456
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_681
timestamp 1636968456
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_693
timestamp 1
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_699
timestamp 1
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_701
timestamp 1636968456
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_713
timestamp 1636968456
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_725
timestamp 1636968456
transform 1 0 67804 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_737
timestamp 1636968456
transform 1 0 68908 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_749
timestamp 1
transform 1 0 70012 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_755
timestamp 1
transform 1 0 70564 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_757
timestamp 1636968456
transform 1 0 70748 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_769
timestamp 1636968456
transform 1 0 71852 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_781
timestamp 1636968456
transform 1 0 72956 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_793
timestamp 1636968456
transform 1 0 74060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_805
timestamp 1
transform 1 0 75164 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_811
timestamp 1
transform 1 0 75716 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_813
timestamp 1636968456
transform 1 0 75900 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_825
timestamp 1636968456
transform 1 0 77004 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_837
timestamp 1
transform 1 0 78108 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_841
timestamp 1
transform 1 0 78476 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_3
timestamp 1
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_14
timestamp 1636968456
transform 1 0 2392 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_26
timestamp 1636968456
transform 1 0 3496 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_38
timestamp 1636968456
transform 1 0 4600 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_50
timestamp 1
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1636968456
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1636968456
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1636968456
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1636968456
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1636968456
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1636968456
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1636968456
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1636968456
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1636968456
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1636968456
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1636968456
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1636968456
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1636968456
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1636968456
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1636968456
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1636968456
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1636968456
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_293
timestamp 1
transform 1 0 28060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_325
timestamp 1
transform 1 0 31004 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_333
timestamp 1
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_344
timestamp 1
transform 1 0 32752 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_372
timestamp 1
transform 1 0 35328 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_384
timestamp 1
transform 1 0 36432 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_401
timestamp 1
transform 1 0 37996 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_409
timestamp 1
transform 1 0 38732 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_432
timestamp 1636968456
transform 1 0 40848 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_444
timestamp 1
transform 1 0 41952 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_469
timestamp 1
transform 1 0 44252 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_481
timestamp 1636968456
transform 1 0 45356 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_493
timestamp 1
transform 1 0 46460 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_501
timestamp 1
transform 1 0 47196 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_505
timestamp 1636968456
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_517
timestamp 1636968456
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_529
timestamp 1636968456
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_541
timestamp 1636968456
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_553
timestamp 1
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_559
timestamp 1
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_561
timestamp 1636968456
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_573
timestamp 1636968456
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_585
timestamp 1636968456
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_597
timestamp 1636968456
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_609
timestamp 1
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_615
timestamp 1
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_617
timestamp 1636968456
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_629
timestamp 1636968456
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_641
timestamp 1636968456
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_653
timestamp 1636968456
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_665
timestamp 1
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_671
timestamp 1
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_673
timestamp 1636968456
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_685
timestamp 1636968456
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_697
timestamp 1636968456
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_709
timestamp 1636968456
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_721
timestamp 1
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_727
timestamp 1
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_729
timestamp 1636968456
transform 1 0 68172 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_741
timestamp 1636968456
transform 1 0 69276 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_753
timestamp 1636968456
transform 1 0 70380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_765
timestamp 1636968456
transform 1 0 71484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_777
timestamp 1
transform 1 0 72588 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_783
timestamp 1
transform 1 0 73140 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_785
timestamp 1636968456
transform 1 0 73324 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_797
timestamp 1636968456
transform 1 0 74428 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_809
timestamp 1636968456
transform 1 0 75532 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_821
timestamp 1636968456
transform 1 0 76636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_833
timestamp 1
transform 1 0 77740 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_839
timestamp 1
transform 1 0 78292 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_841
timestamp 1
transform 1 0 78476 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_3
timestamp 1
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_7
timestamp 1
transform 1 0 1748 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_11
timestamp 1636968456
transform 1 0 2116 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_23
timestamp 1
transform 1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1636968456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1636968456
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1636968456
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1636968456
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1636968456
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1636968456
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1636968456
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1636968456
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1636968456
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1636968456
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1636968456
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1636968456
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1636968456
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1636968456
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1636968456
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1636968456
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1636968456
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1636968456
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1636968456
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_289
timestamp 1
transform 1 0 27692 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_293
timestamp 1
transform 1 0 28060 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_317
timestamp 1
transform 1 0 30268 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_325
timestamp 1
transform 1 0 31004 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_347
timestamp 1636968456
transform 1 0 33028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_359
timestamp 1
transform 1 0 34132 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_371
timestamp 1
transform 1 0 35236 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_387
timestamp 1636968456
transform 1 0 36708 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_399
timestamp 1636968456
transform 1 0 37812 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_411
timestamp 1
transform 1 0 38916 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 1
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 1636968456
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_433
timestamp 1636968456
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_445
timestamp 1636968456
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_463
timestamp 1
transform 1 0 43700 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_474
timestamp 1
transform 1 0 44712 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_482
timestamp 1
transform 1 0 45448 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_490
timestamp 1636968456
transform 1 0 46184 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_502
timestamp 1636968456
transform 1 0 47288 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_514
timestamp 1636968456
transform 1 0 48392 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_526
timestamp 1
transform 1 0 49496 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_533
timestamp 1636968456
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_545
timestamp 1636968456
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_557
timestamp 1636968456
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_569
timestamp 1636968456
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_581
timestamp 1
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_587
timestamp 1
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_589
timestamp 1636968456
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_601
timestamp 1636968456
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_613
timestamp 1636968456
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_625
timestamp 1636968456
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_637
timestamp 1
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_643
timestamp 1
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_645
timestamp 1636968456
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_657
timestamp 1636968456
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_669
timestamp 1636968456
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_681
timestamp 1636968456
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_693
timestamp 1
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_699
timestamp 1
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_701
timestamp 1636968456
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_713
timestamp 1636968456
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_725
timestamp 1636968456
transform 1 0 67804 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_737
timestamp 1636968456
transform 1 0 68908 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_749
timestamp 1
transform 1 0 70012 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_755
timestamp 1
transform 1 0 70564 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_757
timestamp 1636968456
transform 1 0 70748 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_769
timestamp 1636968456
transform 1 0 71852 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_781
timestamp 1636968456
transform 1 0 72956 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_793
timestamp 1636968456
transform 1 0 74060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_805
timestamp 1
transform 1 0 75164 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_811
timestamp 1
transform 1 0 75716 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_813
timestamp 1636968456
transform 1 0 75900 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_825
timestamp 1636968456
transform 1 0 77004 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_837
timestamp 1
transform 1 0 78108 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_841
timestamp 1
transform 1 0 78476 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_3
timestamp 1
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_14
timestamp 1636968456
transform 1 0 2392 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_26
timestamp 1636968456
transform 1 0 3496 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_38
timestamp 1636968456
transform 1 0 4600 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_50
timestamp 1
transform 1 0 5704 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1636968456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1636968456
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1636968456
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1636968456
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1636968456
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1636968456
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1636968456
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1636968456
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1636968456
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1636968456
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1636968456
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1636968456
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1636968456
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1636968456
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1636968456
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1636968456
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1636968456
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1636968456
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1636968456
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1636968456
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_329
timestamp 1
transform 1 0 31372 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_345
timestamp 1636968456
transform 1 0 32844 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_357
timestamp 1636968456
transform 1 0 33948 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_369
timestamp 1
transform 1 0 35052 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_377
timestamp 1
transform 1 0 35788 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_393
timestamp 1
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_401
timestamp 1
transform 1 0 37996 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_406
timestamp 1636968456
transform 1 0 38456 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_418
timestamp 1
transform 1 0 39560 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_426
timestamp 1
transform 1 0 40296 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_442
timestamp 1
transform 1 0 41768 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 1636968456
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_461
timestamp 1
transform 1 0 43516 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_469
timestamp 1
transform 1 0 44252 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_476
timestamp 1
transform 1 0 44896 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_482
timestamp 1
transform 1 0 45448 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_507
timestamp 1636968456
transform 1 0 47748 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_519
timestamp 1636968456
transform 1 0 48852 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_531
timestamp 1636968456
transform 1 0 49956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_543
timestamp 1636968456
transform 1 0 51060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_555
timestamp 1
transform 1 0 52164 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_559
timestamp 1
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_561
timestamp 1636968456
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_573
timestamp 1636968456
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_585
timestamp 1636968456
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_597
timestamp 1636968456
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_609
timestamp 1
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_615
timestamp 1
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_617
timestamp 1636968456
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_629
timestamp 1636968456
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_641
timestamp 1636968456
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_653
timestamp 1636968456
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_665
timestamp 1
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_671
timestamp 1
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_673
timestamp 1636968456
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_685
timestamp 1636968456
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_697
timestamp 1636968456
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_709
timestamp 1636968456
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_721
timestamp 1
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_727
timestamp 1
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_729
timestamp 1636968456
transform 1 0 68172 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_741
timestamp 1636968456
transform 1 0 69276 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_753
timestamp 1636968456
transform 1 0 70380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_765
timestamp 1636968456
transform 1 0 71484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_777
timestamp 1
transform 1 0 72588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_783
timestamp 1
transform 1 0 73140 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_785
timestamp 1636968456
transform 1 0 73324 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_797
timestamp 1636968456
transform 1 0 74428 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_809
timestamp 1636968456
transform 1 0 75532 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_821
timestamp 1636968456
transform 1 0 76636 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_833
timestamp 1
transform 1 0 77740 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_839
timestamp 1
transform 1 0 78292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_841
timestamp 1
transform 1 0 78476 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_3
timestamp 1
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_18
timestamp 1
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_26
timestamp 1
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1636968456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1636968456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1636968456
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1636968456
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1636968456
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1636968456
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1636968456
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1636968456
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1636968456
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1636968456
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1636968456
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1636968456
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1636968456
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1636968456
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1636968456
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1636968456
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1636968456
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1636968456
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1636968456
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1636968456
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1636968456
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1636968456
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_333
timestamp 1
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_358
timestamp 1
transform 1 0 34040 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_371
timestamp 1
transform 1 0 35236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_421
timestamp 1
transform 1 0 39836 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_427
timestamp 1
transform 1 0 40388 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_451
timestamp 1
transform 1 0 42596 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_457
timestamp 1
transform 1 0 43148 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_474
timestamp 1
transform 1 0 44712 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_477
timestamp 1
transform 1 0 44988 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_485
timestamp 1
transform 1 0 45724 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_493
timestamp 1636968456
transform 1 0 46460 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_508
timestamp 1
transform 1 0 47840 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_516
timestamp 1
transform 1 0 48576 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_521
timestamp 1
transform 1 0 49036 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_529
timestamp 1
transform 1 0 49772 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_533
timestamp 1636968456
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_545
timestamp 1636968456
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_557
timestamp 1
transform 1 0 52348 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_564
timestamp 1
transform 1 0 52992 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_570
timestamp 1636968456
transform 1 0 53544 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_582
timestamp 1
transform 1 0 54648 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_589
timestamp 1636968456
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_601
timestamp 1636968456
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_613
timestamp 1
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_620
timestamp 1636968456
transform 1 0 58144 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_632
timestamp 1636968456
transform 1 0 59248 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_648
timestamp 1
transform 1 0 60720 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_654
timestamp 1636968456
transform 1 0 61272 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_666
timestamp 1
transform 1 0 62376 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_675
timestamp 1636968456
transform 1 0 63204 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_687
timestamp 1636968456
transform 1 0 64308 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_699
timestamp 1
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_701
timestamp 1636968456
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_713
timestamp 1636968456
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_725
timestamp 1
transform 1 0 67804 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_731
timestamp 1636968456
transform 1 0 68356 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_743
timestamp 1636968456
transform 1 0 69460 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_755
timestamp 1
transform 1 0 70564 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_757
timestamp 1636968456
transform 1 0 70748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_769
timestamp 1
transform 1 0 71852 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_774
timestamp 1636968456
transform 1 0 72312 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_786
timestamp 1636968456
transform 1 0 73416 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_798
timestamp 1636968456
transform 1 0 74520 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_810
timestamp 1
transform 1 0 75624 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_813
timestamp 1636968456
transform 1 0 75900 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_825
timestamp 1636968456
transform 1 0 77004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_837
timestamp 1
transform 1 0 78108 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_841
timestamp 1
transform 1 0 78476 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_3
timestamp 1
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_7
timestamp 1
transform 1 0 1748 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_11
timestamp 1636968456
transform 1 0 2116 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_23
timestamp 1636968456
transform 1 0 3220 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_35
timestamp 1636968456
transform 1 0 4324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_47
timestamp 1
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1636968456
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1636968456
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1636968456
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1636968456
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1636968456
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1636968456
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1636968456
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1636968456
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1636968456
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1636968456
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1636968456
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1636968456
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1636968456
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1636968456
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 1636968456
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 1636968456
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 1
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1636968456
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1636968456
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1636968456
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1636968456
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_337
timestamp 1
transform 1 0 32108 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_353
timestamp 1
transform 1 0 33580 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_379
timestamp 1
transform 1 0 35972 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_390
timestamp 1
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_393
timestamp 1
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_401
timestamp 1
transform 1 0 37996 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_423
timestamp 1
transform 1 0 40020 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_433
timestamp 1
transform 1 0 40940 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_493
timestamp 1
transform 1 0 46460 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_509
timestamp 1
transform 1 0 47932 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_522
timestamp 1
transform 1 0 49128 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_531
timestamp 1
transform 1 0 49956 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_565
timestamp 1
transform 1 0 53084 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_571
timestamp 1
transform 1 0 53636 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_601
timestamp 1
transform 1 0 56396 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_621
timestamp 1
transform 1 0 58236 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_637
timestamp 1
transform 1 0 59708 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_642
timestamp 1
transform 1 0 60168 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_655
timestamp 1
transform 1 0 61364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_664
timestamp 1
transform 1 0 62192 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_677
timestamp 1
transform 1 0 63388 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_733
timestamp 1
transform 1 0 68540 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_774
timestamp 1
transform 1 0 72312 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_783
timestamp 1
transform 1 0 73140 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_791
timestamp 1636968456
transform 1 0 73876 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_803
timestamp 1636968456
transform 1 0 74980 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_815
timestamp 1636968456
transform 1 0 76084 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_827
timestamp 1636968456
transform 1 0 77188 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_839
timestamp 1
transform 1 0 78292 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_841
timestamp 1
transform 1 0 78476 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1636968456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1636968456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1636968456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1636968456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_53
timestamp 1
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_57
timestamp 1636968456
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_69
timestamp 1636968456
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_81
timestamp 1
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1636968456
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1636968456
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_109
timestamp 1
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_113
timestamp 1636968456
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 1636968456
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 1
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1636968456
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1636968456
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_165
timestamp 1
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_169
timestamp 1636968456
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_181
timestamp 1636968456
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 1
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1636968456
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1636968456
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_221
timestamp 1
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_225
timestamp 1636968456
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_237
timestamp 1636968456
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_249
timestamp 1
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1636968456
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1636968456
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_277
timestamp 1
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_281
timestamp 1636968456
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_293
timestamp 1636968456
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_305
timestamp 1
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1636968456
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1636968456
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_333
timestamp 1
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_337
timestamp 1636968456
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_349
timestamp 1636968456
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_361
timestamp 1
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_365
timestamp 1
transform 1 0 34684 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_373
timestamp 1
transform 1 0 35420 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_384
timestamp 1
transform 1 0 36432 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_393
timestamp 1636968456
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_405
timestamp 1
transform 1 0 38364 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_415
timestamp 1
transform 1 0 39284 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 1
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_421
timestamp 1
transform 1 0 39836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_425
timestamp 1
transform 1 0 40204 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_432
timestamp 1636968456
transform 1 0 40848 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_444
timestamp 1
transform 1 0 41952 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_449
timestamp 1636968456
transform 1 0 42412 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_461
timestamp 1
transform 1 0 43516 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_471
timestamp 1
transform 1 0 44436 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_475
timestamp 1
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_477
timestamp 1
transform 1 0 44988 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_485
timestamp 1
transform 1 0 45724 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_499
timestamp 1
transform 1 0 47012 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_503
timestamp 1
transform 1 0 47380 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_505
timestamp 1636968456
transform 1 0 47564 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_517
timestamp 1636968456
transform 1 0 48668 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_529
timestamp 1
transform 1 0 49772 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_533
timestamp 1636968456
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_545
timestamp 1636968456
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_557
timestamp 1
transform 1 0 52348 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_561
timestamp 1636968456
transform 1 0 52716 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_573
timestamp 1636968456
transform 1 0 53820 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_585
timestamp 1
transform 1 0 54924 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_589
timestamp 1636968456
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_601
timestamp 1636968456
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_613
timestamp 1
transform 1 0 57500 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_617
timestamp 1636968456
transform 1 0 57868 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_629
timestamp 1636968456
transform 1 0 58972 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_641
timestamp 1
transform 1 0 60076 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_645
timestamp 1636968456
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_657
timestamp 1636968456
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_669
timestamp 1
transform 1 0 62652 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_673
timestamp 1636968456
transform 1 0 63020 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_685
timestamp 1636968456
transform 1 0 64124 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_697
timestamp 1
transform 1 0 65228 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_701
timestamp 1636968456
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_713
timestamp 1636968456
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_725
timestamp 1
transform 1 0 67804 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_729
timestamp 1636968456
transform 1 0 68172 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_741
timestamp 1636968456
transform 1 0 69276 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_753
timestamp 1
transform 1 0 70380 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_757
timestamp 1636968456
transform 1 0 70748 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_769
timestamp 1636968456
transform 1 0 71852 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_781
timestamp 1
transform 1 0 72956 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_785
timestamp 1636968456
transform 1 0 73324 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_797
timestamp 1636968456
transform 1 0 74428 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_809
timestamp 1
transform 1 0 75532 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_813
timestamp 1636968456
transform 1 0 75900 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_825
timestamp 1636968456
transform 1 0 77004 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_837
timestamp 1
transform 1 0 78108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_841
timestamp 1
transform 1 0 78476 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform 1 0 14260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 19780 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 18676 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 33212 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 42136 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 39652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 44528 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 10304 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform 1 0 55292 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 32568 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform 1 0 42412 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform 1 0 12144 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 37996 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 29256 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 29532 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 31556 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform 1 0 30360 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform 1 0 9844 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 22080 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 30268 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform 1 0 13432 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 13616 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform 1 0 9292 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 31372 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 19596 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 18216 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 14720 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 29348 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform 1 0 32200 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 20700 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 17480 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform -1 0 14996 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform -1 0 36892 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform -1 0 33120 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform -1 0 21160 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform -1 0 18584 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform -1 0 14812 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform -1 0 20240 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform 1 0 17572 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform -1 0 13524 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform -1 0 40204 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform -1 0 17020 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform -1 0 14352 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform -1 0 52440 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform -1 0 13524 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform -1 0 16192 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform -1 0 11500 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1
transform -1 0 19228 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1
transform -1 0 21068 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1
transform -1 0 48300 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1
transform -1 0 22540 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1
transform 1 0 46000 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1
transform -1 0 15272 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1
transform -1 0 14812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1
transform 1 0 14260 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1
transform -1 0 49588 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1
transform -1 0 19504 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1
transform 1 0 37628 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1
transform -1 0 36432 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1
transform 1 0 9752 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1
transform -1 0 32844 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1
transform -1 0 11408 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1
transform -1 0 12236 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1
transform -1 0 39652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1
transform 1 0 45172 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1
transform -1 0 38732 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1
transform -1 0 50232 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1
transform -1 0 21344 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1
transform -1 0 17480 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1
transform -1 0 50140 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1
transform 1 0 17020 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1
transform 1 0 32936 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1
transform -1 0 17388 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1
transform -1 0 53452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1
transform -1 0 40204 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1
transform 1 0 9476 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1
transform 1 0 35420 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1
transform -1 0 58328 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1
transform -1 0 39928 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1
transform -1 0 45816 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1
transform -1 0 34408 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1
transform -1 0 28060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1
transform -1 0 50048 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1
transform -1 0 55200 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1
transform -1 0 55108 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1
transform -1 0 36800 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1
transform -1 0 31464 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1
transform 1 0 38364 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1
transform -1 0 37996 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1
transform -1 0 44436 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1
transform -1 0 52624 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1
transform -1 0 43700 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1
transform -1 0 52440 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1
transform -1 0 47840 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1
transform -1 0 33396 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1
transform -1 0 50876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1
transform 1 0 41124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1
transform -1 0 35604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1
transform 1 0 32844 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1
transform -1 0 32844 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1
transform -1 0 44620 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1
transform -1 0 42044 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1
transform -1 0 39744 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1
transform 1 0 52716 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1
transform -1 0 50784 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1
transform -1 0 47472 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1
transform -1 0 41400 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1
transform -1 0 50324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1
transform -1 0 56764 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1
transform 1 0 41584 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1
transform -1 0 54556 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1
transform -1 0 41952 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1
transform -1 0 54372 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1
transform -1 0 37260 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1
transform -1 0 42228 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1
transform -1 0 47104 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1
transform -1 0 35420 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1
transform -1 0 42412 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1
transform -1 0 35420 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1
transform -1 0 39560 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1
transform -1 0 58604 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1
transform -1 0 39008 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1
transform 1 0 52992 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1
transform -1 0 37996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1
transform -1 0 54372 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1
transform -1 0 54372 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1
transform -1 0 44712 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1
transform -1 0 42044 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1
transform -1 0 36524 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1
transform -1 0 50048 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1
transform -1 0 53544 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1
transform -1 0 44896 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1
transform -1 0 57776 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1
transform -1 0 36432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1
transform -1 0 44804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1
transform -1 0 34684 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1
transform -1 0 43332 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1
transform -1 0 37996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1
transform -1 0 39928 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1
transform 1 0 55292 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1
transform -1 0 52532 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1
transform -1 0 33672 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1
transform -1 0 35420 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1
transform -1 0 34592 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1
transform -1 0 54740 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1
transform -1 0 31004 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1
transform -1 0 14260 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1
transform -1 0 14812 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1
transform 1 0 50600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 53176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform 1 0 59340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 54464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform -1 0 56672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1
transform -1 0 56856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1
transform 1 0 59984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1
transform 1 0 60628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1
transform 1 0 78108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1
transform -1 0 71208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1
transform 1 0 74152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1
transform 1 0 77372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1
transform 1 0 61272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1
transform 1 0 76084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1
transform -1 0 65412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1
transform -1 0 66056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1
transform 1 0 75440 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1
transform -1 0 67344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1
transform -1 0 72220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1
transform 1 0 74796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1
transform 1 0 73508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1
transform 1 0 71576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1
transform -1 0 67988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1
transform -1 0 58512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1
transform 1 0 77740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1
transform -1 0 69276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1
transform -1 0 52532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1
transform 1 0 69644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1
transform 1 0 70288 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1
transform 1 0 46184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1
transform -1 0 66700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1
transform -1 0 54188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1
transform -1 0 45632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1
transform -1 0 57776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1
transform 1 0 58696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1
transform -1 0 78568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1
transform -1 0 78384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1
transform -1 0 39284 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1
transform -1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1
transform -1 0 48760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1
transform 1 0 78016 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1
transform 1 0 39376 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output47
timestamp 1
transform 1 0 43884 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1
transform 1 0 78016 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output50
timestamp 1
transform 1 0 45172 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output51
timestamp 1
transform 1 0 46460 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1
transform -1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1
transform -1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1
transform 1 0 57868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1
transform 1 0 53544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1
transform 1 0 72864 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1
transform -1 0 51336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1
transform 1 0 61916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1
transform 1 0 51612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1
transform -1 0 68724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1
transform 1 0 63848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1
transform 1 0 49036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1
transform 1 0 49680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1
transform 1 0 63204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1
transform 1 0 64492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1
transform 1 0 76728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1
transform 1 0 78016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1
transform 1 0 62560 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1
transform 1 0 46460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1
transform 1 0 47748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1
transform -1 0 44896 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1
transform 1 0 78016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1
transform 1 0 78016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1
transform 1 0 78200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1
transform 1 0 78200 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1
transform 1 0 78016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_65
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 78844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_66
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 78844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_67
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 78844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_68
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 78844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_69
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 78844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_70
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 78844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_71
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 78844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_72
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 78844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_73
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 78844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_74
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 78844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_75
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 78844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_76
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 78844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_77
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 78844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_78
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 78844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_79
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 78844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_80
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 78844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_81
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 78844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_82
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 78844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_83
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 78844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_84
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 78844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_85
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 78844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_86
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 78844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_87
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 78844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_88
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 78844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_89
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 78844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_90
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 78844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_91
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 78844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_92
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 78844 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_93
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 78844 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_94
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 78844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_95
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 78844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_96
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 78844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_97
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 78844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_98
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 78844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_99
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 78844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_100
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 78844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_101
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 78844 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_102
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 78844 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_103
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 78844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_104
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 78844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_105
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 78844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_106
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 78844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_107
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 78844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_108
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 78844 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_109
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 78844 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_110
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 78844 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_111
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 78844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_112
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 78844 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_113
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 78844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_114
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1
transform -1 0 78844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_115
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1
transform -1 0 78844 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_116
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1
transform -1 0 78844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_117
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1
transform -1 0 78844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_118
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1
transform -1 0 78844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_119
timestamp 1
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1
transform -1 0 78844 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_120
timestamp 1
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1
transform -1 0 78844 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_121
timestamp 1
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1
transform -1 0 78844 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_122
timestamp 1
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1
transform -1 0 78844 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_123
timestamp 1
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1
transform -1 0 78844 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_124
timestamp 1
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1
transform -1 0 78844 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_125
timestamp 1
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1
transform -1 0 78844 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_126
timestamp 1
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1
transform -1 0 78844 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_127
timestamp 1
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1
transform -1 0 78844 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_128
timestamp 1
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1
transform -1 0 78844 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_129
timestamp 1
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1
transform -1 0 78844 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 1
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 1
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 1
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_143
timestamp 1
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_144
timestamp 1
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_145
timestamp 1
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_146
timestamp 1
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_147
timestamp 1
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_148
timestamp 1
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_149
timestamp 1
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_150
timestamp 1
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_151
timestamp 1
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_152
timestamp 1
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_153
timestamp 1
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_154
timestamp 1
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_155
timestamp 1
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_156
timestamp 1
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_157
timestamp 1
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_158
timestamp 1
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_159
timestamp 1
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_160
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_161
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_162
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_163
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_164
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_165
timestamp 1
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_166
timestamp 1
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_167
timestamp 1
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_168
timestamp 1
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_169
timestamp 1
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_170
timestamp 1
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_171
timestamp 1
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_172
timestamp 1
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_173
timestamp 1
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_174
timestamp 1
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_175
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_176
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_177
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_178
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_179
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_180
timestamp 1
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_181
timestamp 1
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_182
timestamp 1
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_183
timestamp 1
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_184
timestamp 1
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_185
timestamp 1
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_186
timestamp 1
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_187
timestamp 1
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_188
timestamp 1
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_189
timestamp 1
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_190
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_191
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_192
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_193
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_194
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_195
timestamp 1
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_196
timestamp 1
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_197
timestamp 1
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_198
timestamp 1
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_199
timestamp 1
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_200
timestamp 1
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_201
timestamp 1
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_202
timestamp 1
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_203
timestamp 1
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_204
timestamp 1
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_205
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_206
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_207
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_208
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_209
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_210
timestamp 1
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_211
timestamp 1
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_212
timestamp 1
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_213
timestamp 1
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_214
timestamp 1
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_215
timestamp 1
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_216
timestamp 1
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_217
timestamp 1
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_218
timestamp 1
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_219
timestamp 1
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_220
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_221
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_222
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_223
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_224
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_225
timestamp 1
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_226
timestamp 1
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_227
timestamp 1
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_228
timestamp 1
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_229
timestamp 1
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_230
timestamp 1
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_231
timestamp 1
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_232
timestamp 1
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_233
timestamp 1
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_234
timestamp 1
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_235
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_236
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_237
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_238
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_239
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_240
timestamp 1
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_241
timestamp 1
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_242
timestamp 1
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_243
timestamp 1
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_244
timestamp 1
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_245
timestamp 1
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_246
timestamp 1
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_247
timestamp 1
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_248
timestamp 1
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_249
timestamp 1
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_250
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_251
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_252
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_253
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_254
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_255
timestamp 1
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_256
timestamp 1
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_257
timestamp 1
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_258
timestamp 1
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_259
timestamp 1
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_260
timestamp 1
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_261
timestamp 1
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_262
timestamp 1
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_263
timestamp 1
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_264
timestamp 1
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_265
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_266
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_267
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_268
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_269
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_270
timestamp 1
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_271
timestamp 1
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_272
timestamp 1
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_273
timestamp 1
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_274
timestamp 1
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_275
timestamp 1
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_276
timestamp 1
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_277
timestamp 1
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_278
timestamp 1
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_279
timestamp 1
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_280
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_281
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_282
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_283
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_284
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_285
timestamp 1
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_286
timestamp 1
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_287
timestamp 1
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_288
timestamp 1
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_289
timestamp 1
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_290
timestamp 1
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_291
timestamp 1
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_292
timestamp 1
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_293
timestamp 1
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_294
timestamp 1
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_295
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_296
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_297
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_298
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_299
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_300
timestamp 1
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_301
timestamp 1
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_302
timestamp 1
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_303
timestamp 1
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_304
timestamp 1
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_305
timestamp 1
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_306
timestamp 1
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_307
timestamp 1
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_308
timestamp 1
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_309
timestamp 1
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_310
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_311
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_312
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_313
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_314
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_315
timestamp 1
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_316
timestamp 1
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_317
timestamp 1
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_318
timestamp 1
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_319
timestamp 1
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_320
timestamp 1
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_321
timestamp 1
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_322
timestamp 1
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_323
timestamp 1
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_324
timestamp 1
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_325
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_326
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_327
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_328
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_329
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_330
timestamp 1
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_331
timestamp 1
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_332
timestamp 1
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_333
timestamp 1
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_334
timestamp 1
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_335
timestamp 1
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_336
timestamp 1
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_337
timestamp 1
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_338
timestamp 1
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_339
timestamp 1
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_340
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_341
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_342
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_343
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_344
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_345
timestamp 1
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_346
timestamp 1
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_347
timestamp 1
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_348
timestamp 1
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_349
timestamp 1
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_350
timestamp 1
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_351
timestamp 1
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_352
timestamp 1
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_353
timestamp 1
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_354
timestamp 1
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_355
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_356
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_357
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_358
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_359
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_360
timestamp 1
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_361
timestamp 1
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_362
timestamp 1
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_363
timestamp 1
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_364
timestamp 1
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_365
timestamp 1
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_366
timestamp 1
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_367
timestamp 1
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_368
timestamp 1
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_369
timestamp 1
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_370
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_371
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_372
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_373
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_374
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_375
timestamp 1
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_376
timestamp 1
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_377
timestamp 1
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_378
timestamp 1
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_379
timestamp 1
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_380
timestamp 1
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_381
timestamp 1
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_382
timestamp 1
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_383
timestamp 1
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_384
timestamp 1
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_385
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_386
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_387
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_388
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_389
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_390
timestamp 1
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_391
timestamp 1
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_392
timestamp 1
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_393
timestamp 1
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_394
timestamp 1
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_395
timestamp 1
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_396
timestamp 1
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_397
timestamp 1
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_398
timestamp 1
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_399
timestamp 1
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_400
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_401
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_402
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_403
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_404
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_405
timestamp 1
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_406
timestamp 1
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_407
timestamp 1
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_408
timestamp 1
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_409
timestamp 1
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_410
timestamp 1
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_411
timestamp 1
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_412
timestamp 1
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_413
timestamp 1
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_414
timestamp 1
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_415
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_416
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_417
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_418
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_419
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_420
timestamp 1
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_421
timestamp 1
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_422
timestamp 1
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_423
timestamp 1
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_424
timestamp 1
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_425
timestamp 1
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_426
timestamp 1
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_427
timestamp 1
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_428
timestamp 1
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_429
timestamp 1
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_430
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_431
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_432
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_433
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_434
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_435
timestamp 1
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_436
timestamp 1
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_437
timestamp 1
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_438
timestamp 1
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_439
timestamp 1
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_440
timestamp 1
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_441
timestamp 1
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_442
timestamp 1
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_443
timestamp 1
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_444
timestamp 1
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_445
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_446
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_447
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_448
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_449
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_450
timestamp 1
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_451
timestamp 1
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_452
timestamp 1
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_453
timestamp 1
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_454
timestamp 1
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_455
timestamp 1
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_456
timestamp 1
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_457
timestamp 1
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_458
timestamp 1
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_459
timestamp 1
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_460
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_461
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_462
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_463
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_464
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_465
timestamp 1
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_466
timestamp 1
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_467
timestamp 1
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_468
timestamp 1
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_469
timestamp 1
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_470
timestamp 1
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_471
timestamp 1
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_472
timestamp 1
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_473
timestamp 1
transform 1 0 73232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_474
timestamp 1
transform 1 0 78384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_475
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_476
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_477
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_478
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_479
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_480
timestamp 1
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_481
timestamp 1
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_482
timestamp 1
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_483
timestamp 1
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_484
timestamp 1
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_485
timestamp 1
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_486
timestamp 1
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_487
timestamp 1
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_488
timestamp 1
transform 1 0 70656 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_489
timestamp 1
transform 1 0 75808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_490
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_491
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_492
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_493
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_494
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_495
timestamp 1
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_496
timestamp 1
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_497
timestamp 1
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_498
timestamp 1
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_499
timestamp 1
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_500
timestamp 1
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_501
timestamp 1
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_502
timestamp 1
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_503
timestamp 1
transform 1 0 73232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_504
timestamp 1
transform 1 0 78384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_505
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_506
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_507
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_508
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_509
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_510
timestamp 1
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_511
timestamp 1
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_512
timestamp 1
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_513
timestamp 1
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_514
timestamp 1
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_515
timestamp 1
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_516
timestamp 1
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_517
timestamp 1
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_518
timestamp 1
transform 1 0 70656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_519
timestamp 1
transform 1 0 75808 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_520
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_521
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_522
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_523
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_524
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_525
timestamp 1
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_526
timestamp 1
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_527
timestamp 1
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_528
timestamp 1
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_529
timestamp 1
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_530
timestamp 1
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_531
timestamp 1
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_532
timestamp 1
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_533
timestamp 1
transform 1 0 73232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_534
timestamp 1
transform 1 0 78384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_535
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_536
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_537
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_538
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_539
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_540
timestamp 1
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_541
timestamp 1
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_542
timestamp 1
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_543
timestamp 1
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_544
timestamp 1
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_545
timestamp 1
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_546
timestamp 1
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_547
timestamp 1
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_548
timestamp 1
transform 1 0 70656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_549
timestamp 1
transform 1 0 75808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_550
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_551
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_552
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_553
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_554
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_555
timestamp 1
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_556
timestamp 1
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_557
timestamp 1
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_558
timestamp 1
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_559
timestamp 1
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_560
timestamp 1
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_561
timestamp 1
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_562
timestamp 1
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_563
timestamp 1
transform 1 0 73232 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_564
timestamp 1
transform 1 0 78384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_565
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_566
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_567
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_568
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_569
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_570
timestamp 1
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_571
timestamp 1
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_572
timestamp 1
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_573
timestamp 1
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_574
timestamp 1
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_575
timestamp 1
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_576
timestamp 1
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_577
timestamp 1
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_578
timestamp 1
transform 1 0 70656 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_579
timestamp 1
transform 1 0 75808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_580
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_581
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_582
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_583
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_584
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_585
timestamp 1
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_586
timestamp 1
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_587
timestamp 1
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_588
timestamp 1
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_589
timestamp 1
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_590
timestamp 1
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_591
timestamp 1
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_592
timestamp 1
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_593
timestamp 1
transform 1 0 73232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_594
timestamp 1
transform 1 0 78384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_595
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_596
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_597
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_598
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_599
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_600
timestamp 1
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_601
timestamp 1
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_602
timestamp 1
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_603
timestamp 1
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_604
timestamp 1
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_605
timestamp 1
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_606
timestamp 1
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_607
timestamp 1
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_608
timestamp 1
transform 1 0 70656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_609
timestamp 1
transform 1 0 75808 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_610
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_611
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_612
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_613
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_614
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_615
timestamp 1
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_616
timestamp 1
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_617
timestamp 1
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_618
timestamp 1
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_619
timestamp 1
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_620
timestamp 1
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_621
timestamp 1
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_622
timestamp 1
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_623
timestamp 1
transform 1 0 73232 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_624
timestamp 1
transform 1 0 78384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_625
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_626
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_627
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_628
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_629
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_630
timestamp 1
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_631
timestamp 1
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_632
timestamp 1
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_633
timestamp 1
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_634
timestamp 1
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_635
timestamp 1
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_636
timestamp 1
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_637
timestamp 1
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_638
timestamp 1
transform 1 0 70656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_639
timestamp 1
transform 1 0 75808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_640
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_641
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_642
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_643
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_644
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_645
timestamp 1
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_646
timestamp 1
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_647
timestamp 1
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_648
timestamp 1
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_649
timestamp 1
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_650
timestamp 1
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_651
timestamp 1
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_652
timestamp 1
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_653
timestamp 1
transform 1 0 73232 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_654
timestamp 1
transform 1 0 78384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_655
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_656
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_657
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_658
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_659
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_660
timestamp 1
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_661
timestamp 1
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_662
timestamp 1
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_663
timestamp 1
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_664
timestamp 1
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_665
timestamp 1
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_666
timestamp 1
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_667
timestamp 1
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_668
timestamp 1
transform 1 0 70656 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_669
timestamp 1
transform 1 0 75808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_670
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_671
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_672
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_673
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_674
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_675
timestamp 1
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_676
timestamp 1
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_677
timestamp 1
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_678
timestamp 1
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_679
timestamp 1
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_680
timestamp 1
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_681
timestamp 1
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_682
timestamp 1
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_683
timestamp 1
transform 1 0 73232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_684
timestamp 1
transform 1 0 78384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_685
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_686
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_687
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_688
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_689
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_690
timestamp 1
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_691
timestamp 1
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_692
timestamp 1
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_693
timestamp 1
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_694
timestamp 1
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_695
timestamp 1
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_696
timestamp 1
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_697
timestamp 1
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_698
timestamp 1
transform 1 0 70656 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_699
timestamp 1
transform 1 0 75808 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_700
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_701
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_702
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_703
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_704
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_705
timestamp 1
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_706
timestamp 1
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_707
timestamp 1
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_708
timestamp 1
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_709
timestamp 1
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_710
timestamp 1
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_711
timestamp 1
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_712
timestamp 1
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_713
timestamp 1
transform 1 0 73232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_714
timestamp 1
transform 1 0 78384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_715
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_716
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_717
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_718
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_719
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_720
timestamp 1
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_721
timestamp 1
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_722
timestamp 1
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_723
timestamp 1
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_724
timestamp 1
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_725
timestamp 1
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_726
timestamp 1
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_727
timestamp 1
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_728
timestamp 1
transform 1 0 70656 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_729
timestamp 1
transform 1 0 75808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_730
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_731
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_732
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_733
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_734
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_735
timestamp 1
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_736
timestamp 1
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_737
timestamp 1
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_738
timestamp 1
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_739
timestamp 1
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_740
timestamp 1
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_741
timestamp 1
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_742
timestamp 1
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_743
timestamp 1
transform 1 0 73232 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_744
timestamp 1
transform 1 0 78384 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_745
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_746
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_747
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_748
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_749
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_750
timestamp 1
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_751
timestamp 1
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_752
timestamp 1
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_753
timestamp 1
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_754
timestamp 1
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_755
timestamp 1
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_756
timestamp 1
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_757
timestamp 1
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_758
timestamp 1
transform 1 0 70656 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_759
timestamp 1
transform 1 0 75808 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_760
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_761
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_762
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_763
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_764
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_765
timestamp 1
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_766
timestamp 1
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_767
timestamp 1
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_768
timestamp 1
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_769
timestamp 1
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_770
timestamp 1
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_771
timestamp 1
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_772
timestamp 1
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_773
timestamp 1
transform 1 0 73232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_774
timestamp 1
transform 1 0 78384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_775
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_776
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_777
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_778
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_779
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_780
timestamp 1
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_781
timestamp 1
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_782
timestamp 1
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_783
timestamp 1
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_784
timestamp 1
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_785
timestamp 1
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_786
timestamp 1
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_787
timestamp 1
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_788
timestamp 1
transform 1 0 70656 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_789
timestamp 1
transform 1 0 75808 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_790
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_791
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_792
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_793
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_794
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_795
timestamp 1
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_796
timestamp 1
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_797
timestamp 1
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_798
timestamp 1
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_799
timestamp 1
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_800
timestamp 1
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_801
timestamp 1
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_802
timestamp 1
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_803
timestamp 1
transform 1 0 73232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_804
timestamp 1
transform 1 0 78384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_805
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_806
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_807
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_808
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_809
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_810
timestamp 1
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_811
timestamp 1
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_812
timestamp 1
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_813
timestamp 1
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_814
timestamp 1
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_815
timestamp 1
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_816
timestamp 1
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_817
timestamp 1
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_818
timestamp 1
transform 1 0 70656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_819
timestamp 1
transform 1 0 75808 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_820
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_821
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_822
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_823
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_824
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_825
timestamp 1
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_826
timestamp 1
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_827
timestamp 1
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_828
timestamp 1
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_829
timestamp 1
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_830
timestamp 1
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_831
timestamp 1
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_832
timestamp 1
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_833
timestamp 1
transform 1 0 73232 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_834
timestamp 1
transform 1 0 78384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_835
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_836
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_837
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_838
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_839
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_840
timestamp 1
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_841
timestamp 1
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_842
timestamp 1
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_843
timestamp 1
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_844
timestamp 1
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_845
timestamp 1
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_846
timestamp 1
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_847
timestamp 1
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_848
timestamp 1
transform 1 0 70656 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_849
timestamp 1
transform 1 0 75808 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_850
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_851
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_852
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_853
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_854
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_855
timestamp 1
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_856
timestamp 1
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_857
timestamp 1
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_858
timestamp 1
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_859
timestamp 1
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_860
timestamp 1
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_861
timestamp 1
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_862
timestamp 1
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_863
timestamp 1
transform 1 0 73232 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_864
timestamp 1
transform 1 0 78384 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_865
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_866
timestamp 1
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_867
timestamp 1
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_868
timestamp 1
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_869
timestamp 1
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_870
timestamp 1
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_871
timestamp 1
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_872
timestamp 1
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_873
timestamp 1
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_874
timestamp 1
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_875
timestamp 1
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_876
timestamp 1
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_877
timestamp 1
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_878
timestamp 1
transform 1 0 70656 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_879
timestamp 1
transform 1 0 75808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_880
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_881
timestamp 1
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_882
timestamp 1
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_883
timestamp 1
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_884
timestamp 1
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_885
timestamp 1
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_886
timestamp 1
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_887
timestamp 1
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_888
timestamp 1
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_889
timestamp 1
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_890
timestamp 1
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_891
timestamp 1
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_892
timestamp 1
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_893
timestamp 1
transform 1 0 73232 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_894
timestamp 1
transform 1 0 78384 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_895
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_896
timestamp 1
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_897
timestamp 1
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_898
timestamp 1
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_899
timestamp 1
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_900
timestamp 1
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_901
timestamp 1
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_902
timestamp 1
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_903
timestamp 1
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_904
timestamp 1
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_905
timestamp 1
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_906
timestamp 1
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_907
timestamp 1
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_908
timestamp 1
transform 1 0 70656 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_909
timestamp 1
transform 1 0 75808 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_910
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_911
timestamp 1
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_912
timestamp 1
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_913
timestamp 1
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_914
timestamp 1
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_915
timestamp 1
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_916
timestamp 1
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_917
timestamp 1
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_918
timestamp 1
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_919
timestamp 1
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_920
timestamp 1
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_921
timestamp 1
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_922
timestamp 1
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_923
timestamp 1
transform 1 0 73232 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_924
timestamp 1
transform 1 0 78384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_925
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_926
timestamp 1
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_927
timestamp 1
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_928
timestamp 1
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_929
timestamp 1
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_930
timestamp 1
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_931
timestamp 1
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_932
timestamp 1
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_933
timestamp 1
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_934
timestamp 1
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_935
timestamp 1
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_936
timestamp 1
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_937
timestamp 1
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_938
timestamp 1
transform 1 0 70656 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_939
timestamp 1
transform 1 0 75808 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_940
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_941
timestamp 1
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_942
timestamp 1
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_943
timestamp 1
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_944
timestamp 1
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_945
timestamp 1
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_946
timestamp 1
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_947
timestamp 1
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_948
timestamp 1
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_949
timestamp 1
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_950
timestamp 1
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_951
timestamp 1
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_952
timestamp 1
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_953
timestamp 1
transform 1 0 73232 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_954
timestamp 1
transform 1 0 78384 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_955
timestamp 1
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_956
timestamp 1
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_957
timestamp 1
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_958
timestamp 1
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_959
timestamp 1
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_960
timestamp 1
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_961
timestamp 1
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_962
timestamp 1
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_963
timestamp 1
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_964
timestamp 1
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_965
timestamp 1
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_966
timestamp 1
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_967
timestamp 1
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_968
timestamp 1
transform 1 0 70656 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_969
timestamp 1
transform 1 0 75808 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_970
timestamp 1
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_971
timestamp 1
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_972
timestamp 1
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_973
timestamp 1
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_974
timestamp 1
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_975
timestamp 1
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_976
timestamp 1
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_977
timestamp 1
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_978
timestamp 1
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_979
timestamp 1
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_980
timestamp 1
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_981
timestamp 1
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_982
timestamp 1
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_983
timestamp 1
transform 1 0 73232 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_984
timestamp 1
transform 1 0 78384 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_985
timestamp 1
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_986
timestamp 1
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_987
timestamp 1
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_988
timestamp 1
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_989
timestamp 1
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_990
timestamp 1
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_991
timestamp 1
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_992
timestamp 1
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_993
timestamp 1
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_994
timestamp 1
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_995
timestamp 1
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_996
timestamp 1
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_997
timestamp 1
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_998
timestamp 1
transform 1 0 70656 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_999
timestamp 1
transform 1 0 75808 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1000
timestamp 1
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1001
timestamp 1
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1002
timestamp 1
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1003
timestamp 1
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1004
timestamp 1
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1005
timestamp 1
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1006
timestamp 1
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1007
timestamp 1
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1008
timestamp 1
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1009
timestamp 1
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1010
timestamp 1
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1011
timestamp 1
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1012
timestamp 1
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1013
timestamp 1
transform 1 0 73232 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1014
timestamp 1
transform 1 0 78384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1015
timestamp 1
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1016
timestamp 1
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1017
timestamp 1
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1018
timestamp 1
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1019
timestamp 1
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1020
timestamp 1
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1021
timestamp 1
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1022
timestamp 1
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1023
timestamp 1
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1024
timestamp 1
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1025
timestamp 1
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1026
timestamp 1
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1027
timestamp 1
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1028
timestamp 1
transform 1 0 70656 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1029
timestamp 1
transform 1 0 75808 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1030
timestamp 1
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1031
timestamp 1
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1032
timestamp 1
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1033
timestamp 1
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1034
timestamp 1
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1035
timestamp 1
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1036
timestamp 1
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1037
timestamp 1
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1038
timestamp 1
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1039
timestamp 1
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1040
timestamp 1
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1041
timestamp 1
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1042
timestamp 1
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1043
timestamp 1
transform 1 0 73232 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1044
timestamp 1
transform 1 0 78384 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1045
timestamp 1
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1046
timestamp 1
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1047
timestamp 1
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1048
timestamp 1
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1049
timestamp 1
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1050
timestamp 1
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1051
timestamp 1
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1052
timestamp 1
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1053
timestamp 1
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1054
timestamp 1
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1055
timestamp 1
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1056
timestamp 1
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1057
timestamp 1
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1058
timestamp 1
transform 1 0 70656 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1059
timestamp 1
transform 1 0 75808 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1060
timestamp 1
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1061
timestamp 1
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1062
timestamp 1
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1063
timestamp 1
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1064
timestamp 1
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1065
timestamp 1
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1066
timestamp 1
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1067
timestamp 1
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1068
timestamp 1
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1069
timestamp 1
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1070
timestamp 1
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1071
timestamp 1
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1072
timestamp 1
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1073
timestamp 1
transform 1 0 73232 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1074
timestamp 1
transform 1 0 78384 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1075
timestamp 1
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1076
timestamp 1
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1077
timestamp 1
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1078
timestamp 1
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1079
timestamp 1
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1080
timestamp 1
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1081
timestamp 1
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1082
timestamp 1
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1083
timestamp 1
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1084
timestamp 1
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1085
timestamp 1
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1086
timestamp 1
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1087
timestamp 1
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1088
timestamp 1
transform 1 0 70656 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1089
timestamp 1
transform 1 0 75808 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1090
timestamp 1
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1091
timestamp 1
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1092
timestamp 1
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1093
timestamp 1
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1094
timestamp 1
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1095
timestamp 1
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1096
timestamp 1
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1097
timestamp 1
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1098
timestamp 1
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1099
timestamp 1
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1100
timestamp 1
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1101
timestamp 1
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1102
timestamp 1
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1103
timestamp 1
transform 1 0 73232 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1104
timestamp 1
transform 1 0 78384 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1105
timestamp 1
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1106
timestamp 1
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1107
timestamp 1
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1108
timestamp 1
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1109
timestamp 1
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1110
timestamp 1
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1111
timestamp 1
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1112
timestamp 1
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1113
timestamp 1
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1114
timestamp 1
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1115
timestamp 1
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1116
timestamp 1
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1117
timestamp 1
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1118
timestamp 1
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1119
timestamp 1
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1120
timestamp 1
transform 1 0 42320 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1121
timestamp 1
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1122
timestamp 1
transform 1 0 47472 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1123
timestamp 1
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1124
timestamp 1
transform 1 0 52624 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1125
timestamp 1
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1126
timestamp 1
transform 1 0 57776 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1127
timestamp 1
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1128
timestamp 1
transform 1 0 62928 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1129
timestamp 1
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1130
timestamp 1
transform 1 0 68080 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1131
timestamp 1
transform 1 0 70656 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1132
timestamp 1
transform 1 0 73232 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1133
timestamp 1
transform 1 0 75808 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1134
timestamp 1
transform 1 0 78384 0 1 36992
box -38 -48 130 592
<< labels >>
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 gpio_in[0]
port 0 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 gpio_in[10]
port 1 nsew signal input
flabel metal2 s 79874 0 79930 800 0 FreeSans 224 90 0 0 gpio_in[11]
port 2 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 gpio_in[12]
port 3 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 gpio_in[13]
port 4 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 gpio_in[14]
port 5 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 gpio_in[15]
port 6 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 gpio_in[16]
port 7 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 gpio_in[17]
port 8 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 gpio_in[18]
port 9 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 gpio_in[19]
port 10 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 gpio_in[1]
port 11 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 gpio_in[20]
port 12 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpio_in[21]
port 13 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 gpio_in[22]
port 14 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 gpio_in[23]
port 15 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 gpio_in[24]
port 16 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 gpio_in[25]
port 17 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 gpio_in[26]
port 18 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 gpio_in[27]
port 19 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gpio_in[28]
port 20 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 gpio_in[29]
port 21 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 gpio_in[2]
port 22 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 gpio_in[30]
port 23 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 gpio_in[31]
port 24 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 gpio_in[32]
port 25 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 gpio_in[33]
port 26 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 gpio_in[34]
port 27 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 gpio_in[35]
port 28 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 gpio_in[36]
port 29 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 gpio_in[37]
port 30 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpio_in[3]
port 31 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gpio_in[4]
port 32 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 gpio_in[5]
port 33 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 gpio_in[6]
port 34 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 gpio_in[7]
port 35 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 gpio_in[8]
port 36 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 gpio_in[9]
port 37 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 gpio_oeb[0]
port 38 nsew signal output
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 gpio_oeb[10]
port 39 nsew signal output
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 gpio_oeb[11]
port 40 nsew signal output
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 gpio_oeb[12]
port 41 nsew signal output
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 gpio_oeb[13]
port 42 nsew signal output
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 gpio_oeb[14]
port 43 nsew signal output
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 gpio_oeb[15]
port 44 nsew signal output
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 gpio_oeb[16]
port 45 nsew signal output
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 gpio_oeb[17]
port 46 nsew signal output
flabel metal2 s 39946 39200 40002 40000 0 FreeSans 224 90 0 0 gpio_oeb[18]
port 47 nsew signal output
flabel metal2 s 73434 39200 73490 40000 0 FreeSans 224 90 0 0 gpio_oeb[19]
port 48 nsew signal output
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 gpio_oeb[1]
port 49 nsew signal output
flabel metal2 s 55402 39200 55458 40000 0 FreeSans 224 90 0 0 gpio_oeb[20]
port 50 nsew signal output
flabel metal2 s 51538 39200 51594 40000 0 FreeSans 224 90 0 0 gpio_oeb[21]
port 51 nsew signal output
flabel metal2 s 41234 39200 41290 40000 0 FreeSans 224 90 0 0 gpio_oeb[22]
port 52 nsew signal output
flabel metal2 s 68282 39200 68338 40000 0 FreeSans 224 90 0 0 gpio_oeb[23]
port 53 nsew signal output
flabel metal2 s 58622 39200 58678 40000 0 FreeSans 224 90 0 0 gpio_oeb[24]
port 54 nsew signal output
flabel metal2 s 48962 39200 49018 40000 0 FreeSans 224 90 0 0 gpio_oeb[25]
port 55 nsew signal output
flabel metal2 s 59266 39200 59322 40000 0 FreeSans 224 90 0 0 gpio_oeb[26]
port 56 nsew signal output
flabel metal2 s 59910 39200 59966 40000 0 FreeSans 224 90 0 0 gpio_oeb[27]
port 57 nsew signal output
flabel metal2 s 45742 39200 45798 40000 0 FreeSans 224 90 0 0 gpio_oeb[28]
port 58 nsew signal output
flabel metal2 s 56046 39200 56102 40000 0 FreeSans 224 90 0 0 gpio_oeb[29]
port 59 nsew signal output
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 gpio_oeb[2]
port 60 nsew signal output
flabel metal2 s 54114 39200 54170 40000 0 FreeSans 224 90 0 0 gpio_oeb[30]
port 61 nsew signal output
flabel metal2 s 56690 39200 56746 40000 0 FreeSans 224 90 0 0 gpio_oeb[31]
port 62 nsew signal output
flabel metal2 s 60554 39200 60610 40000 0 FreeSans 224 90 0 0 gpio_oeb[32]
port 63 nsew signal output
flabel metal2 s 50894 39200 50950 40000 0 FreeSans 224 90 0 0 gpio_oeb[33]
port 64 nsew signal output
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 gpio_oeb[34]
port 65 nsew signal output
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 gpio_oeb[35]
port 66 nsew signal output
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 gpio_oeb[36]
port 67 nsew signal output
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 gpio_oeb[37]
port 68 nsew signal output
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 gpio_oeb[3]
port 69 nsew signal output
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 gpio_oeb[4]
port 70 nsew signal output
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 gpio_oeb[5]
port 71 nsew signal output
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 gpio_oeb[6]
port 72 nsew signal output
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 gpio_oeb[7]
port 73 nsew signal output
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 gpio_oeb[8]
port 74 nsew signal output
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 gpio_oeb[9]
port 75 nsew signal output
flabel metal2 s 43166 39200 43222 40000 0 FreeSans 224 90 0 0 gpio_out[0]
port 76 nsew signal output
flabel metal2 s 61198 39200 61254 40000 0 FreeSans 224 90 0 0 gpio_out[10]
port 77 nsew signal output
flabel metal2 s 42522 39200 42578 40000 0 FreeSans 224 90 0 0 gpio_out[11]
port 78 nsew signal output
flabel metal2 s 44454 39200 44510 40000 0 FreeSans 224 90 0 0 gpio_out[12]
port 79 nsew signal output
flabel metal2 s 52182 39200 52238 40000 0 FreeSans 224 90 0 0 gpio_out[13]
port 80 nsew signal output
flabel metal2 s 69570 39200 69626 40000 0 FreeSans 224 90 0 0 gpio_out[14]
port 81 nsew signal output
flabel metal2 s 61842 39200 61898 40000 0 FreeSans 224 90 0 0 gpio_out[15]
port 82 nsew signal output
flabel metal2 s 62486 39200 62542 40000 0 FreeSans 224 90 0 0 gpio_out[16]
port 83 nsew signal output
flabel metal2 s 63130 39200 63186 40000 0 FreeSans 224 90 0 0 gpio_out[17]
port 84 nsew signal output
flabel metal2 s 38658 39200 38714 40000 0 FreeSans 224 90 0 0 gpio_out[18]
port 85 nsew signal output
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 gpio_out[19]
port 86 nsew signal output
flabel metal2 s 41878 39200 41934 40000 0 FreeSans 224 90 0 0 gpio_out[1]
port 87 nsew signal output
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 gpio_out[20]
port 88 nsew signal output
flabel metal3 s 79200 17008 80000 17128 0 FreeSans 480 0 0 0 gpio_out[21]
port 89 nsew signal output
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 gpio_out[22]
port 90 nsew signal output
flabel metal2 s 43810 39200 43866 40000 0 FreeSans 224 90 0 0 gpio_out[23]
port 91 nsew signal output
flabel metal3 s 79200 23128 80000 23248 0 FreeSans 480 0 0 0 gpio_out[24]
port 92 nsew signal output
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 gpio_out[25]
port 93 nsew signal output
flabel metal2 s 45098 39200 45154 40000 0 FreeSans 224 90 0 0 gpio_out[26]
port 94 nsew signal output
flabel metal2 s 63774 39200 63830 40000 0 FreeSans 224 90 0 0 gpio_out[27]
port 95 nsew signal output
flabel metal2 s 46386 39200 46442 40000 0 FreeSans 224 90 0 0 gpio_out[28]
port 96 nsew signal output
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gpio_out[29]
port 97 nsew signal output
flabel metal2 s 70858 39200 70914 40000 0 FreeSans 224 90 0 0 gpio_out[2]
port 98 nsew signal output
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 gpio_out[30]
port 99 nsew signal output
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 gpio_out[31]
port 100 nsew signal output
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 gpio_out[32]
port 101 nsew signal output
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 gpio_out[33]
port 102 nsew signal output
flabel metal2 s 49606 39200 49662 40000 0 FreeSans 224 90 0 0 gpio_out[34]
port 103 nsew signal output
flabel metal2 s 67638 39200 67694 40000 0 FreeSans 224 90 0 0 gpio_out[35]
port 104 nsew signal output
flabel metal2 s 53470 39200 53526 40000 0 FreeSans 224 90 0 0 gpio_out[36]
port 105 nsew signal output
flabel metal2 s 57978 39200 58034 40000 0 FreeSans 224 90 0 0 gpio_out[37]
port 106 nsew signal output
flabel metal2 s 47030 39200 47086 40000 0 FreeSans 224 90 0 0 gpio_out[3]
port 107 nsew signal output
flabel metal2 s 66994 39200 67050 40000 0 FreeSans 224 90 0 0 gpio_out[4]
port 108 nsew signal output
flabel metal2 s 52826 39200 52882 40000 0 FreeSans 224 90 0 0 gpio_out[5]
port 109 nsew signal output
flabel metal2 s 72146 39200 72202 40000 0 FreeSans 224 90 0 0 gpio_out[6]
port 110 nsew signal output
flabel metal2 s 64418 39200 64474 40000 0 FreeSans 224 90 0 0 gpio_out[7]
port 111 nsew signal output
flabel metal2 s 40590 39200 40646 40000 0 FreeSans 224 90 0 0 gpio_out[8]
port 112 nsew signal output
flabel metal2 s 71502 39200 71558 40000 0 FreeSans 224 90 0 0 gpio_out[9]
port 113 nsew signal output
flabel metal2 s 47674 39200 47730 40000 0 FreeSans 224 90 0 0 irq[0]
port 114 nsew signal output
flabel metal2 s 48318 39200 48374 40000 0 FreeSans 224 90 0 0 irq[1]
port 115 nsew signal output
flabel metal2 s 65062 39200 65118 40000 0 FreeSans 224 90 0 0 irq[2]
port 116 nsew signal output
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 117 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 117 nsew power bidirectional
flabel metal4 s 65648 2128 65968 37584 0 FreeSans 1920 90 0 0 vccd1
port 117 nsew power bidirectional
flabel metal4 s 4868 2128 5188 37584 0 FreeSans 1920 90 0 0 vssd1
port 118 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 37584 0 FreeSans 1920 90 0 0 vssd1
port 118 nsew ground bidirectional
flabel metal4 s 66308 2128 66628 37584 0 FreeSans 1920 90 0 0 vssd1
port 118 nsew ground bidirectional
flabel metal2 s 39302 39200 39358 40000 0 FreeSans 224 90 0 0 wb_clk_i
port 119 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 wb_rst_i
port 120 nsew signal input
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 121 nsew signal output
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 122 nsew signal input
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 123 nsew signal input
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 124 nsew signal input
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 125 nsew signal input
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 126 nsew signal input
flabel metal2 s 59910 0 59966 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 127 nsew signal input
flabel metal2 s 60554 0 60610 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 128 nsew signal input
flabel metal2 s 79230 0 79286 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 129 nsew signal input
flabel metal2 s 70858 0 70914 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 130 nsew signal input
flabel metal2 s 74078 0 74134 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 131 nsew signal input
flabel metal2 s 77298 0 77354 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 132 nsew signal input
flabel metal2 s 61198 0 61254 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 133 nsew signal input
flabel metal2 s 76010 0 76066 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 134 nsew signal input
flabel metal2 s 65062 0 65118 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 135 nsew signal input
flabel metal2 s 65706 0 65762 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 136 nsew signal input
flabel metal2 s 75366 0 75422 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 137 nsew signal input
flabel metal2 s 66994 0 67050 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 138 nsew signal input
flabel metal2 s 72146 0 72202 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 139 nsew signal input
flabel metal2 s 74722 0 74778 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 140 nsew signal input
flabel metal2 s 73434 0 73490 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 141 nsew signal input
flabel metal2 s 71502 0 71558 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 142 nsew signal input
flabel metal2 s 67638 0 67694 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 143 nsew signal input
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 144 nsew signal input
flabel metal2 s 77942 0 77998 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 145 nsew signal input
flabel metal2 s 68926 0 68982 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 146 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 147 nsew signal input
flabel metal2 s 69570 0 69626 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 148 nsew signal input
flabel metal2 s 70214 0 70270 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 149 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 150 nsew signal input
flabel metal2 s 66350 0 66406 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 151 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 152 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 153 nsew signal input
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 154 nsew signal input
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 155 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 156 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 157 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 158 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 159 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 160 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 161 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 162 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 163 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 164 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 165 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 166 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 167 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 168 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 169 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 170 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 171 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 172 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 173 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 174 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 175 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 176 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 177 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 178 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 179 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 180 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 181 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 182 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 183 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 184 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 185 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 186 nsew signal input
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 187 nsew signal output
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 188 nsew signal output
flabel metal2 s 72790 0 72846 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 189 nsew signal output
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 190 nsew signal output
flabel metal2 s 61842 0 61898 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 191 nsew signal output
flabel metal2 s 70214 39200 70270 40000 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 192 nsew signal output
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 193 nsew signal output
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 194 nsew signal output
flabel metal2 s 54758 39200 54814 40000 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 195 nsew signal output
flabel metal2 s 63774 0 63830 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 196 nsew signal output
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 197 nsew signal output
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 198 nsew signal output
flabel metal2 s 50250 39200 50306 40000 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 199 nsew signal output
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 200 nsew signal output
flabel metal2 s 57334 39200 57390 40000 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 201 nsew signal output
flabel metal2 s 63130 0 63186 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 202 nsew signal output
flabel metal2 s 68926 39200 68982 40000 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 203 nsew signal output
flabel metal2 s 64418 0 64474 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 204 nsew signal output
flabel metal2 s 76654 0 76710 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 205 nsew signal output
flabel metal2 s 78586 0 78642 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 206 nsew signal output
flabel metal2 s 62486 0 62542 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 207 nsew signal output
flabel metal2 s 65706 39200 65762 40000 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 208 nsew signal output
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 209 nsew signal output
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 210 nsew signal output
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 211 nsew signal output
flabel metal3 s 79200 6808 80000 6928 0 FreeSans 480 0 0 0 wbs_dat_o[3]
port 212 nsew signal output
flabel metal2 s 66350 39200 66406 40000 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 213 nsew signal output
flabel metal3 s 79200 8168 80000 8288 0 FreeSans 480 0 0 0 wbs_dat_o[5]
port 214 nsew signal output
flabel metal3 s 79200 5448 80000 5568 0 FreeSans 480 0 0 0 wbs_dat_o[6]
port 215 nsew signal output
flabel metal3 s 79200 7488 80000 7608 0 FreeSans 480 0 0 0 wbs_dat_o[7]
port 216 nsew signal output
flabel metal2 s 72790 39200 72846 40000 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 217 nsew signal output
flabel metal3 s 79200 6128 80000 6248 0 FreeSans 480 0 0 0 wbs_dat_o[9]
port 218 nsew signal output
flabel metal3 s 79200 8 80000 128 0 FreeSans 480 0 0 0 wbs_sel_i[0]
port 219 nsew signal input
flabel metal3 s 79200 688 80000 808 0 FreeSans 480 0 0 0 wbs_sel_i[1]
port 220 nsew signal input
flabel metal3 s 79200 1368 80000 1488 0 FreeSans 480 0 0 0 wbs_sel_i[2]
port 221 nsew signal input
flabel metal3 s 79200 2048 80000 2168 0 FreeSans 480 0 0 0 wbs_sel_i[3]
port 222 nsew signal input
flabel metal3 s 79200 4088 80000 4208 0 FreeSans 480 0 0 0 wbs_stb_i
port 223 nsew signal input
flabel metal3 s 79200 4768 80000 4888 0 FreeSans 480 0 0 0 wbs_we_i
port 224 nsew signal input
rlabel metal1 39974 37536 39974 37536 0 vccd1
rlabel metal1 39974 36992 39974 36992 0 vssd1
rlabel metal2 15594 12036 15594 12036 0 _0000_
rlabel metal2 21206 11152 21206 11152 0 _0001_
rlabel metal1 55982 2312 55982 2312 0 _0002_
rlabel metal1 34638 29818 34638 29818 0 _0003_
rlabel metal1 47748 32810 47748 32810 0 _0004_
rlabel metal1 48024 33082 48024 33082 0 _0005_
rlabel metal1 45908 35734 45908 35734 0 _0006_
rlabel metal2 43562 36516 43562 36516 0 _0007_
rlabel metal1 42780 34646 42780 34646 0 _0008_
rlabel metal1 36340 29682 36340 29682 0 _0009_
rlabel metal1 37950 31246 37950 31246 0 _0010_
rlabel metal1 40756 30294 40756 30294 0 _0011_
rlabel metal1 41860 35802 41860 35802 0 _0012_
rlabel metal1 42366 32776 42366 32776 0 _0013_
rlabel metal2 39514 34272 39514 34272 0 _0014_
rlabel metal2 37766 33116 37766 33116 0 _0015_
rlabel metal2 45310 30872 45310 30872 0 _0016_
rlabel metal2 47242 30940 47242 30940 0 _0017_
rlabel metal1 55476 2550 55476 2550 0 _0018_
rlabel metal1 56442 2958 56442 2958 0 _0019_
rlabel metal1 19458 10574 19458 10574 0 _0020_
rlabel metal1 20838 12070 20838 12070 0 _0021_
rlabel metal2 36478 16796 36478 16796 0 _0022_
rlabel metal2 44298 10846 44298 10846 0 _0023_
rlabel metal2 47702 12002 47702 12002 0 _0024_
rlabel metal1 46230 14042 46230 14042 0 _0025_
rlabel metal2 33810 9367 33810 9367 0 _0026_
rlabel metal1 30222 20978 30222 20978 0 _0027_
rlabel metal1 48530 20026 48530 20026 0 _0028_
rlabel metal1 31556 14042 31556 14042 0 _0029_
rlabel metal1 38686 17102 38686 17102 0 _0030_
rlabel metal1 42044 9962 42044 9962 0 _0031_
rlabel metal2 47978 10404 47978 10404 0 _0032_
rlabel metal1 48300 13974 48300 13974 0 _0033_
rlabel metal1 31326 9690 31326 9690 0 _0034_
rlabel metal1 28980 22542 28980 22542 0 _0035_
rlabel metal2 50830 20638 50830 20638 0 _0036_
rlabel metal2 33534 15130 33534 15130 0 _0037_
rlabel metal2 41354 16796 41354 16796 0 _0038_
rlabel metal1 40526 9690 40526 9690 0 _0039_
rlabel metal2 48530 8092 48530 8092 0 _0040_
rlabel metal2 50186 13668 50186 13668 0 _0041_
rlabel metal1 32982 8602 32982 8602 0 _0042_
rlabel metal1 32292 22406 32292 22406 0 _0043_
rlabel metal2 53038 20638 53038 20638 0 _0044_
rlabel metal1 35512 15062 35512 15062 0 _0045_
rlabel metal1 43148 17306 43148 17306 0 _0046_
rlabel metal2 40158 8092 40158 8092 0 _0047_
rlabel metal2 49726 6494 49726 6494 0 _0048_
rlabel metal1 52072 13906 52072 13906 0 _0049_
rlabel metal1 29716 8058 29716 8058 0 _0050_
rlabel metal1 30636 23290 30636 23290 0 _0051_
rlabel metal1 56120 19890 56120 19890 0 _0052_
rlabel metal1 37812 15062 37812 15062 0 _0053_
rlabel metal2 42918 17884 42918 17884 0 _0054_
rlabel metal1 43148 6426 43148 6426 0 _0055_
rlabel metal2 49542 4896 49542 4896 0 _0056_
rlabel metal1 53912 13498 53912 13498 0 _0057_
rlabel metal1 30445 6970 30445 6970 0 _0058_
rlabel metal1 29624 24718 29624 24718 0 _0059_
rlabel metal2 56626 21284 56626 21284 0 _0060_
rlabel metal1 40204 15130 40204 15130 0 _0061_
rlabel metal1 39928 20570 39928 20570 0 _0062_
rlabel metal2 41630 6494 41630 6494 0 _0063_
rlabel metal2 51750 5372 51750 5372 0 _0064_
rlabel metal1 55200 15062 55200 15062 0 _0065_
rlabel metal1 30820 5338 30820 5338 0 _0066_
rlabel metal2 30590 26010 30590 26010 0 _0067_
rlabel metal2 53038 22814 53038 22814 0 _0068_
rlabel metal1 42320 15130 42320 15130 0 _0069_
rlabel metal1 39744 21114 39744 21114 0 _0070_
rlabel metal1 40342 4250 40342 4250 0 _0071_
rlabel metal1 53498 4794 53498 4794 0 _0072_
rlabel metal1 52716 16218 52716 16218 0 _0073_
rlabel metal2 35098 6494 35098 6494 0 _0074_
rlabel metal1 32614 26554 32614 26554 0 _0075_
rlabel metal2 55430 22814 55430 22814 0 _0076_
rlabel metal2 44114 14382 44114 14382 0 _0077_
rlabel metal1 36984 20366 36984 20366 0 _0078_
rlabel metal2 41446 3672 41446 3672 0 _0079_
rlabel metal1 55154 7446 55154 7446 0 _0080_
rlabel metal1 54648 16150 54648 16150 0 _0081_
rlabel via1 34092 6970 34092 6970 0 _0082_
rlabel metal1 33258 23290 33258 23290 0 _0083_
rlabel metal1 55660 24922 55660 24922 0 _0084_
rlabel metal1 45356 12410 45356 12410 0 _0085_
rlabel metal2 34730 21012 34730 21012 0 _0086_
rlabel metal1 43240 4250 43240 4250 0 _0087_
rlabel metal1 53360 7786 53360 7786 0 _0088_
rlabel metal2 56166 18462 56166 18462 0 _0089_
rlabel metal2 32338 4828 32338 4828 0 _0090_
rlabel metal2 33810 24956 33810 24956 0 _0091_
rlabel metal1 53268 24854 53268 24854 0 _0092_
rlabel metal2 43010 13022 43010 13022 0 _0093_
rlabel metal1 32890 20026 32890 20026 0 _0094_
rlabel metal2 45310 3740 45310 3740 0 _0095_
rlabel metal2 51566 7650 51566 7650 0 _0096_
rlabel metal1 54142 18394 54142 18394 0 _0097_
rlabel metal1 35558 4046 35558 4046 0 _0098_
rlabel metal1 33580 27642 33580 27642 0 _0099_
rlabel metal2 51106 24616 51106 24616 0 _0100_
rlabel metal1 40572 12614 40572 12614 0 _0101_
rlabel metal2 33902 18462 33902 18462 0 _0102_
rlabel metal2 49082 4250 49082 4250 0 _0103_
rlabel metal1 52900 9690 52900 9690 0 _0104_
rlabel metal1 50784 18394 50784 18394 0 _0105_
rlabel metal1 35926 2958 35926 2958 0 _0106_
rlabel metal1 35282 27642 35282 27642 0 _0107_
rlabel metal1 54142 26554 54142 26554 0 _0108_
rlabel metal2 38226 11356 38226 11356 0 _0109_
rlabel metal1 34224 16150 34224 16150 0 _0110_
rlabel metal2 46506 5916 46506 5916 0 _0111_
rlabel metal1 55660 9690 55660 9690 0 _0112_
rlabel metal2 48346 18462 48346 18462 0 _0113_
rlabel metal2 37214 4828 37214 4828 0 _0114_
rlabel metal1 36708 27642 36708 27642 0 _0115_
rlabel metal2 51152 26350 51152 26350 0 _0116_
rlabel metal1 36156 10778 36156 10778 0 _0117_
rlabel metal1 32016 16218 32016 16218 0 _0118_
rlabel metal2 49082 6494 49082 6494 0 _0119_
rlabel metal2 54510 11492 54510 11492 0 _0120_
rlabel metal1 45724 17850 45724 17850 0 _0121_
rlabel metal2 38134 5916 38134 5916 0 _0122_
rlabel metal2 38134 27268 38134 27268 0 _0123_
rlabel metal2 49174 26724 49174 26724 0 _0124_
rlabel metal2 34730 13022 34730 13022 0 _0125_
rlabel metal2 32154 17884 32154 17884 0 _0126_
rlabel metal1 45632 9690 45632 9690 0 _0127_
rlabel metal2 52670 11628 52670 11628 0 _0128_
rlabel metal1 44206 16626 44206 16626 0 _0129_
rlabel metal1 38088 9146 38088 9146 0 _0130_
rlabel metal2 38226 25092 38226 25092 0 _0131_
rlabel metal2 48438 24548 48438 24548 0 _0132_
rlabel metal2 33994 11934 33994 11934 0 _0133_
rlabel metal2 31142 19108 31142 19108 0 _0134_
rlabel metal1 47242 8058 47242 8058 0 _0135_
rlabel metal2 50738 12002 50738 12002 0 _0136_
rlabel metal1 47058 16626 47058 16626 0 _0137_
rlabel metal2 38778 7514 38778 7514 0 _0138_
rlabel metal1 36294 24922 36294 24922 0 _0139_
rlabel metal1 47840 23154 47840 23154 0 _0140_
rlabel metal1 31464 12274 31464 12274 0 _0141_
rlabel metal1 20884 14246 20884 14246 0 _0142_
rlabel metal1 18308 18938 18308 18938 0 _0143_
rlabel metal2 49266 28764 49266 28764 0 _0144_
rlabel metal1 48438 26010 48438 26010 0 _0145_
rlabel metal2 42642 29410 42642 29410 0 _0146_
rlabel metal2 40158 28764 40158 28764 0 _0147_
rlabel metal2 40434 26724 40434 26724 0 _0148_
rlabel metal1 45862 23834 45862 23834 0 _0149_
rlabel metal1 17894 16082 17894 16082 0 _0150_
rlabel metal2 12466 17306 12466 17306 0 _0151_
rlabel metal2 11822 15844 11822 15844 0 _0152_
rlabel metal1 14950 17306 14950 17306 0 _0153_
rlabel metal2 14306 15844 14306 15844 0 _0154_
rlabel metal1 15502 14042 15502 14042 0 _0155_
rlabel metal1 13248 12614 13248 12614 0 _0156_
rlabel metal2 11822 14110 11822 14110 0 _0157_
rlabel metal1 21666 18360 21666 18360 0 _0158_
rlabel metal1 36478 33898 36478 33898 0 _0159_
rlabel metal1 38640 36346 38640 36346 0 _0160_
rlabel metal1 36110 36278 36110 36278 0 _0161_
rlabel metal1 34592 36346 34592 36346 0 _0162_
rlabel metal1 34171 34374 34171 34374 0 _0163_
rlabel metal2 34730 32164 34730 32164 0 _0164_
rlabel metal1 33856 33082 33856 33082 0 _0165_
rlabel metal2 31510 35292 31510 35292 0 _0166_
rlabel metal2 33534 36380 33534 36380 0 _0167_
rlabel metal2 30406 33762 30406 33762 0 _0168_
rlabel metal2 28750 34884 28750 34884 0 _0169_
rlabel metal1 27830 33626 27830 33626 0 _0170_
rlabel metal1 27646 31994 27646 31994 0 _0171_
rlabel metal2 27646 30940 27646 30940 0 _0172_
rlabel via1 31424 31994 31424 31994 0 _0173_
rlabel metal2 30130 29410 30130 29410 0 _0174_
rlabel metal1 32798 29070 32798 29070 0 _0175_
rlabel metal1 32936 30022 32936 30022 0 _0176_
rlabel metal1 55798 3128 55798 3128 0 _0177_
rlabel metal1 24978 18394 24978 18394 0 _0178_
rlabel metal1 28428 9622 28428 9622 0 _0179_
rlabel metal2 29762 11492 29762 11492 0 _0180_
rlabel metal1 29716 15402 29716 15402 0 _0181_
rlabel metal1 27002 9010 27002 9010 0 _0182_
rlabel metal1 26956 19210 26956 19210 0 _0183_
rlabel metal2 28382 19108 28382 19108 0 _0184_
rlabel metal1 29900 13498 29900 13498 0 _0185_
rlabel metal2 43102 30498 43102 30498 0 _0186_
rlabel metal2 7590 21250 7590 21250 0 _0187_
rlabel metal1 7820 20502 7820 20502 0 _0188_
rlabel metal2 7314 18904 7314 18904 0 _0189_
rlabel metal2 10442 19992 10442 19992 0 _0190_
rlabel metal2 38318 28934 38318 28934 0 _0191_
rlabel metal1 43976 2618 43976 2618 0 _0192_
rlabel via1 50834 3094 50834 3094 0 _0193_
rlabel metal1 56610 16490 56610 16490 0 _0194_
rlabel metal1 38451 3026 38451 3026 0 _0195_
rlabel metal1 39774 23766 39774 23766 0 _0196_
rlabel metal2 56902 22882 56902 22882 0 _0197_
rlabel metal1 40020 2618 40020 2618 0 _0198_
rlabel metal1 45540 21522 45540 21522 0 _0199_
rlabel metal2 43930 24548 43930 24548 0 _0200_
rlabel metal1 46552 26010 46552 26010 0 _0201_
rlabel metal1 42642 25908 42642 25908 0 _0202_
rlabel metal1 42780 25874 42780 25874 0 _0203_
rlabel metal1 43010 26010 43010 26010 0 _0204_
rlabel metal2 43654 26894 43654 26894 0 _0205_
rlabel metal2 43286 27098 43286 27098 0 _0206_
rlabel metal1 43654 26996 43654 26996 0 _0207_
rlabel metal2 42780 24786 42780 24786 0 _0208_
rlabel metal1 41860 29138 41860 29138 0 _0209_
rlabel metal1 42274 23290 42274 23290 0 _0210_
rlabel metal1 44620 26962 44620 26962 0 _0211_
rlabel metal2 40250 22882 40250 22882 0 _0212_
rlabel metal2 40894 26112 40894 26112 0 _0213_
rlabel metal1 44574 24786 44574 24786 0 _0214_
rlabel metal1 47334 21930 47334 21930 0 _0215_
rlabel metal2 21114 15164 21114 15164 0 _0216_
rlabel metal2 21482 17986 21482 17986 0 _0217_
rlabel metal2 39238 36244 39238 36244 0 _0218_
rlabel metal1 36892 35530 36892 35530 0 _0219_
rlabel metal1 35006 36108 35006 36108 0 _0220_
rlabel metal2 36294 34850 36294 34850 0 _0221_
rlabel metal1 35144 31790 35144 31790 0 _0222_
rlabel metal1 34224 33830 34224 33830 0 _0223_
rlabel metal1 33028 35802 33028 35802 0 _0224_
rlabel metal1 31970 35666 31970 35666 0 _0225_
rlabel metal1 28750 33966 28750 33966 0 _0226_
rlabel metal2 31970 33864 31970 33864 0 _0227_
rlabel metal1 28290 33524 28290 33524 0 _0228_
rlabel metal2 28474 33796 28474 33796 0 _0229_
rlabel metal1 27784 31790 27784 31790 0 _0230_
rlabel metal2 28014 32266 28014 32266 0 _0231_
rlabel metal1 30498 31178 30498 31178 0 _0232_
rlabel metal2 30406 32164 30406 32164 0 _0233_
rlabel metal1 31694 29104 31694 29104 0 _0234_
rlabel metal1 29808 29138 29808 29138 0 _0235_
rlabel metal1 31970 30158 31970 30158 0 _0236_
rlabel metal2 20838 16592 20838 16592 0 _0237_
rlabel metal2 25530 15402 25530 15402 0 _0238_
rlabel metal2 23322 14620 23322 14620 0 _0239_
rlabel metal2 20746 16252 20746 16252 0 _0240_
rlabel metal1 25208 15674 25208 15674 0 _0241_
rlabel metal2 22770 14348 22770 14348 0 _0242_
rlabel metal1 22816 14586 22816 14586 0 _0243_
rlabel metal2 24150 15844 24150 15844 0 _0244_
rlabel metal1 26266 15028 26266 15028 0 _0245_
rlabel metal1 22540 13906 22540 13906 0 _0246_
rlabel metal1 26404 15130 26404 15130 0 _0247_
rlabel metal2 24334 11968 24334 11968 0 _0248_
rlabel metal2 26818 13532 26818 13532 0 _0249_
rlabel metal1 26818 15504 26818 15504 0 _0250_
rlabel metal2 27462 13702 27462 13702 0 _0251_
rlabel via1 24888 13906 24888 13906 0 _0252_
rlabel metal1 27416 16490 27416 16490 0 _0253_
rlabel metal1 28106 17204 28106 17204 0 _0254_
rlabel metal1 23966 16422 23966 16422 0 _0255_
rlabel metal2 25622 14382 25622 14382 0 _0256_
rlabel metal2 25622 16252 25622 16252 0 _0257_
rlabel metal2 21114 15725 21114 15725 0 _0258_
rlabel metal1 27968 16490 27968 16490 0 _0259_
rlabel metal1 27600 17102 27600 17102 0 _0260_
rlabel metal1 27968 13226 27968 13226 0 _0261_
rlabel metal1 25622 15946 25622 15946 0 _0262_
rlabel via1 29026 16082 29026 16082 0 _0263_
rlabel metal1 30130 13260 30130 13260 0 _0264_
rlabel metal1 25668 17782 25668 17782 0 _0265_
rlabel metal1 26726 15878 26726 15878 0 _0266_
rlabel metal1 24518 11662 24518 11662 0 _0267_
rlabel metal2 24794 16422 24794 16422 0 _0268_
rlabel metal1 23644 11526 23644 11526 0 _0269_
rlabel metal1 23460 11322 23460 11322 0 _0270_
rlabel metal2 23322 11900 23322 11900 0 _0271_
rlabel metal1 25162 18122 25162 18122 0 _0272_
rlabel metal1 26036 16694 26036 16694 0 _0273_
rlabel metal1 25484 16762 25484 16762 0 _0274_
rlabel metal1 29164 10574 29164 10574 0 _0275_
rlabel metal1 23138 13906 23138 13906 0 _0276_
rlabel via1 24152 13906 24152 13906 0 _0277_
rlabel metal2 23966 13430 23966 13430 0 _0278_
rlabel metal1 28566 12172 28566 12172 0 _0279_
rlabel metal1 24426 13872 24426 13872 0 _0280_
rlabel metal1 25254 13906 25254 13906 0 _0281_
rlabel metal1 25346 12818 25346 12818 0 _0282_
rlabel metal2 25714 13294 25714 13294 0 _0283_
rlabel metal1 27922 13294 27922 13294 0 _0284_
rlabel metal1 25760 12410 25760 12410 0 _0285_
rlabel metal2 27922 11628 27922 11628 0 _0286_
rlabel metal2 27830 12274 27830 12274 0 _0287_
rlabel metal1 26312 12614 26312 12614 0 _0288_
rlabel metal1 28474 10574 28474 10574 0 _0289_
rlabel metal1 29026 15504 29026 15504 0 _0290_
rlabel metal2 28658 10812 28658 10812 0 _0291_
rlabel metal2 23230 14042 23230 14042 0 _0292_
rlabel metal1 22678 14042 22678 14042 0 _0293_
rlabel metal2 23690 14076 23690 14076 0 _0294_
rlabel metal1 25300 14246 25300 14246 0 _0295_
rlabel metal1 27646 13838 27646 13838 0 _0296_
rlabel metal2 26450 11322 26450 11322 0 _0297_
rlabel metal1 26496 11322 26496 11322 0 _0298_
rlabel metal1 29394 11050 29394 11050 0 _0299_
rlabel metal1 27784 13702 27784 13702 0 _0300_
rlabel metal2 28106 14076 28106 14076 0 _0301_
rlabel metal1 27922 14008 27922 14008 0 _0302_
rlabel metal1 28612 14042 28612 14042 0 _0303_
rlabel metal2 27830 14348 27830 14348 0 _0304_
rlabel metal1 27048 13362 27048 13362 0 _0305_
rlabel metal1 26634 13158 26634 13158 0 _0306_
rlabel metal2 26634 10234 26634 10234 0 _0307_
rlabel via1 27370 18734 27370 18734 0 _0308_
rlabel metal1 26220 16218 26220 16218 0 _0309_
rlabel metal1 25346 18190 25346 18190 0 _0310_
rlabel metal1 27738 17646 27738 17646 0 _0311_
rlabel metal1 26818 17850 26818 17850 0 _0312_
rlabel metal1 26818 18394 26818 18394 0 _0313_
rlabel metal2 28382 18496 28382 18496 0 _0314_
rlabel metal2 30406 13770 30406 13770 0 _0315_
rlabel metal1 43838 24582 43838 24582 0 _0316_
rlabel metal1 40206 23086 40206 23086 0 _0317_
rlabel metal2 46690 20128 46690 20128 0 _0318_
rlabel metal1 48392 22610 48392 22610 0 _0319_
rlabel metal1 44022 20298 44022 20298 0 _0320_
rlabel metal1 45310 21964 45310 21964 0 _0321_
rlabel metal1 41584 25398 41584 25398 0 _0322_
rlabel metal1 41538 25228 41538 25228 0 _0323_
rlabel metal2 48622 15708 48622 15708 0 _0324_
rlabel metal1 44436 22610 44436 22610 0 _0325_
rlabel metal1 40526 13736 40526 13736 0 _0326_
rlabel metal1 42274 25466 42274 25466 0 _0327_
rlabel metal1 10488 20366 10488 20366 0 _0328_
rlabel metal2 9890 20128 9890 20128 0 _0329_
rlabel metal1 7636 20026 7636 20026 0 _0330_
rlabel metal1 7360 20570 7360 20570 0 _0331_
rlabel metal1 7866 20910 7866 20910 0 _0332_
rlabel metal1 7544 19346 7544 19346 0 _0333_
rlabel metal2 10074 20247 10074 20247 0 _0334_
rlabel metal1 47288 19822 47288 19822 0 _0335_
rlabel metal2 51566 23188 51566 23188 0 _0336_
rlabel metal2 38870 19210 38870 19210 0 _0337_
rlabel metal1 36984 18054 36984 18054 0 _0338_
rlabel metal1 37950 22066 37950 22066 0 _0339_
rlabel metal1 38226 18122 38226 18122 0 _0340_
rlabel metal1 38090 19346 38090 19346 0 _0341_
rlabel metal1 36662 13906 36662 13906 0 _0342_
rlabel metal2 38318 21454 38318 21454 0 _0343_
rlabel metal1 36754 18666 36754 18666 0 _0344_
rlabel metal1 36754 20026 36754 20026 0 _0345_
rlabel metal1 39491 18734 39491 18734 0 _0346_
rlabel via2 36662 14365 36662 14365 0 _0347_
rlabel via2 36754 19363 36754 19363 0 _0348_
rlabel metal2 37674 18785 37674 18785 0 _0349_
rlabel metal1 37950 6698 37950 6698 0 _0350_
rlabel metal1 36892 19686 36892 19686 0 _0351_
rlabel metal1 40388 22950 40388 22950 0 _0352_
rlabel metal1 36248 18394 36248 18394 0 _0353_
rlabel metal1 37582 19414 37582 19414 0 _0354_
rlabel metal1 37306 18734 37306 18734 0 _0355_
rlabel metal2 40158 19040 40158 19040 0 _0356_
rlabel metal1 38410 18700 38410 18700 0 _0357_
rlabel metal2 38226 19040 38226 19040 0 _0358_
rlabel metal1 38226 18836 38226 18836 0 _0359_
rlabel metal1 40250 18700 40250 18700 0 _0360_
rlabel metal1 38226 18734 38226 18734 0 _0361_
rlabel metal1 39008 28526 39008 28526 0 _0362_
rlabel metal2 46598 10880 46598 10880 0 _0363_
rlabel metal1 44666 8364 44666 8364 0 _0364_
rlabel metal2 42642 8262 42642 8262 0 _0365_
rlabel metal1 44252 7514 44252 7514 0 _0366_
rlabel metal1 43746 8466 43746 8466 0 _0367_
rlabel metal1 43654 8296 43654 8296 0 _0368_
rlabel metal2 43746 8313 43746 8313 0 _0369_
rlabel metal1 43792 9554 43792 9554 0 _0370_
rlabel metal1 43838 8534 43838 8534 0 _0371_
rlabel metal2 43102 2587 43102 2587 0 _0372_
rlabel metal1 50278 9146 50278 9146 0 _0373_
rlabel metal1 49818 11832 49818 11832 0 _0374_
rlabel metal2 51106 10302 51106 10302 0 _0375_
rlabel metal1 50094 8466 50094 8466 0 _0376_
rlabel metal1 50968 8602 50968 8602 0 _0377_
rlabel metal1 50278 9690 50278 9690 0 _0378_
rlabel metal2 51014 9452 51014 9452 0 _0379_
rlabel metal1 51566 9690 51566 9690 0 _0380_
rlabel metal2 51290 9418 51290 9418 0 _0381_
rlabel metal2 51382 6256 51382 6256 0 _0382_
rlabel metal1 50784 2618 50784 2618 0 _0383_
rlabel metal2 39698 10591 39698 10591 0 _0384_
rlabel metal1 48668 15878 48668 15878 0 _0385_
rlabel metal1 50232 16082 50232 16082 0 _0386_
rlabel metal1 50094 16558 50094 16558 0 _0387_
rlabel metal2 50002 16320 50002 16320 0 _0388_
rlabel metal2 51198 15878 51198 15878 0 _0389_
rlabel viali 51101 16082 51101 16082 0 _0390_
rlabel metal1 50094 15946 50094 15946 0 _0391_
rlabel metal1 48438 15980 48438 15980 0 _0392_
rlabel metal1 48438 16082 48438 16082 0 _0393_
rlabel metal1 49910 16184 49910 16184 0 _0394_
rlabel metal1 50416 15946 50416 15946 0 _0395_
rlabel metal1 35834 8500 35834 8500 0 _0396_
rlabel metal1 36432 6630 36432 6630 0 _0397_
rlabel metal2 35466 8194 35466 8194 0 _0398_
rlabel metal2 37582 8534 37582 8534 0 _0399_
rlabel metal1 37030 8262 37030 8262 0 _0400_
rlabel metal1 36984 8466 36984 8466 0 _0401_
rlabel metal1 37996 9894 37996 9894 0 _0402_
rlabel metal2 37306 8806 37306 8806 0 _0403_
rlabel metal1 37904 8330 37904 8330 0 _0404_
rlabel metal1 38456 22474 38456 22474 0 _0405_
rlabel metal1 36110 23766 36110 23766 0 _0406_
rlabel metal1 36662 22508 36662 22508 0 _0407_
rlabel metal1 39376 22474 39376 22474 0 _0408_
rlabel metal2 39146 22916 39146 22916 0 _0409_
rlabel metal1 40434 23290 40434 23290 0 _0410_
rlabel metal2 36754 22950 36754 22950 0 _0411_
rlabel metal1 36386 23120 36386 23120 0 _0412_
rlabel metal1 36294 23154 36294 23154 0 _0413_
rlabel metal2 36570 22780 36570 22780 0 _0414_
rlabel metal1 37168 22474 37168 22474 0 _0415_
rlabel metal2 39146 23868 39146 23868 0 _0416_
rlabel metal1 50600 21522 50600 21522 0 _0417_
rlabel metal2 51106 23290 51106 23290 0 _0418_
rlabel metal2 51566 22780 51566 22780 0 _0419_
rlabel metal1 49772 22202 49772 22202 0 _0420_
rlabel metal1 51290 22440 51290 22440 0 _0421_
rlabel metal1 51336 21658 51336 21658 0 _0422_
rlabel metal1 50554 22644 50554 22644 0 _0423_
rlabel metal1 51290 22712 51290 22712 0 _0424_
rlabel metal1 56258 22678 56258 22678 0 _0425_
rlabel metal1 37076 12954 37076 12954 0 _0426_
rlabel metal1 36892 13498 36892 13498 0 _0427_
rlabel metal1 39698 13328 39698 13328 0 _0428_
rlabel metal2 37858 13124 37858 13124 0 _0429_
rlabel metal1 39155 13430 39155 13430 0 _0430_
rlabel metal1 40618 13804 40618 13804 0 _0431_
rlabel metal2 40434 13600 40434 13600 0 _0432_
rlabel metal2 39422 13600 39422 13600 0 _0433_
rlabel metal1 37030 13430 37030 13430 0 _0434_
rlabel metal1 38410 13362 38410 13362 0 _0435_
rlabel metal1 40434 2482 40434 2482 0 _0436_
rlabel metal1 48162 28050 48162 28050 0 _0437_
rlabel metal1 43148 28526 43148 28526 0 _0438_
rlabel metal2 45954 27064 45954 27064 0 _0439_
rlabel metal2 46046 27472 46046 27472 0 _0440_
rlabel metal2 21482 14212 21482 14212 0 _0441_
rlabel metal1 17618 25228 17618 25228 0 _0442_
rlabel metal1 34040 32742 34040 32742 0 _0443_
rlabel metal1 40250 31280 40250 31280 0 _0444_
rlabel metal1 64860 3128 64860 3128 0 _0445_
rlabel metal1 59938 2856 59938 2856 0 _0446_
rlabel metal2 55062 2176 55062 2176 0 _0447_
rlabel metal1 59662 3094 59662 3094 0 _0448_
rlabel metal2 68494 3196 68494 3196 0 _0449_
rlabel metal2 72634 3434 72634 3434 0 _0450_
rlabel metal1 74520 2958 74520 2958 0 _0451_
rlabel metal2 72266 2788 72266 2788 0 _0452_
rlabel metal1 71576 3094 71576 3094 0 _0453_
rlabel metal2 72542 3298 72542 3298 0 _0454_
rlabel metal1 58558 3536 58558 3536 0 _0455_
rlabel metal2 58466 3162 58466 3162 0 _0456_
rlabel via1 22126 16626 22126 16626 0 _0457_
rlabel metal2 20378 17238 20378 17238 0 _0458_
rlabel metal2 28750 14042 28750 14042 0 _0459_
rlabel metal2 19734 13889 19734 13889 0 _0460_
rlabel metal1 17871 11798 17871 11798 0 _0461_
rlabel metal1 19964 12410 19964 12410 0 _0462_
rlabel metal1 19550 12716 19550 12716 0 _0463_
rlabel metal2 14122 15640 14122 15640 0 _0464_
rlabel metal2 16146 15810 16146 15810 0 _0465_
rlabel metal2 17066 16592 17066 16592 0 _0466_
rlabel metal2 14306 14586 14306 14586 0 _0467_
rlabel metal1 14444 14382 14444 14382 0 _0468_
rlabel metal1 14766 12954 14766 12954 0 _0469_
rlabel metal1 17204 15130 17204 15130 0 _0470_
rlabel metal1 17894 16150 17894 16150 0 _0471_
rlabel metal1 17618 13906 17618 13906 0 _0472_
rlabel metal2 17986 14246 17986 14246 0 _0473_
rlabel metal1 18124 12206 18124 12206 0 _0474_
rlabel metal2 19090 12988 19090 12988 0 _0475_
rlabel metal2 17434 11934 17434 11934 0 _0476_
rlabel metal1 18124 11866 18124 11866 0 _0477_
rlabel metal1 17112 11730 17112 11730 0 _0478_
rlabel metal1 20838 12784 20838 12784 0 _0479_
rlabel metal1 9752 18258 9752 18258 0 _0480_
rlabel metal1 15502 25840 15502 25840 0 _0481_
rlabel metal1 16330 25738 16330 25738 0 _0482_
rlabel metal1 15318 29716 15318 29716 0 _0483_
rlabel metal1 15640 30022 15640 30022 0 _0484_
rlabel metal1 14214 25364 14214 25364 0 _0485_
rlabel metal2 13202 24922 13202 24922 0 _0486_
rlabel metal2 14582 25568 14582 25568 0 _0487_
rlabel metal2 14582 29104 14582 29104 0 _0488_
rlabel metal2 13386 28900 13386 28900 0 _0489_
rlabel metal2 15134 27166 15134 27166 0 _0490_
rlabel metal1 11362 20944 11362 20944 0 _0491_
rlabel metal1 15180 24582 15180 24582 0 _0492_
rlabel metal2 14490 24956 14490 24956 0 _0493_
rlabel metal1 12374 24752 12374 24752 0 _0494_
rlabel metal1 13064 24242 13064 24242 0 _0495_
rlabel metal1 10350 24378 10350 24378 0 _0496_
rlabel metal2 10626 23970 10626 23970 0 _0497_
rlabel metal1 12558 27030 12558 27030 0 _0498_
rlabel metal2 12466 27234 12466 27234 0 _0499_
rlabel metal1 10350 26792 10350 26792 0 _0500_
rlabel metal2 10994 26996 10994 26996 0 _0501_
rlabel metal1 10718 27642 10718 27642 0 _0502_
rlabel metal1 10526 27098 10526 27098 0 _0503_
rlabel metal1 10764 28730 10764 28730 0 _0504_
rlabel metal1 10718 28084 10718 28084 0 _0505_
rlabel metal1 12604 30294 12604 30294 0 _0506_
rlabel metal1 10994 29172 10994 29172 0 _0507_
rlabel metal1 13018 30192 13018 30192 0 _0508_
rlabel metal1 10994 30736 10994 30736 0 _0509_
rlabel metal2 13340 30226 13340 30226 0 _0510_
rlabel metal1 13435 30226 13435 30226 0 _0511_
rlabel metal1 16008 28730 16008 28730 0 _0512_
rlabel metal1 15916 28526 15916 28526 0 _0513_
rlabel metal1 15932 28458 15932 28458 0 _0514_
rlabel metal2 15686 28492 15686 28492 0 _0515_
rlabel metal1 15456 30906 15456 30906 0 _0516_
rlabel metal1 16698 31824 16698 31824 0 _0517_
rlabel metal1 17618 30804 17618 30804 0 _0518_
rlabel via1 17720 29546 17720 29546 0 _0519_
rlabel metal2 18446 30022 18446 30022 0 _0520_
rlabel metal2 19274 29818 19274 29818 0 _0521_
rlabel metal1 19274 29512 19274 29512 0 _0522_
rlabel metal2 20470 27812 20470 27812 0 _0523_
rlabel metal2 20654 27812 20654 27812 0 _0524_
rlabel metal2 19458 27642 19458 27642 0 _0525_
rlabel metal2 19090 25466 19090 25466 0 _0526_
rlabel metal2 16974 23324 16974 23324 0 _0527_
rlabel metal2 17250 23868 17250 23868 0 _0528_
rlabel metal1 17296 22066 17296 22066 0 _0529_
rlabel metal1 17526 24922 17526 24922 0 _0530_
rlabel metal1 17158 24684 17158 24684 0 _0531_
rlabel metal1 31786 30838 31786 30838 0 _0532_
rlabel metal2 30314 32810 30314 32810 0 _0533_
rlabel metal2 32062 33082 32062 33082 0 _0534_
rlabel metal1 35619 32878 35619 32878 0 _0535_
rlabel metal1 38778 35802 38778 35802 0 _0536_
rlabel metal1 35926 36686 35926 36686 0 _0537_
rlabel metal1 35650 35802 35650 35802 0 _0538_
rlabel metal2 35466 32742 35466 32742 0 _0539_
rlabel metal1 36800 33490 36800 33490 0 _0540_
rlabel metal2 41446 33133 41446 33133 0 _0541_
rlabel metal1 36202 30022 36202 30022 0 _0542_
rlabel metal1 36494 30294 36494 30294 0 _0543_
rlabel metal1 37122 30906 37122 30906 0 _0544_
rlabel metal1 37628 30906 37628 30906 0 _0545_
rlabel metal1 40710 31144 40710 31144 0 _0546_
rlabel metal1 40702 33626 40702 33626 0 _0547_
rlabel via1 40718 31450 40718 31450 0 _0548_
rlabel metal1 41400 35462 41400 35462 0 _0549_
rlabel metal1 41178 35802 41178 35802 0 _0550_
rlabel metal1 44666 32912 44666 32912 0 _0551_
rlabel metal2 44482 32572 44482 32572 0 _0552_
rlabel metal1 44160 32402 44160 32402 0 _0553_
rlabel metal2 43838 33354 43838 33354 0 _0554_
rlabel metal1 44114 32980 44114 32980 0 _0555_
rlabel metal2 56074 23120 56074 23120 0 _0556_
rlabel metal1 44482 31926 44482 31926 0 _0557_
rlabel metal2 48070 32266 48070 32266 0 _0558_
rlabel metal1 39682 33558 39682 33558 0 _0559_
rlabel metal2 41170 33728 41170 33728 0 _0560_
rlabel metal1 39606 33898 39606 33898 0 _0561_
rlabel metal2 38962 33524 38962 33524 0 _0562_
rlabel via1 46590 32742 46590 32742 0 _0563_
rlabel metal1 37766 33082 37766 33082 0 _0564_
rlabel metal1 45264 31382 45264 31382 0 _0565_
rlabel metal1 45678 31382 45678 31382 0 _0566_
rlabel metal1 48024 32402 48024 32402 0 _0567_
rlabel metal1 46920 31314 46920 31314 0 _0568_
rlabel metal2 47610 32708 47610 32708 0 _0569_
rlabel metal1 47656 32470 47656 32470 0 _0570_
rlabel metal1 46322 32538 46322 32538 0 _0571_
rlabel metal1 46046 36210 46046 36210 0 _0572_
rlabel metal2 47518 33082 47518 33082 0 _0573_
rlabel metal1 46000 35258 46000 35258 0 _0574_
rlabel metal1 44022 36006 44022 36006 0 _0575_
rlabel metal2 43562 34510 43562 34510 0 _0576_
rlabel metal2 43378 34612 43378 34612 0 _0577_
rlabel metal1 42918 33388 42918 33388 0 _0578_
rlabel metal2 46138 34102 46138 34102 0 _0579_
rlabel metal1 18630 12852 18630 12852 0 _0580_
rlabel metal1 21206 12240 21206 12240 0 _0581_
rlabel metal2 20378 15266 20378 15266 0 _0582_
rlabel metal1 27991 14994 27991 14994 0 _0583_
rlabel metal1 20976 16082 20976 16082 0 _0584_
rlabel metal1 26450 17306 26450 17306 0 _0585_
rlabel metal1 33718 4624 33718 4624 0 _0586_
rlabel metal1 28336 17170 28336 17170 0 _0587_
rlabel via2 33626 17187 33626 17187 0 _0588_
rlabel metal2 31050 17442 31050 17442 0 _0589_
rlabel metal1 29164 14994 29164 14994 0 _0590_
rlabel metal2 28198 17510 28198 17510 0 _0591_
rlabel metal1 32706 17544 32706 17544 0 _0592_
rlabel metal1 36754 17204 36754 17204 0 _0593_
rlabel metal1 44068 10778 44068 10778 0 _0594_
rlabel metal2 47978 11798 47978 11798 0 _0595_
rlabel metal1 46690 13940 46690 13940 0 _0596_
rlabel metal1 34960 10098 34960 10098 0 _0597_
rlabel metal2 34270 23834 34270 23834 0 _0598_
rlabel metal1 30774 21420 30774 21420 0 _0599_
rlabel metal2 48898 20298 48898 20298 0 _0600_
rlabel metal1 32246 13974 32246 13974 0 _0601_
rlabel metal2 38410 16966 38410 16966 0 _0602_
rlabel metal2 42090 10948 42090 10948 0 _0603_
rlabel metal1 48254 10098 48254 10098 0 _0604_
rlabel metal1 48484 14382 48484 14382 0 _0605_
rlabel metal2 31878 9350 31878 9350 0 _0606_
rlabel metal1 29900 21998 29900 21998 0 _0607_
rlabel metal2 50922 20468 50922 20468 0 _0608_
rlabel metal1 33764 13702 33764 13702 0 _0609_
rlabel metal2 41354 17340 41354 17340 0 _0610_
rlabel metal1 41078 9486 41078 9486 0 _0611_
rlabel metal2 48898 8908 48898 8908 0 _0612_
rlabel metal1 50462 13328 50462 13328 0 _0613_
rlabel metal1 32890 8466 32890 8466 0 _0614_
rlabel metal1 32430 22644 32430 22644 0 _0615_
rlabel metal2 52854 20434 52854 20434 0 _0616_
rlabel metal1 35466 14586 35466 14586 0 _0617_
rlabel metal2 43470 17340 43470 17340 0 _0618_
rlabel metal1 40802 8466 40802 8466 0 _0619_
rlabel metal1 49680 6766 49680 6766 0 _0620_
rlabel metal2 52210 14076 52210 14076 0 _0621_
rlabel metal2 30406 8058 30406 8058 0 _0622_
rlabel metal1 31050 23052 31050 23052 0 _0623_
rlabel metal2 55154 20604 55154 20604 0 _0624_
rlabel metal1 37628 14586 37628 14586 0 _0625_
rlabel metal2 42642 18564 42642 18564 0 _0626_
rlabel metal1 43286 6324 43286 6324 0 _0627_
rlabel metal2 49726 5372 49726 5372 0 _0628_
rlabel metal1 54096 13294 54096 13294 0 _0629_
rlabel metal2 31050 7548 31050 7548 0 _0630_
rlabel metal1 30912 24378 30912 24378 0 _0631_
rlabel metal1 56350 20978 56350 20978 0 _0632_
rlabel metal1 40296 14994 40296 14994 0 _0633_
rlabel metal2 40066 19958 40066 19958 0 _0634_
rlabel metal1 42182 6732 42182 6732 0 _0635_
rlabel metal1 52026 5236 52026 5236 0 _0636_
rlabel metal1 55614 15436 55614 15436 0 _0637_
rlabel metal2 31234 5644 31234 5644 0 _0638_
rlabel metal1 30958 25466 30958 25466 0 _0639_
rlabel metal1 53268 22202 53268 22202 0 _0640_
rlabel metal2 42090 14790 42090 14790 0 _0641_
rlabel metal1 39008 20570 39008 20570 0 _0642_
rlabel metal1 40940 4114 40940 4114 0 _0643_
rlabel metal2 53682 5338 53682 5338 0 _0644_
rlabel metal1 52762 16082 52762 16082 0 _0645_
rlabel metal2 35374 6324 35374 6324 0 _0646_
rlabel metal2 32430 26180 32430 26180 0 _0647_
rlabel metal2 55154 23052 55154 23052 0 _0648_
rlabel metal2 44022 14790 44022 14790 0 _0649_
rlabel metal1 36754 20468 36754 20468 0 _0650_
rlabel metal1 41354 4080 41354 4080 0 _0651_
rlabel metal1 54694 7446 54694 7446 0 _0652_
rlabel metal2 54786 16762 54786 16762 0 _0653_
rlabel metal1 33810 6426 33810 6426 0 _0654_
rlabel metal1 33626 23052 33626 23052 0 _0655_
rlabel metal1 55660 24378 55660 24378 0 _0656_
rlabel metal1 45632 13158 45632 13158 0 _0657_
rlabel metal2 35006 20604 35006 20604 0 _0658_
rlabel metal1 43516 4114 43516 4114 0 _0659_
rlabel metal2 53498 7990 53498 7990 0 _0660_
rlabel metal1 54648 17850 54648 17850 0 _0661_
rlabel metal2 33166 5372 33166 5372 0 _0662_
rlabel metal1 34270 25228 34270 25228 0 _0663_
rlabel metal1 53452 24378 53452 24378 0 _0664_
rlabel metal1 42964 13294 42964 13294 0 _0665_
rlabel metal1 33626 19788 33626 19788 0 _0666_
rlabel metal1 45494 4114 45494 4114 0 _0667_
rlabel metal2 51750 7820 51750 7820 0 _0668_
rlabel metal1 53728 17850 53728 17850 0 _0669_
rlabel metal2 35558 4794 35558 4794 0 _0670_
rlabel metal1 34454 26554 34454 26554 0 _0671_
rlabel metal1 51566 24922 51566 24922 0 _0672_
rlabel metal1 40526 11866 40526 11866 0 _0673_
rlabel metal1 34178 18700 34178 18700 0 _0674_
rlabel metal1 47564 4590 47564 4590 0 _0675_
rlabel metal2 53038 9724 53038 9724 0 _0676_
rlabel metal1 51060 18258 51060 18258 0 _0677_
rlabel metal2 36478 4556 36478 4556 0 _0678_
rlabel metal1 35374 27098 35374 27098 0 _0679_
rlabel metal1 53544 26010 53544 26010 0 _0680_
rlabel metal2 38410 11900 38410 11900 0 _0681_
rlabel metal2 34546 17340 34546 17340 0 _0682_
rlabel metal1 46506 6358 46506 6358 0 _0683_
rlabel metal2 55062 9248 55062 9248 0 _0684_
rlabel metal2 48438 18292 48438 18292 0 _0685_
rlabel metal2 37490 5372 37490 5372 0 _0686_
rlabel metal2 36938 27268 36938 27268 0 _0687_
rlabel metal2 51474 26044 51474 26044 0 _0688_
rlabel metal1 36524 10642 36524 10642 0 _0689_
rlabel metal2 32430 16524 32430 16524 0 _0690_
rlabel metal1 47426 6732 47426 6732 0 _0691_
rlabel metal2 54786 10948 54786 10948 0 _0692_
rlabel metal1 46230 17306 46230 17306 0 _0693_
rlabel metal1 38318 6290 38318 6290 0 _0694_
rlabel metal1 38502 26010 38502 26010 0 _0695_
rlabel metal2 49910 26146 49910 26146 0 _0696_
rlabel metal1 35098 13260 35098 13260 0 _0697_
rlabel metal1 32476 18258 32476 18258 0 _0698_
rlabel metal2 45954 8806 45954 8806 0 _0699_
rlabel metal1 52946 11152 52946 11152 0 _0700_
rlabel metal1 46322 15878 46322 15878 0 _0701_
rlabel metal1 38640 8602 38640 8602 0 _0702_
rlabel metal1 38502 24752 38502 24752 0 _0703_
rlabel metal1 48714 24106 48714 24106 0 _0704_
rlabel metal1 33856 12206 33856 12206 0 _0705_
rlabel metal2 32890 19006 32890 19006 0 _0706_
rlabel metal1 47058 7820 47058 7820 0 _0707_
rlabel metal2 51014 11526 51014 11526 0 _0708_
rlabel metal1 46368 16218 46368 16218 0 _0709_
rlabel metal1 38686 7820 38686 7820 0 _0710_
rlabel metal1 36754 24752 36754 24752 0 _0711_
rlabel metal1 48760 23290 48760 23290 0 _0712_
rlabel metal1 31556 12818 31556 12818 0 _0713_
rlabel metal1 20608 15538 20608 15538 0 _0714_
rlabel metal2 20562 15164 20562 15164 0 _0715_
rlabel via1 46125 26282 46125 26282 0 _0716_
rlabel metal1 42780 28662 42780 28662 0 _0717_
rlabel metal2 44574 27438 44574 27438 0 _0718_
rlabel metal1 45954 27914 45954 27914 0 _0719_
rlabel metal1 46552 28118 46552 28118 0 _0720_
rlabel metal1 46046 29104 46046 29104 0 _0721_
rlabel metal2 46506 28730 46506 28730 0 _0722_
rlabel metal1 46368 28526 46368 28526 0 _0723_
rlabel metal1 46644 28662 46644 28662 0 _0724_
rlabel metal1 44643 32810 44643 32810 0 _0725_
rlabel metal1 44896 31790 44896 31790 0 _0726_
rlabel metal1 48438 28186 48438 28186 0 _0727_
rlabel metal2 44850 25330 44850 25330 0 _0728_
rlabel metal2 44114 25534 44114 25534 0 _0729_
rlabel metal1 44244 24922 44244 24922 0 _0730_
rlabel metal2 31786 20162 31786 20162 0 clknet_0_wb_clk_i
rlabel metal1 17342 12138 17342 12138 0 clknet_1_0__leaf_wb_clk_i
rlabel metal2 45126 33694 45126 33694 0 clknet_1_1__leaf_wb_clk_i
rlabel metal2 9522 17986 9522 17986 0 clknet_leaf_0_wb_clk_i
rlabel metal2 34270 30464 34270 30464 0 clknet_leaf_10_wb_clk_i
rlabel metal2 36202 36448 36202 36448 0 clknet_leaf_11_wb_clk_i
rlabel metal2 42274 36448 42274 36448 0 clknet_leaf_12_wb_clk_i
rlabel metal1 55269 25330 55269 25330 0 clknet_leaf_13_wb_clk_i
rlabel metal1 57132 23086 57132 23086 0 clknet_leaf_14_wb_clk_i
rlabel metal1 40066 21556 40066 21556 0 clknet_leaf_15_wb_clk_i
rlabel metal2 38594 19074 38594 19074 0 clknet_leaf_16_wb_clk_i
rlabel metal1 45310 18292 45310 18292 0 clknet_leaf_17_wb_clk_i
rlabel metal1 51704 16626 51704 16626 0 clknet_leaf_18_wb_clk_i
rlabel metal2 51842 11492 51842 11492 0 clknet_leaf_19_wb_clk_i
rlabel metal1 16790 17102 16790 17102 0 clknet_leaf_1_wb_clk_i
rlabel metal1 55890 2482 55890 2482 0 clknet_leaf_20_wb_clk_i
rlabel metal1 49404 6222 49404 6222 0 clknet_leaf_21_wb_clk_i
rlabel metal2 34822 6528 34822 6528 0 clknet_leaf_22_wb_clk_i
rlabel metal2 33626 9792 33626 9792 0 clknet_leaf_23_wb_clk_i
rlabel metal1 30314 12206 30314 12206 0 clknet_leaf_24_wb_clk_i
rlabel metal2 21482 10336 21482 10336 0 clknet_leaf_25_wb_clk_i
rlabel metal1 29670 6834 29670 6834 0 clknet_leaf_26_wb_clk_i
rlabel metal2 17158 11730 17158 11730 0 clknet_leaf_27_wb_clk_i
rlabel metal1 25622 19822 25622 19822 0 clknet_leaf_2_wb_clk_i
rlabel metal1 14260 21454 14260 21454 0 clknet_leaf_3_wb_clk_i
rlabel metal1 7590 21556 7590 21556 0 clknet_leaf_4_wb_clk_i
rlabel metal1 11730 31790 11730 31790 0 clknet_leaf_5_wb_clk_i
rlabel metal1 19596 31858 19596 31858 0 clknet_leaf_6_wb_clk_i
rlabel metal2 30222 34544 30222 34544 0 clknet_leaf_7_wb_clk_i
rlabel metal2 23598 25568 23598 25568 0 clknet_leaf_8_wb_clk_i
rlabel metal1 32108 21998 32108 21998 0 clknet_leaf_9_wb_clk_i
rlabel metal1 1380 16082 1380 16082 0 gpio_in[34]
rlabel metal2 1426 13787 1426 13787 0 gpio_in[35]
rlabel metal1 1334 14382 1334 14382 0 gpio_in[36]
rlabel metal2 1426 15249 1426 15249 0 gpio_in[37]
rlabel metal3 751 22508 751 22508 0 gpio_oeb[0]
rlabel metal3 820 34068 820 34068 0 gpio_oeb[10]
rlabel metal1 1610 26554 1610 26554 0 gpio_oeb[11]
rlabel metal3 820 25228 820 25228 0 gpio_oeb[12]
rlabel metal1 1610 23834 1610 23834 0 gpio_oeb[13]
rlabel metal1 1610 29274 1610 29274 0 gpio_oeb[14]
rlabel metal3 820 33388 820 33388 0 gpio_oeb[15]
rlabel metal1 1610 34714 1610 34714 0 gpio_oeb[16]
rlabel metal3 820 35428 820 35428 0 gpio_oeb[17]
rlabel metal1 40158 36890 40158 36890 0 gpio_oeb[18]
rlabel metal1 73186 36890 73186 36890 0 gpio_oeb[19]
rlabel metal3 820 31348 820 31348 0 gpio_oeb[1]
rlabel metal1 55338 36890 55338 36890 0 gpio_oeb[20]
rlabel metal1 51520 36890 51520 36890 0 gpio_oeb[21]
rlabel metal1 41216 36890 41216 36890 0 gpio_oeb[22]
rlabel metal1 68356 36890 68356 36890 0 gpio_oeb[23]
rlabel metal1 58604 36890 58604 36890 0 gpio_oeb[24]
rlabel metal2 48990 38056 48990 38056 0 gpio_oeb[25]
rlabel metal1 59248 36890 59248 36890 0 gpio_oeb[26]
rlabel metal2 59938 38056 59938 38056 0 gpio_oeb[27]
rlabel metal1 45724 36890 45724 36890 0 gpio_oeb[28]
rlabel metal1 55982 36890 55982 36890 0 gpio_oeb[29]
rlabel metal3 958 23188 958 23188 0 gpio_oeb[2]
rlabel metal1 54050 36890 54050 36890 0 gpio_oeb[30]
rlabel metal1 56672 36890 56672 36890 0 gpio_oeb[31]
rlabel metal1 60536 36890 60536 36890 0 gpio_oeb[32]
rlabel metal1 50876 36890 50876 36890 0 gpio_oeb[33]
rlabel metal3 820 36108 820 36108 0 gpio_oeb[34]
rlabel metal3 820 24548 820 24548 0 gpio_oeb[35]
rlabel metal3 820 27948 820 27948 0 gpio_oeb[36]
rlabel metal1 1840 36346 1840 36346 0 gpio_oeb[37]
rlabel metal3 820 25908 820 25908 0 gpio_oeb[3]
rlabel metal3 820 27268 820 27268 0 gpio_oeb[4]
rlabel metal3 820 29988 820 29988 0 gpio_oeb[5]
rlabel metal3 820 30668 820 30668 0 gpio_oeb[6]
rlabel metal3 820 28628 820 28628 0 gpio_oeb[7]
rlabel metal1 1610 31994 1610 31994 0 gpio_oeb[8]
rlabel metal3 820 32708 820 32708 0 gpio_oeb[9]
rlabel metal1 43056 36890 43056 36890 0 gpio_out[0]
rlabel metal2 61226 38056 61226 38056 0 gpio_out[10]
rlabel metal1 42596 36890 42596 36890 0 gpio_out[11]
rlabel metal1 44850 36890 44850 36890 0 gpio_out[12]
rlabel metal1 52164 36890 52164 36890 0 gpio_out[13]
rlabel metal1 69552 36890 69552 36890 0 gpio_out[14]
rlabel metal1 61778 36890 61778 36890 0 gpio_out[15]
rlabel metal1 62468 36890 62468 36890 0 gpio_out[16]
rlabel metal1 63204 36890 63204 36890 0 gpio_out[17]
rlabel metal1 38778 37434 38778 37434 0 gpio_out[18]
rlabel metal2 42550 1520 42550 1520 0 gpio_out[19]
rlabel metal1 41860 36890 41860 36890 0 gpio_out[1]
rlabel metal2 48346 1520 48346 1520 0 gpio_out[20]
rlabel via2 78246 17051 78246 17051 0 gpio_out[21]
rlabel metal2 39376 2822 39376 2822 0 gpio_out[22]
rlabel metal1 44022 37366 44022 37366 0 gpio_out[23]
rlabel metal2 78246 23341 78246 23341 0 gpio_out[24]
rlabel metal2 43838 1520 43838 1520 0 gpio_out[25]
rlabel metal2 45126 38328 45126 38328 0 gpio_out[26]
rlabel metal1 63756 36890 63756 36890 0 gpio_out[27]
rlabel metal1 46552 37434 46552 37434 0 gpio_out[28]
rlabel metal2 32890 1520 32890 1520 0 gpio_out[29]
rlabel metal1 70840 36890 70840 36890 0 gpio_out[2]
rlabel metal3 751 21828 751 21828 0 gpio_out[30]
rlabel metal3 751 21148 751 21148 0 gpio_out[31]
rlabel metal3 751 19788 751 19788 0 gpio_out[32]
rlabel metal3 1096 20468 1096 20468 0 gpio_out[33]
rlabel metal1 49542 36890 49542 36890 0 gpio_out[34]
rlabel metal1 67620 36890 67620 36890 0 gpio_out[35]
rlabel metal2 53498 38056 53498 38056 0 gpio_out[36]
rlabel metal2 58006 38056 58006 38056 0 gpio_out[37]
rlabel metal1 47012 36890 47012 36890 0 gpio_out[3]
rlabel metal1 66976 36890 66976 36890 0 gpio_out[4]
rlabel metal2 52854 38056 52854 38056 0 gpio_out[5]
rlabel metal1 72128 36890 72128 36890 0 gpio_out[6]
rlabel metal1 64400 36890 64400 36890 0 gpio_out[7]
rlabel metal1 40664 36890 40664 36890 0 gpio_out[8]
rlabel metal1 71484 36890 71484 36890 0 gpio_out[9]
rlabel metal2 47702 38056 47702 38056 0 irq[0]
rlabel metal1 48300 36890 48300 36890 0 irq[1]
rlabel metal1 65044 36890 65044 36890 0 irq[2]
rlabel metal2 8142 15708 8142 15708 0 net1
rlabel metal1 59340 3026 59340 3026 0 net10
rlabel metal1 31142 8908 31142 8908 0 net100
rlabel metal1 35834 15436 35834 15436 0 net101
rlabel metal1 34730 13362 34730 13362 0 net102
rlabel metal1 37628 4998 37628 4998 0 net103
rlabel metal1 38364 15538 38364 15538 0 net104
rlabel metal1 34822 20230 34822 20230 0 net105
rlabel metal1 31004 24718 31004 24718 0 net106
rlabel metal1 39652 16966 39652 16966 0 net107
rlabel metal1 29716 23086 29716 23086 0 net108
rlabel metal1 48944 14790 48944 14790 0 net109
rlabel metal1 59938 2618 59938 2618 0 net11
rlabel metal1 44758 14790 44758 14790 0 net110
rlabel metal1 56166 15572 56166 15572 0 net111
rlabel metal1 52578 9350 52578 9350 0 net112
rlabel metal1 54740 18870 54740 18870 0 net113
rlabel metal2 55246 23936 55246 23936 0 net114
rlabel metal1 53314 23120 53314 23120 0 net115
rlabel metal2 55982 15300 55982 15300 0 net116
rlabel metal1 39238 34170 39238 34170 0 net117
rlabel metal2 44574 19550 44574 19550 0 net118
rlabel metal1 33166 10608 33166 10608 0 net119
rlabel metal1 60214 2550 60214 2550 0 net12
rlabel metal2 34178 14076 34178 14076 0 net120
rlabel metal1 38272 8534 38272 8534 0 net121
rlabel metal2 39790 14722 39790 14722 0 net122
rlabel metal2 31418 25534 31418 25534 0 net123
rlabel metal1 34178 21998 34178 21998 0 net124
rlabel metal1 37950 20502 37950 20502 0 net125
rlabel metal1 36754 18258 36754 18258 0 net126
rlabel metal1 45724 7786 45724 7786 0 net127
rlabel metal2 47978 14620 47978 14620 0 net128
rlabel metal1 54004 6290 54004 6290 0 net129
rlabel metal1 74294 3128 74294 3128 0 net13
rlabel metal1 51336 14314 51336 14314 0 net130
rlabel metal2 53038 17442 53038 17442 0 net131
rlabel metal1 55361 24106 55361 24106 0 net132
rlabel metal2 50370 19414 50370 19414 0 net133
rlabel metal2 52486 8806 52486 8806 0 net134
rlabel metal2 43378 2210 43378 2210 0 net135
rlabel metal1 33879 13906 33879 13906 0 net136
rlabel metal1 37076 12342 37076 12342 0 net137
rlabel metal1 37628 15402 37628 15402 0 net138
rlabel metal2 37306 13804 37306 13804 0 net139
rlabel metal2 71162 2397 71162 2397 0 net14
rlabel metal1 33028 19346 33028 19346 0 net140
rlabel metal2 32614 25619 32614 25619 0 net141
rlabel metal1 35282 20944 35282 20944 0 net142
rlabel metal1 33258 21114 33258 21114 0 net143
rlabel metal1 45402 4556 45402 4556 0 net144
rlabel metal2 42090 8602 42090 8602 0 net145
rlabel metal2 51106 5814 51106 5814 0 net146
rlabel metal2 48530 10880 48530 10880 0 net147
rlabel metal1 55706 24208 55706 24208 0 net148
rlabel metal1 52900 19822 52900 19822 0 net149
rlabel metal1 74152 2618 74152 2618 0 net15
rlabel metal1 51474 17646 51474 17646 0 net150
rlabel metal2 33166 14688 33166 14688 0 net151
rlabel metal2 29762 16932 29762 16932 0 net152
rlabel metal1 44850 2516 44850 2516 0 net153
rlabel metal1 64354 3026 64354 3026 0 net154
rlabel metal1 58558 4114 58558 4114 0 net155
rlabel metal1 10902 17129 10902 17129 0 net156
rlabel metal1 11999 16150 11999 16150 0 net157
rlabel metal2 22034 9962 22034 9962 0 net158
rlabel metal1 32338 13498 32338 13498 0 net159
rlabel metal1 75900 3094 75900 3094 0 net16
rlabel metal1 19511 10642 19511 10642 0 net160
rlabel metal1 10297 21930 10297 21930 0 net161
rlabel metal1 14858 21114 14858 21114 0 net162
rlabel metal1 19596 22678 19596 22678 0 net163
rlabel metal1 23329 25942 23329 25942 0 net164
rlabel metal2 31602 34476 31602 34476 0 net165
rlabel metal1 30314 30226 30314 30226 0 net166
rlabel metal1 34369 8874 34369 8874 0 net167
rlabel metal2 41262 8874 41262 8874 0 net168
rlabel metal1 38962 3400 38962 3400 0 net169
rlabel metal1 61318 2516 61318 2516 0 net17
rlabel metal1 44429 16558 44429 16558 0 net170
rlabel metal1 44620 12818 44620 12818 0 net171
rlabel metal2 46598 9248 46598 9248 0 net172
rlabel metal2 52946 4590 52946 4590 0 net173
rlabel metal1 53169 12138 53169 12138 0 net174
rlabel metal1 46690 18217 46690 18217 0 net175
rlabel metal1 55805 18326 55805 18326 0 net176
rlabel metal2 33442 21216 33442 21216 0 net177
rlabel metal2 41170 20706 41170 20706 0 net178
rlabel metal2 37490 36414 37490 36414 0 net179
rlabel metal1 73094 2856 73094 2856 0 net18
rlabel metal1 43049 34646 43049 34646 0 net180
rlabel metal1 45041 36822 45041 36822 0 net181
rlabel metal1 56396 22610 56396 22610 0 net182
rlabel metal1 51375 24106 51375 24106 0 net183
rlabel metal1 49358 32946 49358 32946 0 net184
rlabel metal1 37720 21930 37720 21930 0 net185
rlabel metal1 19596 12206 19596 12206 0 net186
rlabel metal1 24731 16082 24731 16082 0 net187
rlabel metal2 27554 14093 27554 14093 0 net188
rlabel metal2 40526 36992 40526 36992 0 net189
rlabel metal2 65366 2176 65366 2176 0 net19
rlabel metal1 73370 36754 73370 36754 0 net190
rlabel metal1 55476 36754 55476 36754 0 net191
rlabel metal1 51704 36754 51704 36754 0 net192
rlabel metal1 41400 36754 41400 36754 0 net193
rlabel metal2 68310 36550 68310 36550 0 net194
rlabel metal1 58788 36754 58788 36754 0 net195
rlabel metal2 48806 36550 48806 36550 0 net196
rlabel metal1 59432 36754 59432 36754 0 net197
rlabel metal1 60444 36686 60444 36686 0 net198
rlabel metal1 46046 36686 46046 36686 0 net199
rlabel metal2 7682 14212 7682 14212 0 net2
rlabel metal1 66056 2278 66056 2278 0 net20
rlabel metal1 56120 36754 56120 36754 0 net200
rlabel metal1 54188 36754 54188 36754 0 net201
rlabel metal1 56856 36754 56856 36754 0 net202
rlabel metal2 60674 36550 60674 36550 0 net203
rlabel metal1 51060 36754 51060 36754 0 net204
rlabel metal2 43102 36550 43102 36550 0 net205
rlabel metal1 42044 36754 42044 36754 0 net206
rlabel metal1 71024 36754 71024 36754 0 net207
rlabel metal1 47196 36754 47196 36754 0 net208
rlabel metal1 67160 36754 67160 36754 0 net209
rlabel metal1 74888 2618 74888 2618 0 net21
rlabel metal2 52946 36550 52946 36550 0 net210
rlabel metal2 72266 36550 72266 36550 0 net211
rlabel metal1 64584 36754 64584 36754 0 net212
rlabel metal2 40894 36992 40894 36992 0 net213
rlabel metal1 71668 36754 71668 36754 0 net214
rlabel metal2 61042 36550 61042 36550 0 net215
rlabel metal2 42550 36550 42550 36550 0 net216
rlabel metal1 44850 36346 44850 36346 0 net217
rlabel metal1 52348 36754 52348 36754 0 net218
rlabel metal1 69736 36754 69736 36754 0 net219
rlabel metal1 67298 2516 67298 2516 0 net22
rlabel metal1 61916 36754 61916 36754 0 net220
rlabel metal1 62652 36754 62652 36754 0 net221
rlabel metal2 63158 36550 63158 36550 0 net222
rlabel metal1 63940 36754 63940 36754 0 net223
rlabel metal1 49680 36754 49680 36754 0 net224
rlabel metal1 67804 36754 67804 36754 0 net225
rlabel metal2 53314 36550 53314 36550 0 net226
rlabel metal2 58098 36550 58098 36550 0 net227
rlabel metal2 47794 36550 47794 36550 0 net228
rlabel metal1 48484 36754 48484 36754 0 net229
rlabel metal1 72312 2414 72312 2414 0 net23
rlabel metal1 65228 36754 65228 36754 0 net230
rlabel metal1 66516 36754 66516 36754 0 net231
rlabel metal1 73048 36686 73048 36686 0 net232
rlabel metal1 70380 36754 70380 36754 0 net233
rlabel metal1 54832 36754 54832 36754 0 net234
rlabel metal1 50416 36754 50416 36754 0 net235
rlabel metal1 57500 36754 57500 36754 0 net236
rlabel metal1 69092 36754 69092 36754 0 net237
rlabel metal1 65872 36754 65872 36754 0 net238
rlabel metal1 2070 23120 2070 23120 0 net239
rlabel metal1 72726 2482 72726 2482 0 net24
rlabel metal2 2070 31484 2070 31484 0 net240
rlabel metal2 2162 23358 2162 23358 0 net241
rlabel metal1 2116 25874 2116 25874 0 net242
rlabel metal1 2116 27438 2116 27438 0 net243
rlabel metal1 2116 30226 2116 30226 0 net244
rlabel metal1 2116 30702 2116 30702 0 net245
rlabel metal1 2116 28526 2116 28526 0 net246
rlabel metal2 2070 32062 2070 32062 0 net247
rlabel metal1 2116 32878 2116 32878 0 net248
rlabel metal1 2116 33966 2116 33966 0 net249
rlabel metal1 72634 2550 72634 2550 0 net25
rlabel metal2 2070 26622 2070 26622 0 net250
rlabel metal1 2116 25262 2116 25262 0 net251
rlabel metal2 2070 23868 2070 23868 0 net252
rlabel metal2 2070 29308 2070 29308 0 net253
rlabel metal1 2116 33490 2116 33490 0 net254
rlabel metal2 2070 34748 2070 34748 0 net255
rlabel metal1 2116 35666 2116 35666 0 net256
rlabel metal1 2070 36176 2070 36176 0 net257
rlabel metal1 2116 24786 2116 24786 0 net258
rlabel metal1 2116 28050 2116 28050 0 net259
rlabel metal1 71392 2618 71392 2618 0 net26
rlabel metal2 2162 36414 2162 36414 0 net260
rlabel metal2 14582 20060 14582 20060 0 net261
rlabel metal1 18768 18734 18768 18734 0 net262
rlabel metal1 17935 19414 17935 19414 0 net263
rlabel metal1 31602 30260 31602 30260 0 net264
rlabel metal2 21298 18428 21298 18428 0 net265
rlabel metal1 41032 2414 41032 2414 0 net266
rlabel metal1 38686 2414 38686 2414 0 net267
rlabel metal1 43654 2414 43654 2414 0 net268
rlabel metal1 9476 24174 9476 24174 0 net269
rlabel metal1 68494 2550 68494 2550 0 net27
rlabel metal1 56534 3468 56534 3468 0 net270
rlabel metal2 31602 29308 31602 29308 0 net271
rlabel metal2 42826 30668 42826 30668 0 net272
rlabel metal1 13110 19856 13110 19856 0 net273
rlabel metal1 36800 34034 36800 34034 0 net274
rlabel metal1 28198 31314 28198 31314 0 net275
rlabel metal1 28980 33626 28980 33626 0 net276
rlabel metal1 30820 31450 30820 31450 0 net277
rlabel metal1 31096 32402 31096 32402 0 net278
rlabel metal2 10258 18938 10258 18938 0 net279
rlabel metal1 58604 2618 58604 2618 0 net28
rlabel metal1 21298 25908 21298 25908 0 net280
rlabel metal1 28980 35054 28980 35054 0 net281
rlabel metal2 13662 24378 13662 24378 0 net282
rlabel metal1 12696 14246 12696 14246 0 net283
rlabel metal2 9890 18428 9890 18428 0 net284
rlabel metal1 29394 30260 29394 30260 0 net285
rlabel metal1 18262 16490 18262 16490 0 net286
rlabel metal1 17434 16218 17434 16218 0 net287
rlabel metal1 13662 30294 13662 30294 0 net288
rlabel metal1 28566 32878 28566 32878 0 net289
rlabel metal1 72680 2822 72680 2822 0 net29
rlabel metal1 33028 36754 33028 36754 0 net290
rlabel metal1 19964 27438 19964 27438 0 net291
rlabel metal1 16514 14042 16514 14042 0 net292
rlabel metal1 14122 12818 14122 12818 0 net293
rlabel metal1 35696 31858 35696 31858 0 net294
rlabel metal1 32154 12886 32154 12886 0 net295
rlabel metal1 19458 23698 19458 23698 0 net296
rlabel metal1 17342 31790 17342 31790 0 net297
rlabel metal1 13340 27438 13340 27438 0 net298
rlabel metal1 17802 30702 17802 30702 0 net299
rlabel metal1 8418 14994 8418 14994 0 net3
rlabel metal1 70242 2550 70242 2550 0 net30
rlabel metal1 18308 30702 18308 30702 0 net300
rlabel metal2 12834 30906 12834 30906 0 net301
rlabel metal1 38502 28526 38502 28526 0 net302
rlabel metal2 15594 17408 15594 17408 0 net303
rlabel metal2 13294 17884 13294 17884 0 net304
rlabel metal1 51520 11730 51520 11730 0 net305
rlabel metal1 12558 15334 12558 15334 0 net306
rlabel metal1 14766 15572 14766 15572 0 net307
rlabel metal1 10764 29138 10764 29138 0 net308
rlabel metal1 17066 21998 17066 21998 0 net309
rlabel metal2 52486 2074 52486 2074 0 net31
rlabel metal1 20148 25874 20148 25874 0 net310
rlabel metal1 47518 16218 47518 16218 0 net311
rlabel metal1 20976 29274 20976 29274 0 net312
rlabel metal1 46736 7854 46736 7854 0 net313
rlabel metal1 14536 24786 14536 24786 0 net314
rlabel metal2 13110 22780 13110 22780 0 net315
rlabel metal1 15042 22202 15042 22202 0 net316
rlabel metal1 48760 23698 48760 23698 0 net317
rlabel metal1 18722 30226 18722 30226 0 net318
rlabel metal1 38364 7854 38364 7854 0 net319
rlabel metal1 67160 2822 67160 2822 0 net32
rlabel metal1 35604 36754 35604 36754 0 net320
rlabel metal2 10626 20060 10626 20060 0 net321
rlabel metal2 32154 18938 32154 18938 0 net322
rlabel metal2 10718 22916 10718 22916 0 net323
rlabel metal2 11454 30906 11454 30906 0 net324
rlabel metal1 38778 33490 38778 33490 0 net325
rlabel metal1 45724 16762 45724 16762 0 net326
rlabel metal1 37536 35734 37536 35734 0 net327
rlabel metal1 48990 24208 48990 24208 0 net328
rlabel metal1 20608 28186 20608 28186 0 net329
rlabel metal1 70058 2618 70058 2618 0 net33
rlabel metal1 16008 28050 16008 28050 0 net330
rlabel metal1 48530 10064 48530 10064 0 net331
rlabel metal2 17710 12172 17710 12172 0 net332
rlabel metal1 34086 32912 34086 32912 0 net333
rlabel metal1 16100 30702 16100 30702 0 net334
rlabel metal1 52394 7310 52394 7310 0 net335
rlabel metal1 39146 8942 39146 8942 0 net336
rlabel metal2 10534 28220 10534 28220 0 net337
rlabel metal1 36386 34544 36386 34544 0 net338
rlabel metal1 57592 3502 57592 3502 0 net339
rlabel metal2 46414 2142 46414 2142 0 net34
rlabel metal1 38042 17204 38042 17204 0 net340
rlabel metal1 44850 14926 44850 14926 0 net341
rlabel metal1 33580 5134 33580 5134 0 net342
rlabel metal1 27140 9690 27140 9690 0 net343
rlabel metal1 49128 14382 49128 14382 0 net344
rlabel metal1 53774 9554 53774 9554 0 net345
rlabel metal1 54096 8398 54096 8398 0 net346
rlabel metal1 35834 6766 35834 6766 0 net347
rlabel metal1 30728 7854 30728 7854 0 net348
rlabel metal1 39100 20910 39100 20910 0 net349
rlabel metal1 66608 2618 66608 2618 0 net35
rlabel metal1 37168 20434 37168 20434 0 net350
rlabel metal1 43332 14926 43332 14926 0 net351
rlabel metal2 52026 25092 52026 25092 0 net352
rlabel metal1 42688 11118 42688 11118 0 net353
rlabel metal1 51474 20910 51474 20910 0 net354
rlabel metal1 46690 9554 46690 9554 0 net355
rlabel metal1 32338 9554 32338 9554 0 net356
rlabel metal1 49956 26350 49956 26350 0 net357
rlabel metal1 41860 6766 41860 6766 0 net358
rlabel metal1 34684 18734 34684 18734 0 net359
rlabel metal1 54372 2618 54372 2618 0 net36
rlabel metal1 33580 7310 33580 7310 0 net360
rlabel metal1 31740 7378 31740 7378 0 net361
rlabel metal1 43608 13294 43608 13294 0 net362
rlabel metal2 40894 8602 40894 8602 0 net363
rlabel metal1 38870 11662 38870 11662 0 net364
rlabel metal1 53452 26350 53452 26350 0 net365
rlabel metal1 50048 5134 50048 5134 0 net366
rlabel metal1 46598 17646 46598 17646 0 net367
rlabel metal1 40480 20434 40480 20434 0 net368
rlabel metal1 49404 8466 49404 8466 0 net369
rlabel metal2 54878 2244 54878 2244 0 net37
rlabel metal1 55200 9520 55200 9520 0 net370
rlabel metal1 42320 17646 42320 17646 0 net371
rlabel metal1 53544 16082 53544 16082 0 net372
rlabel metal1 40986 14926 40986 14926 0 net373
rlabel metal1 52992 13906 52992 13906 0 net374
rlabel metal1 36248 15470 36248 15470 0 net375
rlabel metal1 41446 9554 41446 9554 0 net376
rlabel metal1 46092 12206 46092 12206 0 net377
rlabel metal1 34040 8466 34040 8466 0 net378
rlabel metal1 40986 3978 40986 3978 0 net379
rlabel metal1 58650 3366 58650 3366 0 net38
rlabel metal1 34454 15470 34454 15470 0 net380
rlabel metal1 38548 15470 38548 15470 0 net381
rlabel metal1 57270 22610 57270 22610 0 net382
rlabel metal1 38042 5134 38042 5134 0 net383
rlabel metal1 53728 18190 53728 18190 0 net384
rlabel metal1 37030 10642 37030 10642 0 net385
rlabel metal1 53498 20910 53498 20910 0 net386
rlabel metal1 53452 11118 53452 11118 0 net387
rlabel metal1 43838 35054 43838 35054 0 net388
rlabel metal1 41124 12750 41124 12750 0 net389
rlabel metal1 58558 2278 58558 2278 0 net39
rlabel metal1 35604 13294 35604 13294 0 net390
rlabel metal1 49036 18734 49036 18734 0 net391
rlabel metal1 52578 5202 52578 5202 0 net392
rlabel metal2 43746 17340 43746 17340 0 net393
rlabel metal2 56166 16388 56166 16388 0 net394
rlabel metal1 35328 20434 35328 20434 0 net395
rlabel metal1 43976 4046 43976 4046 0 net396
rlabel metal1 33948 19822 33948 19822 0 net397
rlabel metal1 41722 4114 41722 4114 0 net398
rlabel metal1 37030 4114 37030 4114 0 net399
rlabel metal1 1610 15368 1610 15368 0 net4
rlabel metal2 59386 3876 59386 3876 0 net40
rlabel metal1 39008 6222 39008 6222 0 net400
rlabel metal1 56028 20910 56028 20910 0 net401
rlabel metal1 51658 18190 51658 18190 0 net402
rlabel metal2 32982 10438 32982 10438 0 net403
rlabel metal1 34086 9588 34086 9588 0 net404
rlabel metal2 33902 10404 33902 10404 0 net405
rlabel metal1 53774 23086 53774 23086 0 net406
rlabel metal1 29348 33966 29348 33966 0 net407
rlabel metal1 13340 30362 13340 30362 0 net408
rlabel metal1 14214 23834 14214 23834 0 net409
rlabel metal1 58742 3434 58742 3434 0 net41
rlabel metal1 39284 37162 39284 37162 0 net42
rlabel metal1 43976 2482 43976 2482 0 net43
rlabel metal1 49220 2550 49220 2550 0 net44
rlabel metal1 77970 17170 77970 17170 0 net45
rlabel metal1 39422 2890 39422 2890 0 net46
rlabel metal1 43976 37162 43976 37162 0 net47
rlabel metal2 58558 23494 58558 23494 0 net48
rlabel metal1 41354 2924 41354 2924 0 net49
rlabel metal1 55269 2414 55269 2414 0 net5
rlabel metal2 44390 36754 44390 36754 0 net50
rlabel metal2 46138 37026 46138 37026 0 net51
rlabel metal1 32752 2822 32752 2822 0 net52
rlabel metal2 7038 21488 7038 21488 0 net53
rlabel metal1 7498 20434 7498 20434 0 net54
rlabel metal1 1702 19788 1702 19788 0 net55
rlabel metal1 4301 20910 4301 20910 0 net56
rlabel metal1 57914 2448 57914 2448 0 net57
rlabel metal1 53544 2822 53544 2822 0 net58
rlabel metal1 47104 2822 47104 2822 0 net59
rlabel metal1 53728 2550 53728 2550 0 net6
rlabel metal2 72910 2890 72910 2890 0 net60
rlabel metal1 51244 2822 51244 2822 0 net61
rlabel metal1 61870 2414 61870 2414 0 net62
rlabel metal2 51658 2618 51658 2618 0 net63
rlabel metal2 68678 2618 68678 2618 0 net64
rlabel metal1 63802 2414 63802 2414 0 net65
rlabel metal1 45816 2822 45816 2822 0 net66
rlabel metal1 49036 2822 49036 2822 0 net67
rlabel metal1 49772 2414 49772 2414 0 net68
rlabel metal2 63250 2618 63250 2618 0 net69
rlabel metal2 59386 2108 59386 2108 0 net7
rlabel metal1 64446 2414 64446 2414 0 net70
rlabel metal1 76682 2822 76682 2822 0 net71
rlabel metal2 78062 2618 78062 2618 0 net72
rlabel metal1 62514 2414 62514 2414 0 net73
rlabel metal1 46460 2822 46460 2822 0 net74
rlabel metal2 47794 2618 47794 2618 0 net75
rlabel metal1 72818 3094 72818 3094 0 net76
rlabel metal1 78016 7378 78016 7378 0 net77
rlabel metal2 78062 8262 78062 8262 0 net78
rlabel metal1 78154 5678 78154 5678 0 net79
rlabel metal1 54694 2516 54694 2516 0 net8
rlabel metal1 78246 7888 78246 7888 0 net80
rlabel metal2 78062 6460 78062 6460 0 net81
rlabel metal1 36386 4080 36386 4080 0 net82
rlabel metal2 36662 20604 36662 20604 0 net83
rlabel metal2 39514 18649 39514 18649 0 net84
rlabel metal1 49082 13294 49082 13294 0 net85
rlabel metal2 52854 11458 52854 11458 0 net86
rlabel metal1 51244 25874 51244 25874 0 net87
rlabel metal1 46046 17680 46046 17680 0 net88
rlabel metal1 55246 22576 55246 22576 0 net89
rlabel metal1 59248 2822 59248 2822 0 net9
rlabel metal1 29946 14382 29946 14382 0 net90
rlabel metal1 30544 24786 30544 24786 0 net91
rlabel metal1 34316 25874 34316 25874 0 net92
rlabel metal1 47380 19754 47380 19754 0 net93
rlabel metal1 45126 20910 45126 20910 0 net94
rlabel metal1 41630 8500 41630 8500 0 net95
rlabel metal2 36202 14212 36202 14212 0 net96
rlabel metal1 38732 14382 38732 14382 0 net97
rlabel metal2 47794 17578 47794 17578 0 net98
rlabel metal2 54234 14416 54234 14416 0 net99
rlabel metal2 54326 3332 54326 3332 0 team_11_WB.EN_VAL_REG
rlabel metal2 18078 17578 18078 17578 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[0\]
rlabel metal1 12190 17544 12190 17544 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[1\]
rlabel metal2 20654 16864 20654 16864 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[2\]
rlabel metal2 15502 18394 15502 18394 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[3\]
rlabel metal2 14674 15674 14674 15674 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[4\]
rlabel metal1 16146 13872 16146 13872 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[5\]
rlabel metal2 13846 13056 13846 13056 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[6\]
rlabel metal2 12374 14688 12374 14688 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[7\]
rlabel metal1 19136 17102 19136 17102 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[0\]
rlabel metal2 14306 17646 14306 17646 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[1\]
rlabel metal1 12972 16218 12972 16218 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[2\]
rlabel metal1 16330 17782 16330 17782 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[3\]
rlabel metal1 15732 16014 15732 16014 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[4\]
rlabel metal1 17020 14450 17020 14450 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[5\]
rlabel metal1 14674 11866 14674 11866 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[6\]
rlabel metal2 13478 14688 13478 14688 0 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[7\]
rlabel metal2 31970 3808 31970 3808 0 team_11_WB.instance_to_wrap.kp.buffertop.nrst
rlabel metal1 12604 22066 12604 22066 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[0\]
rlabel metal2 9522 28356 9522 28356 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[10\]
rlabel metal1 11040 29682 11040 29682 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[11\]
rlabel metal1 12466 30260 12466 30260 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[12\]
rlabel metal1 13754 31246 13754 31246 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[13\]
rlabel via2 14582 30141 14582 30141 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[14\]
rlabel metal2 17986 28866 17986 28866 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[15\]
rlabel metal1 17526 28526 17526 28526 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[16\]
rlabel metal1 15640 30294 15640 30294 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[17\]
rlabel metal2 18538 31994 18538 31994 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[18\]
rlabel metal1 19780 31246 19780 31246 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[19\]
rlabel metal1 14582 23086 14582 23086 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[1\]
rlabel metal2 19090 29886 19090 29886 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[20\]
rlabel metal2 22402 29478 22402 29478 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[21\]
rlabel metal1 20562 27302 20562 27302 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[22\]
rlabel metal1 20378 27506 20378 27506 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[23\]
rlabel metal1 20562 26282 20562 26282 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[24\]
rlabel metal1 20792 25874 20792 25874 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[25\]
rlabel metal2 21114 24004 21114 24004 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[26\]
rlabel metal2 17710 25313 17710 25313 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[27\]
rlabel metal2 17986 25568 17986 25568 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[28\]
rlabel metal2 17342 24956 17342 24956 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[29\]
rlabel metal1 15180 24786 15180 24786 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[2\]
rlabel metal2 13478 24548 13478 24548 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[3\]
rlabel metal1 10672 21862 10672 21862 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[4\]
rlabel metal2 10902 24480 10902 24480 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[5\]
rlabel metal1 9844 24718 9844 24718 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[6\]
rlabel metal2 12466 25840 12466 25840 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[7\]
rlabel metal2 14674 27098 14674 27098 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[8\]
rlabel metal2 12926 25840 12926 25840 0 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[9\]
rlabel metal2 13938 21726 13938 21726 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[0\]
rlabel metal1 10074 28118 10074 28118 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[10\]
rlabel metal1 10166 29070 10166 29070 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[11\]
rlabel metal1 10442 30906 10442 30906 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[12\]
rlabel metal1 12282 30906 12282 30906 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[13\]
rlabel metal1 13248 29206 13248 29206 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[14\]
rlabel metal1 16514 28118 16514 28118 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[15\]
rlabel via1 16139 27642 16139 27642 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[16\]
rlabel metal1 15410 31654 15410 31654 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[17\]
rlabel metal1 17296 31994 17296 31994 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[18\]
rlabel metal2 18538 31076 18538 31076 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[19\]
rlabel metal1 14214 22066 14214 22066 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[1\]
rlabel metal2 20470 29342 20470 29342 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[20\]
rlabel metal1 20654 29546 20654 29546 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[21\]
rlabel metal1 21252 27098 21252 27098 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[22\]
rlabel metal2 18538 27166 18538 27166 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[23\]
rlabel metal1 22494 25806 22494 25806 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[24\]
rlabel metal1 19274 25194 19274 25194 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[25\]
rlabel metal1 19734 23698 19734 23698 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[26\]
rlabel metal2 17618 23902 17618 23902 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[27\]
rlabel metal1 16790 22202 16790 22202 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[28\]
rlabel metal1 16928 24786 16928 24786 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[29\]
rlabel metal2 14766 24684 14766 24684 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[2\]
rlabel metal2 11914 24412 11914 24412 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[3\]
rlabel metal1 11460 22202 11460 22202 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[4\]
rlabel metal2 9062 23902 9062 23902 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[5\]
rlabel metal2 9062 24548 9062 24548 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[6\]
rlabel metal1 13708 26894 13708 26894 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[7\]
rlabel metal1 13156 27574 13156 27574 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[8\]
rlabel metal1 10212 26282 10212 26282 0 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[9\]
rlabel metal2 24150 12036 24150 12036 0 team_11_WB.instance_to_wrap.kp.controlstop.mode
rlabel metal1 32154 3026 32154 3026 0 team_11_WB.instance_to_wrap.kp.controlstop.msg_tx_ctrl
rlabel metal1 28658 14926 28658 14926 0 team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl
rlabel metal1 17181 12410 17181 12410 0 team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[0\]
rlabel metal1 18768 12206 18768 12206 0 team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[1\]
rlabel metal2 19228 11220 19228 11220 0 team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[2\]
rlabel metal1 19826 10778 19826 10778 0 team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[3\]
rlabel metal2 23874 18564 23874 18564 0 team_11_WB.instance_to_wrap.kp.controlstop.upper
rlabel metal1 14168 20366 14168 20366 0 team_11_WB.instance_to_wrap.kp.debouncertop.keyvalid
rlabel metal1 18998 19244 18998 19244 0 team_11_WB.instance_to_wrap.kp.debouncertop.next_receive_ready
rlabel metal1 18216 18802 18216 18802 0 team_11_WB.instance_to_wrap.kp.debouncertop.receive_ready
rlabel metal2 36570 18972 36570 18972 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[0\]
rlabel metal1 36662 5236 36662 5236 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[100\]
rlabel metal1 38226 25874 38226 25874 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[101\]
rlabel metal1 51658 25806 51658 25806 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[102\]
rlabel metal1 36064 13906 36064 13906 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[103\]
rlabel metal1 35374 17646 35374 17646 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[104\]
rlabel metal2 45678 8126 45678 8126 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[105\]
rlabel metal2 55062 11322 55062 11322 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[106\]
rlabel via1 47886 17646 47886 17646 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[107\]
rlabel metal1 38502 8432 38502 8432 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[108\]
rlabel metal1 37858 24718 37858 24718 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[109\]
rlabel metal1 24196 13158 24196 13158 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[10\]
rlabel metal1 49634 24106 49634 24106 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[110\]
rlabel metal1 34822 12614 34822 12614 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[111\]
rlabel metal1 34960 19278 34960 19278 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[112\]
rlabel metal1 47058 10064 47058 10064 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[113\]
rlabel metal1 50876 9554 50876 9554 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[114\]
rlabel metal1 45540 16626 45540 16626 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[115\]
rlabel metal2 39330 7344 39330 7344 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[116\]
rlabel metal1 39721 25126 39721 25126 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[117\]
rlabel metal1 49082 23154 49082 23154 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[118\]
rlabel metal2 39882 13022 39882 13022 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[119\]
rlabel metal2 45494 15487 45494 15487 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[11\]
rlabel metal1 32798 19380 32798 19380 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[120\]
rlabel metal1 45678 8568 45678 8568 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[121\]
rlabel metal2 52302 11900 52302 11900 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[122\]
rlabel metal1 48622 16456 48622 16456 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[123\]
rlabel metal2 37674 8398 37674 8398 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[124\]
rlabel metal2 37582 24276 37582 24276 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[125\]
rlabel metal1 49174 22950 49174 22950 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[126\]
rlabel metal1 33074 12716 33074 12716 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[127\]
rlabel via2 34362 9571 34362 9571 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[12\]
rlabel metal2 30222 22508 30222 22508 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[13\]
rlabel via2 29486 18173 29486 18173 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[14\]
rlabel via2 34086 13923 34086 13923 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[15\]
rlabel metal1 37030 17680 37030 17680 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[16\]
rlabel metal2 43378 10880 43378 10880 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[17\]
rlabel metal1 49128 10778 49128 10778 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[18\]
rlabel metal2 50416 14382 50416 14382 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[19\]
rlabel metal2 29854 9129 29854 9129 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[1\]
rlabel metal1 33304 10030 33304 10030 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[20\]
rlabel metal1 33166 22610 33166 22610 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[21\]
rlabel metal2 50002 21216 50002 21216 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[22\]
rlabel metal1 34914 14790 34914 14790 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[23\]
rlabel via1 38961 16558 38961 16558 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[24\]
rlabel metal1 41262 8500 41262 8500 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[25\]
rlabel metal1 50094 9622 50094 9622 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[26\]
rlabel metal1 48070 14484 48070 14484 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[27\]
rlabel metal1 33718 9146 33718 9146 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[28\]
rlabel metal1 30452 22610 30452 22610 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[29\]
rlabel metal2 31234 11305 31234 11305 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[2\]
rlabel viali 50738 21522 50738 21522 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[30\]
rlabel metal2 36570 14076 36570 14076 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[31\]
rlabel metal1 44666 17714 44666 17714 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[32\]
rlabel metal1 43010 9520 43010 9520 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[33\]
rlabel via1 50462 10030 50462 10030 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[34\]
rlabel metal1 50830 14382 50830 14382 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[35\]
rlabel via1 32228 8942 32228 8942 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[36\]
rlabel metal1 33386 22610 33386 22610 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[37\]
rlabel metal1 52256 19822 52256 19822 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[38\]
rlabel viali 36109 14382 36109 14382 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[39\]
rlabel metal1 33442 15538 33442 15538 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[3\]
rlabel metal1 39790 19312 39790 19312 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[40\]
rlabel via1 41537 8466 41537 8466 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[41\]
rlabel metal1 50324 7378 50324 7378 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[42\]
rlabel viali 51198 14382 51198 14382 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[43\]
rlabel metal2 32798 7956 32798 7956 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[44\]
rlabel metal2 30958 24310 30958 24310 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[45\]
rlabel metal1 52026 23018 52026 23018 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[46\]
rlabel viali 37858 14382 37858 14382 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[47\]
rlabel metal1 38318 20400 38318 20400 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[48\]
rlabel metal1 41124 6766 41124 6766 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[49\]
rlabel metal2 33258 10047 33258 10047 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[4\]
rlabel via1 50737 5678 50737 5678 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[50\]
rlabel metal2 52302 15810 52302 15810 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[51\]
rlabel metal1 35282 5610 35282 5610 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[52\]
rlabel metal1 31648 24174 31648 24174 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[53\]
rlabel metal2 54602 22797 54602 22797 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[54\]
rlabel metal1 42550 14450 42550 14450 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[55\]
rlabel metal1 37950 21590 37950 21590 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[56\]
rlabel metal2 40526 6885 40526 6885 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[57\]
rlabel via1 51584 10030 51584 10030 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[58\]
rlabel metal2 53774 16337 53774 16337 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[59\]
rlabel metal1 39054 22610 39054 22610 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[5\]
rlabel metal1 32660 6358 32660 6358 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[60\]
rlabel metal1 35006 23630 35006 23630 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[61\]
rlabel metal1 55476 23290 55476 23290 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[62\]
rlabel via1 41538 14382 41538 14382 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[63\]
rlabel metal1 36018 20808 36018 20808 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[64\]
rlabel via1 41924 5678 41924 5678 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[65\]
rlabel metal1 53774 7344 53774 7344 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[66\]
rlabel metal2 55062 16286 55062 16286 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[67\]
rlabel via1 34822 5678 34822 5678 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[68\]
rlabel metal1 34914 25194 34914 25194 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[69\]
rlabel metal2 29854 19873 29854 19873 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[6\]
rlabel metal1 55338 24820 55338 24820 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[70\]
rlabel metal2 46874 12444 46874 12444 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[71\]
rlabel metal1 37122 21454 37122 21454 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[72\]
rlabel metal1 44666 4794 44666 4794 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[73\]
rlabel metal2 51658 8670 51658 8670 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[74\]
rlabel metal1 53038 17646 53038 17646 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[75\]
rlabel metal1 34730 5270 34730 5270 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[76\]
rlabel metal2 34546 25772 34546 25772 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[77\]
rlabel metal1 51014 24854 51014 24854 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[78\]
rlabel metal1 40158 11662 40158 11662 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[79\]
rlabel metal1 32568 13974 32568 13974 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[7\]
rlabel metal1 34592 20366 34592 20366 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[80\]
rlabel via1 43120 5202 43120 5202 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[81\]
rlabel metal1 52302 9928 52302 9928 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[82\]
rlabel metal1 51060 18326 51060 18326 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[83\]
rlabel metal2 36432 5202 36432 5202 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[84\]
rlabel metal1 35374 25262 35374 25262 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[85\]
rlabel metal2 52578 23902 52578 23902 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[86\]
rlabel via1 38226 13294 38226 13294 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[87\]
rlabel metal2 35374 17884 35374 17884 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[88\]
rlabel metal2 44850 6766 44850 6766 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[89\]
rlabel metal2 37030 16592 37030 16592 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[8\]
rlabel metal1 55016 10030 55016 10030 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[90\]
rlabel metal2 52486 18598 52486 18598 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[91\]
rlabel metal1 37122 5610 37122 5610 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[92\]
rlabel metal1 36662 26928 36662 26928 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[93\]
rlabel metal1 52164 26350 52164 26350 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[94\]
rlabel metal1 36708 13158 36708 13158 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[95\]
rlabel metal2 34822 16694 34822 16694 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[96\]
rlabel metal1 44712 5882 44712 5882 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[97\]
rlabel viali 52026 10030 52026 10030 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[98\]
rlabel metal1 50371 18224 50371 18224 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[99\]
rlabel metal1 29532 12070 29532 12070 0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[9\]
rlabel metal2 10810 19040 10810 19040 0 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[0\]
rlabel metal2 10718 18156 10718 18156 0 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[1\]
rlabel metal1 9752 17238 9752 17238 0 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[2\]
rlabel metal2 13018 19550 13018 19550 0 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[3\]
rlabel metal2 8326 15844 8326 15844 0 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[4\]
rlabel metal1 8050 13974 8050 13974 0 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[5\]
rlabel metal1 9338 13192 9338 13192 0 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[6\]
rlabel metal1 9384 14926 9384 14926 0 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[7\]
rlabel metal2 11546 20706 11546 20706 0 team_11_WB.instance_to_wrap.kp.keypadtop.next_keyvalid
rlabel metal2 38226 35938 38226 35938 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[0\]
rlabel metal2 29946 32946 29946 32946 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[10\]
rlabel metal2 29486 33626 29486 33626 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[11\]
rlabel metal1 29210 32300 29210 32300 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[12\]
rlabel metal1 29854 31722 29854 31722 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[13\]
rlabel metal1 29900 31110 29900 31110 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[14\]
rlabel metal1 30452 30158 30452 30158 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[15\]
rlabel metal2 32154 30464 32154 30464 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[16\]
rlabel metal1 32844 30566 32844 30566 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[17\]
rlabel metal2 39514 36312 39514 36312 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[1\]
rlabel metal1 36554 36822 36554 36822 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[2\]
rlabel metal1 35972 36890 35972 36890 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[3\]
rlabel via1 35374 34510 35374 34510 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[4\]
rlabel metal1 35650 33524 35650 33524 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[5\]
rlabel metal2 33074 33422 33074 33422 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[6\]
rlabel metal1 32614 33864 32614 33864 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[7\]
rlabel metal1 32154 36346 32154 36346 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[8\]
rlabel metal1 32430 34000 32430 34000 0 team_11_WB.instance_to_wrap.sending.cnt_20ms\[9\]
rlabel metal1 35972 30022 35972 30022 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[0\]
rlabel metal1 45494 32436 45494 32436 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[10\]
rlabel metal1 45402 32232 45402 32232 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[11\]
rlabel metal1 44988 35258 44988 35258 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[12\]
rlabel metal1 44758 36550 44758 36550 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[13\]
rlabel metal2 44298 33286 44298 33286 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[14\]
rlabel metal2 37674 30192 37674 30192 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[1\]
rlabel metal2 37490 30906 37490 30906 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[2\]
rlabel metal1 39928 30158 39928 30158 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[3\]
rlabel metal2 42182 33388 42182 33388 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[4\]
rlabel viali 41814 33493 41814 33493 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[5\]
rlabel metal2 42458 33728 42458 33728 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[6\]
rlabel metal1 41860 33286 41860 33286 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[7\]
rlabel metal1 44666 33558 44666 33558 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[8\]
rlabel metal1 46368 31994 46368 31994 0 team_11_WB.instance_to_wrap.sending.cnt_500hz\[9\]
rlabel metal2 47518 28866 47518 28866 0 team_11_WB.instance_to_wrap.sending.currentState\[0\]
rlabel metal1 45402 29138 45402 29138 0 team_11_WB.instance_to_wrap.sending.currentState\[1\]
rlabel metal1 45770 26384 45770 26384 0 team_11_WB.instance_to_wrap.sending.currentState\[2\]
rlabel metal2 40894 28866 40894 28866 0 team_11_WB.instance_to_wrap.sending.currentState\[3\]
rlabel metal2 41262 26622 41262 26622 0 team_11_WB.instance_to_wrap.sending.currentState\[4\]
rlabel metal1 46322 28424 46322 28424 0 team_11_WB.instance_to_wrap.sending.currentState\[5\]
rlabel metal2 45908 36380 45908 36380 0 team_11_WB.instance_to_wrap.sending.lcd_en
rlabel metal1 44298 36142 44298 36142 0 team_11_WB.instance_to_wrap.sending.lcd_rs
rlabel metal2 34086 20179 34086 20179 0 wb_clk_i
rlabel metal1 50646 2380 50646 2380 0 wb_rst_i
rlabel metal2 57362 1656 57362 1656 0 wbs_ack_o
rlabel metal2 52854 1520 52854 1520 0 wbs_adr_i[0]
rlabel metal2 59294 1520 59294 1520 0 wbs_adr_i[10]
rlabel metal1 54188 2414 54188 2414 0 wbs_adr_i[11]
rlabel metal2 56258 748 56258 748 0 wbs_adr_i[12]
rlabel metal1 56626 3536 56626 3536 0 wbs_adr_i[13]
rlabel metal2 59938 1520 59938 1520 0 wbs_adr_i[14]
rlabel metal2 60582 1520 60582 1520 0 wbs_adr_i[15]
rlabel metal1 78798 3026 78798 3026 0 wbs_adr_i[16]
rlabel metal2 70886 1520 70886 1520 0 wbs_adr_i[17]
rlabel metal2 74106 1520 74106 1520 0 wbs_adr_i[18]
rlabel metal2 77326 1520 77326 1520 0 wbs_adr_i[19]
rlabel metal2 61226 1520 61226 1520 0 wbs_adr_i[1]
rlabel metal2 76038 1520 76038 1520 0 wbs_adr_i[20]
rlabel metal2 65090 1520 65090 1520 0 wbs_adr_i[21]
rlabel metal2 65734 1520 65734 1520 0 wbs_adr_i[22]
rlabel metal2 75394 1520 75394 1520 0 wbs_adr_i[23]
rlabel metal2 67022 1520 67022 1520 0 wbs_adr_i[24]
rlabel metal1 72036 2414 72036 2414 0 wbs_adr_i[25]
rlabel metal2 74750 1520 74750 1520 0 wbs_adr_i[26]
rlabel metal1 73646 2346 73646 2346 0 wbs_adr_i[27]
rlabel metal2 71530 1520 71530 1520 0 wbs_adr_i[28]
rlabel metal2 67666 1520 67666 1520 0 wbs_adr_i[29]
rlabel metal1 58144 2414 58144 2414 0 wbs_adr_i[2]
rlabel metal2 77970 1588 77970 1588 0 wbs_adr_i[30]
rlabel metal2 68954 1520 68954 1520 0 wbs_adr_i[31]
rlabel metal2 52210 1520 52210 1520 0 wbs_adr_i[3]
rlabel metal2 69598 1520 69598 1520 0 wbs_adr_i[4]
rlabel metal2 70242 1520 70242 1520 0 wbs_adr_i[5]
rlabel metal2 45126 1622 45126 1622 0 wbs_adr_i[6]
rlabel metal2 66240 2278 66240 2278 0 wbs_adr_i[7]
rlabel metal1 53958 2346 53958 2346 0 wbs_adr_i[8]
rlabel metal2 45218 2244 45218 2244 0 wbs_adr_i[9]
rlabel metal1 57546 2448 57546 2448 0 wbs_cyc_i
rlabel metal1 58834 2346 58834 2346 0 wbs_dat_i[0]
rlabel metal2 53498 1520 53498 1520 0 wbs_dat_o[0]
rlabel metal2 47058 1520 47058 1520 0 wbs_dat_o[10]
rlabel metal2 72818 1520 72818 1520 0 wbs_dat_o[11]
rlabel metal2 50922 1520 50922 1520 0 wbs_dat_o[12]
rlabel metal2 61870 1520 61870 1520 0 wbs_dat_o[13]
rlabel metal1 70196 36890 70196 36890 0 wbs_dat_o[14]
rlabel metal2 51566 1520 51566 1520 0 wbs_dat_o[15]
rlabel metal2 68310 1520 68310 1520 0 wbs_dat_o[16]
rlabel metal1 54694 36890 54694 36890 0 wbs_dat_o[17]
rlabel metal2 63802 1520 63802 1520 0 wbs_dat_o[18]
rlabel metal2 45770 1520 45770 1520 0 wbs_dat_o[19]
rlabel metal2 48990 1520 48990 1520 0 wbs_dat_o[1]
rlabel metal1 50232 36890 50232 36890 0 wbs_dat_o[20]
rlabel metal2 49634 1520 49634 1520 0 wbs_dat_o[21]
rlabel metal1 57316 36890 57316 36890 0 wbs_dat_o[22]
rlabel metal2 63158 1520 63158 1520 0 wbs_dat_o[23]
rlabel metal1 68908 36890 68908 36890 0 wbs_dat_o[24]
rlabel metal2 64446 1520 64446 1520 0 wbs_dat_o[25]
rlabel metal2 76682 1520 76682 1520 0 wbs_dat_o[26]
rlabel metal2 78614 1520 78614 1520 0 wbs_dat_o[27]
rlabel metal2 62514 1520 62514 1520 0 wbs_dat_o[28]
rlabel metal1 65596 36890 65596 36890 0 wbs_dat_o[29]
rlabel metal2 46414 959 46414 959 0 wbs_dat_o[2]
rlabel metal2 47702 1520 47702 1520 0 wbs_dat_o[30]
rlabel metal2 43194 1656 43194 1656 0 wbs_dat_o[31]
rlabel metal2 78246 7021 78246 7021 0 wbs_dat_o[3]
rlabel metal2 66240 36890 66240 36890 0 wbs_dat_o[4]
rlabel metal2 78246 8279 78246 8279 0 wbs_dat_o[5]
rlabel via2 78430 5525 78430 5525 0 wbs_dat_o[6]
rlabel metal2 78430 7633 78430 7633 0 wbs_dat_o[7]
rlabel metal1 72680 36890 72680 36890 0 wbs_dat_o[8]
rlabel via2 78246 6171 78246 6171 0 wbs_dat_o[9]
rlabel metal2 78522 4369 78522 4369 0 wbs_stb_i
rlabel metal2 78338 5015 78338 5015 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 80000 40000
<< end >>
