* NGSPICE file created from team_08_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

.subckt team_08_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4]
+ la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_0_94_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7963_ _0487_ _0493_ vssd1 vssd1 vccd1 vccd1 _3502_ sky130_fd_sc_hd__or2_1
X_6914_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[9\]
+ _2708_ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__and2_1
X_7894_ net160 _3443_ _3445_ net166 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9242__SET_B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout162_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8906__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9633_ net484 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_76_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6845_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[9\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__or4_1
XFILLER_0_64_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6917__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9564_ net432 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_92_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6776_ net684 _2615_ _2617_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5727_ _1620_ _1622_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__or2_1
X_9495_ net370 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
X_8515_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ _3333_ _3352_ vssd1 vssd1 vccd1 vccd1 _3995_ sky130_fd_sc_hd__nor3_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7981__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8446_ _3925_ _3926_ vssd1 vssd1 vccd1 vccd1 _3927_ sky130_fd_sc_hd__or2_1
X_5658_ _0798_ _1602_ _1610_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5589_ _1485_ _1541_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_96_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8377_ _3858_ _3843_ _2875_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__a2bb2o_1
X_4609_ net261 _0566_ _0568_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[4\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7328_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[18\]
+ _2995_ vssd1 vssd1 vccd1 vccd1 _2996_ sky130_fd_sc_hd__or2_1
XANTENNA__4829__B _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8842__B1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7259_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[10\]
+ _2942_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9529__404 vssd1 vssd1 vccd1 vccd1 _9529__404/HI net404 sky130_fd_sc_hd__conb_1
XANTENNA__9432__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7221__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8373__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4580__A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7581__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8987__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7884__A1 _3403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4755__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8061__A1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4960_ _0737_ net145 vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__nand2_4
X_4891_ _0806_ _0843_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6630_ _2519_ _2520_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[24\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6561_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[12\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[14\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[15\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2476_ sky130_fd_sc_hd__and4bb_1
X_5512_ _0907_ _1464_ _1462_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8300_ _0500_ _3501_ _3508_ _3515_ vssd1 vssd1 vccd1 vccd1 _3793_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9280_ clknet_leaf_13_wb_clk_i _0123_ net213 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6492_ _0516_ _0535_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__and2_1
X_5443_ _0883_ _1395_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__nand2_1
XANTENNA__7875__B2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8231_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[15\]
+ _2992_ vssd1 vssd1 vccd1 vccd1 _3734_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6210__A _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5374_ _1309_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__nor2_1
X_8162_ _0654_ _3678_ _3681_ net161 net237 vssd1 vssd1 vccd1 vccd1 _3682_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7088__C1 _2828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7113_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[8\] _2844_
+ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout138 _0817_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_4
X_8093_ _0644_ _3621_ vssd1 vssd1 vccd1 vccd1 _3622_ sky130_fd_sc_hd__or2_2
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout127 _3214_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_4
Xfanout105 _3271_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_4
Xfanout116 _3225_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_4
X_7044_ _2790_ _2791_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout149 net151 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6063__B1 _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4576__A1_N net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8995_ clknet_leaf_3_wb_clk_i _0159_ net202 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7946_ net332 net329 vssd1 vssd1 vccd1 vccd1 _3486_ sky130_fd_sc_hd__nand2_1
X_7877_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[13\]
+ _3431_ _3403_ vssd1 vssd1 vccd1 vccd1 _3434_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9616_ net480 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
X_6828_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[7\]
+ net562 _2648_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6366__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6759_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__or4b_1
X_9547_ net415 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6118__B2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9478_ net353 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XANTENNA__8600__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5943__B _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8429_ _3319_ net94 _3322_ vssd1 vssd1 vccd1 vccd1 _3910_ sky130_fd_sc_hd__a21o_1
XANTENNA__6120__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold170 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[4\]
+ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8043__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6357__A1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6357__B2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5090_ _1038_ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4916__C _0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5992_ _1907_ _1941_ _1940_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_8780_ net174 _3335_ _3886_ _4257_ vssd1 vssd1 vccd1 vccd1 _4258_ sky130_fd_sc_hd__a31o_1
X_7800_ net290 _3377_ _3385_ net292 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__a22o_1
X_4943_ _0894_ _0895_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7731_ net124 net117 _3307_ vssd1 vssd1 vccd1 vccd1 _3321_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7662_ _3246_ _3248_ _3251_ vssd1 vssd1 vccd1 vccd1 _3252_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4874_ _0824_ _0825_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7545__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9401_ clknet_leaf_32_wb_clk_i _0348_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_6613_ net618 _2507_ net262 vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7593_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\]
+ net184 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\]
+ net176 vssd1 vssd1 vccd1 vccd1 _3183_ sky130_fd_sc_hd__nand4_1
XFILLER_0_28_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9332_ clknet_leaf_53_wb_clk_i _0015_ net201 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_6544_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[18\] _2461_
+ vssd1 vssd1 vccd1 vccd1 _2462_ sky130_fd_sc_hd__and2_1
XANTENNA__8420__A _3329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9263_ clknet_leaf_10_wb_clk_i _0085_ net226 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6475_ net158 vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5426_ _1372_ _1375_ _1377_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8214_ _2989_ _3722_ vssd1 vssd1 vccd1 vccd1 _3723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9194_ clknet_leaf_11_wb_clk_i _0028_ net226 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5357_ _1303_ _1307_ _1308_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__or3_1
X_8145_ _0657_ _3480_ _3667_ net278 vssd1 vssd1 vccd1 vccd1 _3668_ sky130_fd_sc_hd__a211o_1
X_5288_ _1236_ _1240_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__nand2_1
X_8076_ _0706_ _3605_ vssd1 vssd1 vccd1 vccd1 _3606_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7027_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[5\] team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8978_ net311 vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__inv_2
X_7929_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[2\] _3469_ vssd1
+ vssd1 vccd1 vccd1 _3470_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8500__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4857__X _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7067__A2 _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6009__B _0926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5848__B _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4752__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4590_ net191 _0405_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__nand2_2
XFILLER_0_49_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6260_ _2059_ _2118_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4646__A_N _0573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8894__B net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6191_ _1394_ _2143_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__nor2_1
X_5211_ _1147_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5142_ _1093_ _1094_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5073_ _1023_ _1025_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__xor2_1
X_8901_ _3271_ _4376_ _4377_ vssd1 vssd1 vccd1 vccd1 _4378_ sky130_fd_sc_hd__a21oi_1
X_8832_ _3933_ _4308_ _4309_ _3286_ vssd1 vssd1 vccd1 vccd1 _4310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5975_ _1924_ _1927_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__nand2_1
X_8763_ net95 _4239_ vssd1 vssd1 vccd1 vccd1 _4241_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4926_ _0818_ _0878_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout242_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8694_ _3305_ _4113_ _4165_ _4166_ _4172_ vssd1 vssd1 vccd1 vccd1 _4173_ sky130_fd_sc_hd__a41o_1
X_7714_ _3301_ _3303_ _3295_ vssd1 vssd1 vccd1 vccd1 _3304_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4857_ _0781_ _0790_ _0605_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__a21o_4
XFILLER_0_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7645_ _3231_ _3233_ vssd1 vssd1 vccd1 vccd1 _3235_ sky130_fd_sc_hd__nand2_2
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9210__RESET_B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7576_ net257 _3174_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_60_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8730__A2 _3789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4788_ _0718_ _0740_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__nand2_1
X_6527_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[11\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[12\]
+ _2447_ vssd1 vssd1 vccd1 vccd1 _2451_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9315_ clknet_leaf_3_wb_clk_i _0286_ net202 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9246_ clknet_leaf_11_wb_clk_i _0097_ net217 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6458_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[3\]
+ _2400_ vssd1 vssd1 vccd1 vccd1 _2401_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5409_ _1358_ _1360_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__and2_1
X_9177_ clknet_leaf_10_wb_clk_i _0040_ net227 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6389_ team_08_WB.instance_to_wrap.allocation.game.game.score\[5\] _2339_ vssd1 vssd1
+ vccd1 vccd1 _2340_ sky130_fd_sc_hd__or2_2
XFILLER_0_101_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8128_ _0698_ _3643_ vssd1 vssd1 vccd1 vccd1 _3654_ sky130_fd_sc_hd__or2_1
XANTENNA__8246__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8309__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5014__A _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8059_ net603 net242 _3020_ _3456_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_67_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8325__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8549__A2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9369__RESET_B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7509__B1 _3022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8182__B1 _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5760_ _1661_ _1709_ _1710_ _1712_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8522__X _4001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8960__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5691_ _1610_ _1643_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4711_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[2\] _0647_
+ _0664_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4642_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[7\] vssd1
+ vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7430_ _0441_ net308 vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7361_ _0637_ net275 vssd1 vssd1 vccd1 vccd1 _3015_ sky130_fd_sc_hd__nor2_2
X_4573_ net316 _0535_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6312_ _0450_ _0451_ vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__nor2_1
X_7292_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[22\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[21\]
+ _2964_ vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__and3_1
X_9100_ clknet_leaf_53_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[30\]
+ net200 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6243_ _1693_ _2130_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9031_ clknet_leaf_52_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[13\]
+ net207 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_6174_ _2125_ _2126_ _1834_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5125_ _1033_ _1035_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5056_ _0824_ _0835_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5769__A _0919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5121__X _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8815_ net329 net189 vssd1 vssd1 vccd1 vccd1 _4293_ sky130_fd_sc_hd__and2b_1
X_5958_ _0724_ _0860_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_62_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8746_ _4203_ _4204_ _4207_ _4209_ _4223_ vssd1 vssd1 vccd1 vccd1 _4224_ sky130_fd_sc_hd__o221a_1
X_9603__467 vssd1 vssd1 vccd1 vccd1 _9603__467/HI net467 sky130_fd_sc_hd__conb_1
X_4909_ _0810_ _0860_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5889_ _1839_ _1840_ _1838_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__a21bo_1
X_8677_ net283 _3621_ vssd1 vssd1 vccd1 vccd1 _4156_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8703__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7628_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[8\]
+ _3204_ _3217_ vssd1 vssd1 vccd1 vccd1 _3218_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7559_ net258 _3165_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8467__A1 _3279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9229_ clknet_leaf_21_wb_clk_i _0057_ net240 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4567__B _0505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[1\]
+ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.clk1
+ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[3\]
+ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[16\] vssd1
+ vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold96 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[15\] vssd1 vssd1
+ vccd1 vccd1 net594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[6\] vssd1 vssd1
+ vccd1 vccd1 net583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8458__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9122__Q team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6930_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6861_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[4\]
+ _2670_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8394__B1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9580_ net444 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5812_ _1763_ _1764_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__nand2b_1
X_6792_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[10\]
+ _2625_ _2627_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8600_ net109 _3596_ vssd1 vssd1 vccd1 vccd1 _4079_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5743_ _0754_ _0910_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__nor2_1
XANTENNA__5747__A2 _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8531_ _0663_ net113 vssd1 vssd1 vccd1 vccd1 _4010_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5674_ _1618_ _1625_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8462_ net154 _3904_ _3909_ _3312_ net174 vssd1 vssd1 vccd1 vccd1 _3943_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4625_ _0581_ _0582_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7413_ _0440_ _3055_ _3056_ _0438_ net302 vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__o2111ai_1
X_8393_ _3867_ _3872_ vssd1 vssd1 vccd1 vccd1 _3874_ sky130_fd_sc_hd__nand2_1
X_4556_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[3\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[5\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7344_ net536 _2998_ vssd1 vssd1 vccd1 vccd1 _3007_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout205_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7275_ net577 _2954_ _2956_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__a21oi_1
X_4487_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[1\] vssd1
+ vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6226_ _1248_ _2148_ _1191_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_55_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9014_ clknet_leaf_6_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[4\]
+ net212 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__6880__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6157_ _2108_ _2109_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5108_ _1037_ _1060_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_51_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout195_X net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7698__B _3241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6088_ _2039_ _2040_ _2038_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_51_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5039_ net123 _0946_ _0948_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7420__B1_N team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_cactus
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8924__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4850__B _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7219__A _0423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8137__B1 _3662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8729_ _4204_ _4206_ _4203_ vssd1 vssd1 vccd1 vccd1 _4207_ sky130_fd_sc_hd__or3b_1
XANTENNA__6123__A _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9538__494 vssd1 vssd1 vccd1 vccd1 net494 _9538__494/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_75_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6623__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5390_ _1342_ _1340_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_22_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4488__A team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7060_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[1\]
+ _2789_ _2792_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__a22o_1
Xfanout309 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_2
XANTENNA__5665__A1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6011_ _1961_ _1962_ _1963_ vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8603__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7962_ _0487_ _0493_ vssd1 vssd1 vccd1 vccd1 _3501_ sky130_fd_sc_hd__nor2_1
X_6913_ net272 _2707_ _2708_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__nor3_1
X_9632_ net264 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
X_7893_ _3444_ vssd1 vssd1 vccd1 vccd1 _3445_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6844_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__or4b_1
XFILLER_0_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8423__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9563_ net431 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6775_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[4\]
+ _2615_ net274 vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8142__B net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9494_ net369 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
XFILLER_0_91_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5726_ _1676_ _1677_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout322_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8514_ _3332_ _3954_ _3963_ vssd1 vssd1 vccd1 vccd1 _3994_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8445_ net154 net94 _3885_ _3321_ _3324_ vssd1 vssd1 vccd1 vccd1 _3926_ sky130_fd_sc_hd__o221a_1
X_5657_ _1608_ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__nand2_1
XANTENNA__6878__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout110_X net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5588_ _1483_ _1484_ _1476_ _1479_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_96_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8376_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[7\] _3855_ vssd1
+ vssd1 vccd1 vccd1 _3858_ sky130_fd_sc_hd__xor2_1
X_4608_ _0501_ _0567_ _0540_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7327_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[17\]
+ _2994_ vssd1 vssd1 vccd1 vccd1 _2995_ sky130_fd_sc_hd__or2_1
X_4539_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[11\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[13\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_53_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8842__A1 _0423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7258_ _2944_ _2945_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6209_ _2160_ _2161_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7189_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[12\] _2894_ vssd1
+ vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9609__473 vssd1 vssd1 vccd1 vccd1 _9609__473/HI net473 sky130_fd_sc_hd__conb_1
XFILLER_0_67_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4861__A _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7581__B2 _2368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5692__A _0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5895__A1 _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input40_X net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4755__B _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8061__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4890_ _0841_ _0842_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6560_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[9\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[11\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__and4bb_1
X_5511_ _1462_ _1463_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6491_ _0638_ _0639_ _2427_ net294 vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
X_5442_ _0849_ _0862_ _0848_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8230_ _3732_ _3733_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__nand2_1
XANTENNA__6210__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5373_ _1277_ _1325_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8161_ _3679_ _3680_ vssd1 vssd1 vccd1 vccd1 _3681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8092_ net288 _0643_ vssd1 vssd1 vccd1 vccd1 _3621_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7112_ _0454_ _2844_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_91_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout128 _0939_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_4
XANTENNA__9235__RESET_B net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7043_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[0\]
+ _0458_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__or3_1
Xfanout106 _3252_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__buf_4
Xfanout117 net120 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_4
Xfanout139 _0701_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_4
XANTENNA_fanout272_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8994_ clknet_leaf_4_wb_clk_i _0158_ net204 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4952__Y _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7945_ _0494_ _3483_ vssd1 vssd1 vccd1 vccd1 _3485_ sky130_fd_sc_hd__xor2_1
XANTENNA__4681__A _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7876_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[12\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[13\] _3428_
+ vssd1 vssd1 vccd1 vccd1 _3433_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout158_X net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9615_ net479 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
X_6827_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[7\]
+ _2648_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9546_ net414 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_98_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6758_ net524 _2602_ _2604_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5709_ _1660_ _1661_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__and2_1
X_6689_ _0464_ _2556_ _2559_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6118__A2 _0926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9477_ net352 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_6_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8428_ _3315_ _3879_ vssd1 vssd1 vccd1 vccd1 _3909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6120__B _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8359_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[1\] _2874_ _3846_
+ _0561_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold171 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[3\]
+ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7079__B1 _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[10\] vssd1
+ vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold182 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__9321__SET_B net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8047__B net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8043__A2 _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8063__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7306__A1 _0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5868__Y _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5991_ net143 _1943_ _0744_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__o21a_1
X_4942_ _0889_ _0893_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7730_ _3318_ _3319_ vssd1 vssd1 vccd1 vccd1 _3320_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7661_ _3245_ _3250_ vssd1 vssd1 vccd1 vccd1 _3251_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4873_ _0825_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__inv_2
X_9400_ clknet_leaf_31_wb_clk_i _0347_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_6612_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[17\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[18\]
+ _2505_ vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7592_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[11\]
+ _3180_ _3181_ vssd1 vssd1 vccd1 vccd1 _3182_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9331_ clknet_leaf_53_wb_clk_i _0014_ net201 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6543_ _2461_ _2428_ _2460_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[17\]
+ sky130_fd_sc_hd__and3b_1
X_9262_ clknet_leaf_10_wb_clk_i _0084_ net227 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_6474_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[24\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[23\]
+ _2416_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[25\]
+ vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_93_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5425_ _1372_ _1375_ _1377_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8213_ net661 _2988_ vssd1 vssd1 vccd1 vccd1 _3722_ sky130_fd_sc_hd__nand2_1
X_9193_ clknet_leaf_16_wb_clk_i _0027_ net228 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5356_ _1303_ _1307_ _1308_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__o21ai_1
XANTENNA__8258__C1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8144_ _0654_ net161 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _3667_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5287_ _1239_ _1237_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_11_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8075_ net183 _0704_ vssd1 vssd1 vccd1 vccd1 _3605_ sky130_fd_sc_hd__and2b_1
XANTENNA__5350__A_N _0999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7026_ _0429_ net3 vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7987__A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8977_ net311 vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__inv_2
XANTENNA__7784__A1 _2368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7928_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[1\] team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3469_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7859_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[8\] _3416_
+ vssd1 vssd1 vccd1 vccd1 _3421_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9529_ net404 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_80_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5970__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4586__A _0551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5210_ _1148_ _1162_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__nand2_1
X_9473__348 vssd1 vssd1 vccd1 vccd1 _9473__348/HI net348 sky130_fd_sc_hd__conb_1
X_6190_ _2140_ _2142_ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__and2_1
XANTENNA__4496__A team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5141_ _0746_ _1091_ _1092_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8255__A2 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5072_ _0959_ _0966_ _0964_ _0861_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__a211o_1
X_9514__389 vssd1 vssd1 vccd1 vccd1 _9514__389/HI net389 sky130_fd_sc_hd__conb_1
X_8900_ _3271_ _4376_ _2275_ vssd1 vssd1 vccd1 vccd1 _4377_ sky130_fd_sc_hd__o21a_1
XANTENNA__7215__B1 _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7766__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8831_ _3300_ _3860_ _3869_ vssd1 vssd1 vccd1 vccd1 _4309_ sky130_fd_sc_hd__nor3_1
XFILLER_0_94_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8762_ _4239_ net95 net100 _4238_ vssd1 vssd1 vccd1 vccd1 _4240_ sky130_fd_sc_hd__a2bb2o_1
X_5974_ _1924_ _1925_ _1926_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7713_ net153 _3302_ vssd1 vssd1 vccd1 vccd1 _3303_ sky130_fd_sc_hd__nor2_1
X_4925_ _0876_ _0877_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8693_ _4161_ _4162_ _4170_ _4171_ vssd1 vssd1 vccd1 vccd1 _4172_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_23_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4856_ _0781_ _0790_ _0605_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout235_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7644_ _3231_ _3233_ vssd1 vssd1 vccd1 vccd1 _3234_ sky130_fd_sc_hd__and2_2
X_7575_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr2\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr2\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.clk1 vssd1
+ vssd1 vccd1 vccd1 _3174_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4787_ _0724_ net144 vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9314_ clknet_leaf_3_wb_clk_i _0285_ net202 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_6526_ _2449_ _2450_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[11\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9250__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9245_ clknet_leaf_15_wb_clk_i _0096_ net215 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6457_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2400_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8494__A2 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5408_ _1358_ _1360_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__nor2_1
X_9176_ clknet_leaf_19_wb_clk_i _0035_ net229 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6388_ team_08_WB.instance_to_wrap.allocation.game.game.score\[3\] team_08_WB.instance_to_wrap.allocation.game.game.score\[4\]
+ _2338_ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__or3_1
X_5339_ _1281_ _1284_ _1291_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__a21o_1
X_8127_ _0698_ _3643_ vssd1 vssd1 vccd1 vccd1 _3653_ sky130_fd_sc_hd__nand2_1
XANTENNA__8246__A2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8309__C _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8058_ _3586_ _3591_ _3592_ net239 net589 vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__o32a_1
X_7009_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[5\] team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_67_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5301__Y _1254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8325__B net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7509__A1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8341__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8060__B net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6385__C_N _2324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7693__B1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7404__B net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _1608_ _1609_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4710_ _0664_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7419__X _3064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4641_ _0576_ _0598_ _0575_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__a21o_1
XANTENNA__9079__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4572_ _0540_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__inv_2
X_7360_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[7\] _2975_
+ _3013_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__a21bo_1
X_9555__423 vssd1 vssd1 vccd1 vccd1 _9555__423/HI net423 sky130_fd_sc_hd__conb_1
XFILLER_0_80_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6311_ _2261_ _2262_ _2263_ _0635_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__o22ai_1
X_7291_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[21\]
+ _2964_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[22\]
+ vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6242_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[19\]
+ _2193_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__and2_1
X_9030_ clknet_leaf_52_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[12\]
+ net207 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4497__Y _0134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7684__B1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6993__X net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6173_ _1832_ _1833_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5124_ net130 _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4954__A _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5055_ _1006_ _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout185_A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8814_ _4290_ _4291_ vssd1 vssd1 vccd1 vccd1 _4292_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_9_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5488__C _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5957_ _1908_ _1909_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4960__Y _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8745_ _4211_ _4221_ _4222_ vssd1 vssd1 vccd1 vccd1 _4223_ sky130_fd_sc_hd__or3_1
XANTENNA__5785__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4908_ _0809_ _0859_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout140_X net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8676_ _3864_ _4112_ _4113_ _4154_ _4152_ vssd1 vssd1 vccd1 vccd1 _4155_ sky130_fd_sc_hd__a41o_1
X_5888_ _1838_ _1839_ _1840_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout238_X net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7627_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[9\]
+ net126 vssd1 vssd1 vccd1 vccd1 _3217_ sky130_fd_sc_hd__xnor2_2
X_4839_ net140 vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7558_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr1\[1\] team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr1\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.clk1 vssd1
+ vssd1 vccd1 vccd1 _3165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9495__370 vssd1 vssd1 vccd1 vccd1 _9495__370/HI net370 sky130_fd_sc_hd__conb_1
XFILLER_0_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7489_ _0439_ net309 _0442_ net306 vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__a22o_1
X_6509_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[6\] _2437_
+ vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__and2_1
XANTENNA__8467__A2 _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9228_ clknet_leaf_18_wb_clk_i _0056_ net230 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9159_ _0134_ _0405_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ sky130_fd_sc_hd__dfxtp_4
Xhold20 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[8\] vssd1
+ vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[20\] vssd1
+ vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4864__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold64 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 _3157_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.clk1
+ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[8\]
+ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[19\]
+ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4583__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5695__A _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8155__B2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5141__A1 _0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7418__B1 _3022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8091__B1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9585__449 vssd1 vssd1 vccd1 vccd1 _9585__449/HI net449 sky130_fd_sc_hd__conb_1
XFILLER_0_89_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6860_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[4\]
+ _2670_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8394__A1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5811_ _0924_ _1716_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__xnor2_1
X_6791_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[10\]
+ _2625_ net274 vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5742_ _1649_ _1650_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8530_ net118 _3674_ vssd1 vssd1 vccd1 vccd1 _4009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5673_ _1625_ _1618_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8461_ _3876_ _3903_ _3934_ _3941_ _3929_ vssd1 vssd1 vccd1 vccd1 _3942_ sky130_fd_sc_hd__a311o_1
XFILLER_0_53_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4624_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[4\] vssd1
+ vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8392_ _3872_ vssd1 vssd1 vccd1 vccd1 _3873_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9479__354 vssd1 vssd1 vccd1 vccd1 _9479__354/HI net354 sky130_fd_sc_hd__conb_1
X_7412_ net302 _0438_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__nand2_1
X_4555_ _0523_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__inv_2
X_7343_ _2997_ _3006_ _3002_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_38_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout100_A _3265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4486_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__inv_2
X_7274_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[16\]
+ _2954_ net180 vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__o21ai_1
X_9013_ clknet_leaf_8_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[3\]
+ net223 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6225_ _1138_ _2150_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_55_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _2100_ _2101_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5107_ _1058_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__nor2_1
XANTENNA__8082__B1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6087_ _2035_ _2037_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4659__A_N team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5038_ _0901_ _0951_ _0990_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6989_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2754_ sky130_fd_sc_hd__xnor2_1
X_8728_ net97 _4202_ _4205_ net103 vssd1 vssd1 vccd1 vccd1 _4206_ sky130_fd_sc_hd__o22ai_1
XANTENNA__8137__A1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6123__B _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8659_ _4120_ _4133_ _4135_ net150 _4124_ vssd1 vssd1 vccd1 vccd1 _4138_ sky130_fd_sc_hd__o221a_1
XANTENNA__7896__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4859__A _0573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7360__A2 _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XANTENNA__4865__Y _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input30_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4882__B1 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4594__A _0425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4769__A _0719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8851__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6010_ _0718_ _0928_ _0930_ net168 vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7961_ _0487_ _0493_ vssd1 vssd1 vccd1 vccd1 _3500_ sky130_fd_sc_hd__nand2_1
X_7892_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[17\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[18\] _3439_
+ vssd1 vssd1 vccd1 vccd1 _3444_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6912_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[8\]
+ _2704_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__and3_1
X_9631_ net266 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
X_6843_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__or2_1
XANTENNA__9094__RESET_B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8423__B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9562_ net430 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_99_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6774_ _0465_ _2613_ _2616_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5725_ _1677_ _1676_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__and2b_1
X_9493_ net368 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_72_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8513_ _3958_ _3973_ _3992_ _3341_ vssd1 vssd1 vccd1 vccd1 _3993_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5656_ _0798_ _1601_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout315_A team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8444_ _3319_ net94 _3324_ vssd1 vssd1 vccd1 vccd1 _3925_ sky130_fd_sc_hd__a21oi_1
X_4607_ _0484_ _0497_ _0500_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__and3_1
X_5587_ _1537_ _1539_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_96_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8375_ _3857_ _3843_ _2875_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_5_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7326_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[16\]
+ _2993_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__or2_1
X_4538_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[3\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[4\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout103_X net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8842__A2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7257_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[10\]
+ _2942_ net179 vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4469_ net310 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6208_ _1196_ _1251_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_70_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7188_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[12\] _2894_ vssd1
+ vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_5_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _2090_ _2091_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__or2_1
XANTENNA__7802__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8614__A _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4861__B _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6134__A _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5344__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5895__A2 _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8599__A1_N net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8524__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5867__B _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8349__B2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8349__A1 _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5510_ _0814_ net145 _1461_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6490_ _0463_ _2425_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__nand2_1
X_5441_ _1345_ _1391_ _1392_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5372_ net128 _1276_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__or2_1
X_8160_ net286 _2388_ vssd1 vssd1 vccd1 vccd1 _3680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8285__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8091_ _3617_ _3618_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 _3620_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7111_ _2844_ _2845_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__nor2_1
Xfanout129 net132 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_91_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7042_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[3\] vssd1
+ vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__nand2b_1
Xfanout107 _3252_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_2
Xfanout118 net119 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_2
XFILLER_0_38_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8993_ clknet_leaf_2_wb_clk_i _0157_ net204 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4962__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7944_ _0494_ _3483_ vssd1 vssd1 vccd1 vccd1 _3484_ sky130_fd_sc_hd__and2_1
XANTENNA__6653__S _2532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7875_ _3431_ _3432_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[12\]
+ net166 vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__a2bb2o_1
X_9614_ net478 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_65_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6826_ net673 _2648_ _2650_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6757_ net524 _2602_ net268 vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9545_ net413 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_18_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5708_ _0791_ _0929_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__nor2_1
XANTENNA__5793__A _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6688_ net274 _2558_ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9476_ net351 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_21_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5639_ _1588_ _1590_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8427_ _3278_ _3355_ _3907_ vssd1 vssd1 vccd1 vccd1 _3908_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8358_ _3469_ _3845_ _3842_ vssd1 vssd1 vccd1 vccd1 _3846_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5017__B _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7309_ _2977_ _2980_ vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__nand2_1
Xhold150 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[4\] vssd1 vssd1
+ vccd1 vccd1 net659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold172 net69 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__dlygate4sd3_1
X_8289_ _3779_ _3781_ _3782_ vssd1 vssd1 vccd1 vccd1 _3783_ sky130_fd_sc_hd__or3b_1
Xhold194 team_08_WB.instance_to_wrap.allocation.game.game.score\[0\] vssd1 vssd1 vccd1
+ vccd1 net692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7003__A1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7306__A2 _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8078__X _3608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5990_ _0717_ _0860_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4941_ _0889_ _0893_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4872_ net167 _0762_ _0774_ _0796_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__o22a_4
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7660_ _3217_ _3249_ vssd1 vssd1 vccd1 vccd1 _3250_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6611_ _2507_ _2508_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[17\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9330_ clknet_leaf_53_wb_clk_i _0013_ net201 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_7591_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[16\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[15\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\]
+ _0455_ vssd1 vssd1 vccd1 vccd1 _3181_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6542_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[17\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[16\]
+ _2457_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9261_ clknet_leaf_10_wb_clk_i _0083_ net227 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6473_ _2403_ _2414_ _2415_ _2412_ vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5424_ _1355_ _1376_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__xnor2_1
X_9192_ clknet_leaf_17_wb_clk_i _0026_ net228 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8212_ _3034_ _3721_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__nand2_1
X_8143_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\] net243
+ _3480_ _3666_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5355_ _1252_ _1254_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5286_ _1236_ _1238_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__nand2_1
X_8074_ _3597_ _3601_ _3604_ net243 net605 vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__o32a_1
X_7025_ _2774_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.tft_dc
+ net3 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__mux2_1
XANTENNA__7987__B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8435__Y _3916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout268_X net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout170_X net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8164__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8976_ net311 vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__inv_2
X_7927_ _3464_ _3465_ _3467_ _2268_ vssd1 vssd1 vccd1 vccd1 _3468_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7858_ net159 _3419_ _3420_ net165 net680 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_26_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6809_ net270 _2633_ _2639_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8733__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7789_ _3373_ _3375_ _2380_ vssd1 vssd1 vccd1 vccd1 _3376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9528_ net403 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_36_Left_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9459_ clknet_leaf_44_wb_clk_i _0397_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_cactus
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8500__A4 _3895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5970__B _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_45_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4873__Y _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5698__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8724__A1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5140_ _0746_ _1091_ _1092_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__and3_1
X_5071_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_63_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8830_ net108 net106 _3930_ _3932_ vssd1 vssd1 vccd1 vccd1 _4308_ sky130_fd_sc_hd__a31o_1
X_5973_ _0723_ _0928_ _1889_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__a21o_1
X_8761_ net316 _4233_ _4235_ vssd1 vssd1 vccd1 vccd1 _4239_ sky130_fd_sc_hd__o21a_1
X_4924_ _0745_ _0830_ _0832_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_35_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7712_ net124 net120 vssd1 vssd1 vccd1 vccd1 _3302_ sky130_fd_sc_hd__nand2_2
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8692_ _4157_ _4164_ vssd1 vssd1 vccd1 vccd1 _4171_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_23_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4855_ _0784_ net140 vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_72_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7643_ _3221_ _3232_ vssd1 vssd1 vccd1 vccd1 _3233_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout130_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4786_ _0736_ _0737_ _0634_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__a21o_1
X_7574_ _3172_ _3173_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6525_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[11\] _2447_
+ net156 vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9313_ clknet_leaf_1_wb_clk_i _0284_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_win
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__9316__Q team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9244_ clknet_leaf_12_wb_clk_i _0091_ net218 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6456_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[3\] _2325_
+ _2381_ _2399_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a22o_1
XANTENNA__5135__X _1088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5407_ _1312_ _1359_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4687__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9175_ _0150_ _0412_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_6387_ team_08_WB.instance_to_wrap.allocation.game.game.score\[2\] _2326_ _2336_
+ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5338_ _1288_ _1289_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_81_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9290__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8126_ net608 net243 _3644_ _3652_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__o22a_1
X_8057_ net314 _2426_ net277 vssd1 vssd1 vccd1 vccd1 _3592_ sky130_fd_sc_hd__a21o_1
X_7008_ _0467_ _0468_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] _2764_
+ _2766_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__a311o_1
X_5269_ _1219_ _1221_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__nor2_4
XFILLER_0_98_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8954__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8959_ net281 net154 net127 net286 _4117_ vssd1 vssd1 vccd1 vccd1 _4436_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_90_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7701__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout290 team_08_WB.instance_to_wrap.allocation.game.cactus1size.state\[1\] vssd1
+ vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8945__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4640_ _0579_ _0597_ _0578_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6310_ net293 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__nor2_1
X_4571_ _0523_ _0539_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__and2_2
XFILLER_0_40_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7290_ net579 _2964_ _2966_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6241_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[19\]
+ _2193_ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7154__Y _2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9048__RESET_B net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6172_ _1879_ _2124_ _1878_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5123_ _0995_ _1072_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4794__X _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8707__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4954__B _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5054_ _1005_ _0998_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__and2b_1
X_8813_ net328 net187 vssd1 vssd1 vccd1 vccd1 _4291_ sky130_fd_sc_hd__or2_1
XANTENNA__8936__B2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8936__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout178_A _0674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4970__A _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5956_ _1860_ _1861_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_62_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8744_ _3775_ _4212_ net186 vssd1 vssd1 vccd1 vccd1 _4222_ sky130_fd_sc_hd__a21oi_1
X_4907_ _0738_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__nor2_4
X_5887_ _0715_ _0909_ _1791_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8675_ _4111_ _4149_ _4153_ vssd1 vssd1 vccd1 vccd1 _4154_ sky130_fd_sc_hd__and3_1
X_4838_ _0781_ _0790_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7626_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[9\]
+ net124 vssd1 vssd1 vccd1 vccd1 _3216_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4769_ _0719_ _0720_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__nor2_1
XANTENNA__4969__X _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7557_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr1\[0\] net549
+ _3164_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7488_ net301 _3047_ _3127_ _3124_ net302 vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__a311o_1
X_6508_ _2437_ _2438_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[5\]
+ sky130_fd_sc_hd__nor2_1
X_9227_ clknet_leaf_18_wb_clk_i _0055_ net230 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6439_ _0428_ _2385_ vssd1 vssd1 vccd1 vccd1 _2386_ sky130_fd_sc_hd__nor2_2
XFILLER_0_101_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9158_ clknet_leaf_37_wb_clk_i net544 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.cs
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8109_ net296 _3633_ _3634_ _3635_ vssd1 vssd1 vccd1 vccd1 _3637_ sky130_fd_sc_hd__a31o_1
Xhold21 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__9435__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9089_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[19\]
+ net222 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold10 _0252_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4864__B _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold43 _3169_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold98 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[7\]
+ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[4\] vssd1 vssd1
+ vccd1 vccd1 net585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8927__A1 _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5363__A_N _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5695__B _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8155__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8863__B1 _3271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6047__A _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7150__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5886__A _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5810_ _0924_ _1762_ _1761_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__o21a_1
XANTENNA__4790__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6790_ _2625_ _2626_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__nor2_1
XANTENNA__8262__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5741_ _1652_ _1653_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8460_ _3938_ _3940_ _3908_ vssd1 vssd1 vccd1 vccd1 _3941_ sky130_fd_sc_hd__a21oi_1
X_5672_ _1623_ _1624_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__xor2_1
XFILLER_0_72_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7354__B1 _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7411_ net307 _3041_ net304 vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__a21o_1
X_4623_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[4\] vssd1
+ vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__and2b_1
X_8391_ _3861_ _3871_ vssd1 vssd1 vccd1 vccd1 _3872_ sky130_fd_sc_hd__or2_2
XFILLER_0_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4554_ _0517_ _0522_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7342_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[19\]
+ _2996_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__and2_1
XANTENNA__4880__A_N _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7273_ net180 _2953_ _2955_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6224_ _1086_ _2152_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__xor2_1
XANTENNA__5126__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4485_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__inv_2
X_9012_ clknet_leaf_7_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[2\]
+ net212 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[2\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_55_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4965__A _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6155_ _2106_ _2107_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__or2_1
X_5106_ _1043_ _1057_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__nor2_1
X_6086_ net167 _0921_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5037_ _0958_ _0989_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6988_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2753_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8727_ net319 _4197_ vssd1 vssd1 vccd1 vccd1 _4205_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5939_ _1846_ _1889_ _1891_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8658_ net149 _4135_ _4136_ net136 vssd1 vssd1 vccd1 vccd1 _4137_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__7896__A1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7609_ _3182_ _3184_ vssd1 vssd1 vccd1 vccd1 _3199_ sky130_fd_sc_hd__and2_1
X_8589_ net155 _4067_ _4064_ net177 vssd1 vssd1 vccd1 vccd1 _4068_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_79_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4859__B _0602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__6320__B2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_101_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4882__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input23_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7584__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7887__B2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6311__A1 _2261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7960_ _2393_ _3481_ _3499_ net233 net588 vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__o32a_1
X_7891_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[18\]
+ _3441_ vssd1 vssd1 vccd1 vccd1 _3443_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4791__Y _0744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6911_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[7\]
+ _2704_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__a21oi_1
X_9630_ net483 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6842_ net528 _2658_ _2660_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__a21oi_1
X_9561_ net429 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
X_6773_ net274 _2615_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5724_ _0939_ _1617_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__xnor2_1
X_9492_ net367 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8720__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8512_ _3991_ vssd1 vssd1 vccd1 vccd1 _3992_ sky130_fd_sc_hd__inv_2
XANTENNA__7878__B2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5655_ _1557_ _1604_ _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9303__336 vssd1 vssd1 vccd1 vccd1 _9303__336/HI net336 sky130_fd_sc_hd__conb_1
X_8443_ _3290_ _3897_ vssd1 vssd1 vccd1 vccd1 _3924_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8374_ _3855_ _3856_ vssd1 vssd1 vccd1 vccd1 _3857_ sky130_fd_sc_hd__and2_1
X_4606_ _0423_ _0546_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5586_ _1527_ _1530_ _1537_ _1538_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_96_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7325_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[15\]
+ _2992_ vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4537_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[1\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__or2_1
XANTENNA__4966__Y _0919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7256_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[10\]
+ _2942_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__and2_1
X_4468_ net305 vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__inv_2
X_6207_ _2157_ _2159_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__xnor2_1
X_7187_ _2874_ _2894_ _2895_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__nor3_1
XANTENNA__4695__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8842__A3 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _2076_ _2077_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _2019_ _2021_ vssd1 vssd1 vccd1 vccd1 _2022_ sky130_fd_sc_hd__nor2_1
XANTENNA__7802__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8614__B _3178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6134__B _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4589__B _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8818__B1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8805__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8524__B net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8540__A _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5440_ _1345_ _1392_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4499__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5371_ net128 _1323_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8285__A1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8090_ _3617_ _3618_ vssd1 vssd1 vccd1 vccd1 _3619_ sky130_fd_sc_hd__nor2_1
X_7110_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[5\]
+ _2842_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[6\]
+ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_91_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7041_ _2787_ _2788_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__nor2_2
Xfanout108 net109 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_4
Xfanout119 net120 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_2
XFILLER_0_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8992_ clknet_leaf_2_wb_clk_i _0156_ net204 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7943_ _3464_ _3482_ vssd1 vssd1 vccd1 vccd1 _3483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7874_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[12\]
+ _3428_ net160 vssd1 vssd1 vccd1 vccd1 _3432_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout160_A _3403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9613_ net477 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
X_6825_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[7\]
+ _2648_ net275 vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9544_ net412 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
X_6756_ _2602_ _2603_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5707_ _0810_ _0812_ _0931_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5793__B _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9475_ net350 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_73_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6687_ _0464_ _2556_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5638_ _1590_ _1588_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout213_X net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8426_ net101 _3353_ _3280_ vssd1 vssd1 vccd1 vccd1 _3907_ sky130_fd_sc_hd__a21o_1
X_5569_ _1507_ _1519_ _1521_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4977__X _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8357_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[1\] team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3845_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_72_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold140 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7079__A2 _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8276__B2 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8276__A1 _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7308_ _2972_ _2976_ vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__nor2_1
Xhold162 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[15\] vssd1
+ vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[17\] vssd1 vssd1
+ vccd1 vccd1 net693 sky130_fd_sc_hd__dlygate4sd3_1
X_8288_ _2307_ net161 _2425_ net327 net225 vssd1 vssd1 vccd1 vccd1 _3782_ sky130_fd_sc_hd__o221a_1
Xhold173 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[18\] vssd1
+ vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__dlygate4sd3_1
X_7239_ net639 _2930_ net181 vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6145__A _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7423__B _3064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6450__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4940_ _0891_ _0892_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4871_ _0778_ _0822_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_19_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5894__A _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4553__D_N net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6610_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[17\] _2505_
+ _2478_ vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__o21ai_1
X_7590_ net184 net173 vssd1 vssd1 vccd1 vccd1 _3180_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6541_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[16\] _2457_
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[17\] vssd1 vssd1
+ vccd1 vccd1 _2460_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9260_ clknet_leaf_10_wb_clk_i _0082_ net227 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6472_ _2406_ _2409_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_41_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5423_ _0940_ _1323_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__xnor2_1
X_9191_ clknet_leaf_16_wb_clk_i _0021_ net227 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8211_ _2988_ _3720_ net121 vssd1 vssd1 vccd1 vccd1 _3721_ sky130_fd_sc_hd__a21o_1
X_5354_ _1304_ _1306_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__and2b_1
X_8142_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[1\]
+ net277 vssd1 vssd1 vccd1 vccd1 _3666_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5285_ _1233_ _1235_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nand2b_1
X_8073_ _0661_ _0702_ _2419_ _3603_ vssd1 vssd1 vccd1 vccd1 _3604_ sky130_fd_sc_hd__a22o_1
X_7024_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.wr team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.wr
+ net293 vssd1 vssd1 vccd1 vccd1 _2774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8975_ net311 vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__inv_2
X_7926_ net196 _3466_ vssd1 vssd1 vccd1 vccd1 _3467_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout163_X net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7857_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[7\]
+ _3416_ vssd1 vssd1 vccd1 vccd1 _3420_ sky130_fd_sc_hd__or2_1
X_6808_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ _2638_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__o21ba_1
XANTENNA__8194__B1 _2532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7788_ _2361_ _3374_ _2371_ _2359_ vssd1 vssd1 vccd1 vccd1 _3375_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6739_ net631 _2590_ net268 vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9527_ net402 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_18_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9458_ clknet_leaf_44_wb_clk_i _0396_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_dino
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8409_ net171 net94 _3888_ _3882_ vssd1 vssd1 vccd1 vccd1 _3890_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9389_ clknet_leaf_20_wb_clk_i _0336_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__8249__B2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_100_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_48_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7932__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5219__A _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _1021_ _1022_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7384__C_N team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5226__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8412__A1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5972_ _0761_ _0926_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8963__A2 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8760_ net313 _4235_ vssd1 vssd1 vccd1 vccd1 _4238_ sky130_fd_sc_hd__xor2_1
XANTENNA__7766__A3 _3355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4923_ _0852_ _0861_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7711_ _3286_ _3300_ vssd1 vssd1 vccd1 vccd1 _3301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8691_ _4165_ _4169_ vssd1 vssd1 vccd1 vccd1 _4170_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4854_ _0794_ _0801_ _0799_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__a21o_1
X_7642_ _3218_ _3223_ _3220_ vssd1 vssd1 vccd1 vccd1 _3232_ sky130_fd_sc_hd__a21oi_1
X_4785_ _0736_ _0737_ _0634_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__a21oi_4
X_7573_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.clk1
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr2\[0\] team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr2\[1\]
+ net257 vssd1 vssd1 vccd1 vccd1 _3173_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout123_A _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6524_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[11\] _2447_
+ vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__and2_1
X_9312_ clknet_leaf_2_wb_clk_i _0283_ net202 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.game.score\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9243_ clknet_leaf_19_wb_clk_i _0270_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.clk1
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6455_ _2374_ _2397_ vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__nor2_1
X_5406_ _1055_ _1311_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__and2_1
X_9174_ _0149_ _0411_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_6386_ team_08_WB.instance_to_wrap.allocation.game.game.score\[2\] _2326_ vssd1 vssd1
+ vccd1 vccd1 _2337_ sky130_fd_sc_hd__nor2_1
X_5337_ _1267_ _1287_ _1289_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__a21o_1
X_8125_ net299 _0652_ _3650_ _3651_ vssd1 vssd1 vccd1 vccd1 _3652_ sky130_fd_sc_hd__a31o_1
XANTENNA__8296__A_N net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5268_ _1218_ _1217_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__and2b_1
X_8056_ net314 net198 _3511_ _3590_ vssd1 vssd1 vccd1 vccd1 _3591_ sky130_fd_sc_hd__o211a_1
X_7007_ _2759_ _2763_ _2766_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__or3_1
XFILLER_0_98_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5199_ _1149_ _1151_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5217__A1 _1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4990__X _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8958_ _4433_ _4434_ vssd1 vssd1 vccd1 vccd1 _4435_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_84_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7909_ net561 _0713_ _2841_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8889_ _3873_ _4198_ _4365_ _4366_ vssd1 vssd1 vccd1 vccd1 _4367_ sky130_fd_sc_hd__or4_1
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7693__A2 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5045__Y _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7701__B net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5061__X _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[8\] vssd1
+ vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_2
Xfanout291 team_08_WB.instance_to_wrap.allocation.game.cactus1size.state\[1\] vssd1
+ vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8813__A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4570_ _0526_ _0529_ _0531_ _0533_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9520__395 vssd1 vssd1 vccd1 vccd1 _9520__395/HI net395 sky130_fd_sc_hd__conb_1
XFILLER_0_52_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4788__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6240_ _1642_ _2131_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7684__A2 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6171_ _1921_ _2123_ _1920_ vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_97_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5122_ _0919_ _0937_ _0935_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5412__A _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5053_ _0998_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8282__X _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8812_ _0422_ _0425_ vssd1 vssd1 vccd1 vccd1 _4290_ sky130_fd_sc_hd__nor2_1
XANTENNA__9387__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4970__B _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4958__B1 _0809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5955_ _1844_ _1887_ _1907_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_62_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8149__B1 _2393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8743_ _4213_ _4220_ vssd1 vssd1 vccd1 vccd1 _4221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4906_ _0634_ _0736_ _0737_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout240_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5886_ _0724_ _0905_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8674_ _4141_ _4146_ vssd1 vssd1 vccd1 vccd1 _4153_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4837_ _0602_ _0604_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__xnor2_4
XANTENNA__9327__Q team_08_WB.instance_to_wrap.allocation.game.controller.state\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7625_ _3210_ _3213_ vssd1 vssd1 vccd1 vccd1 _3215_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4768_ _0719_ _0720_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__and2_2
X_7556_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr1\[0\] _3163_
+ net257 vssd1 vssd1 vccd1 vccd1 _3164_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout126_X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4699_ net294 _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__nor2_1
X_7487_ _3126_ vssd1 vssd1 vccd1 vccd1 _3127_ sky130_fd_sc_hd__inv_2
X_6507_ net626 _2435_ _2429_ vssd1 vssd1 vccd1 vccd1 _2438_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9226_ clknet_leaf_20_wb_clk_i _0054_ net240 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6438_ net287 net285 vssd1 vssd1 vccd1 vccd1 _2385_ sky130_fd_sc_hd__nand2_2
X_9157_ clknet_leaf_36_wb_clk_i _0257_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.tft_sdi
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8108_ _3635_ vssd1 vssd1 vccd1 vccd1 _3636_ sky130_fd_sc_hd__inv_2
X_6369_ net287 _0648_ vssd1 vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__nand2_1
XANTENNA__5438__B2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__dlygate4sd3_1
X_9088_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[18\]
+ net222 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold11 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[6\]
+ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8617__B net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8039_ _3548_ _3552_ _3571_ _3574_ vssd1 vssd1 vccd1 vccd1 _3575_ sky130_fd_sc_hd__or4_1
Xhold44 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[2\]
+ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[4\]
+ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 _0180_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold88 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.wr vssd1
+ vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[0\]
+ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[2\] vssd1 vssd1
+ vccd1 vccd1 net597 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8927__A2 _3179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9463__338 vssd1 vssd1 vccd1 vccd1 _9463__338/HI net338 sky130_fd_sc_hd__conb_1
XFILLER_0_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9504__379 vssd1 vssd1 vccd1 vccd1 _9504__379/HI net379 sky130_fd_sc_hd__conb_1
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7666__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6874__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7712__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8527__B _3241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6047__B _0926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8918__A2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4790__B _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5886__B _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5740_ _1692_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5671_ _0940_ _1571_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7410_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[2\]
+ _3042_ _3054_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_26_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4789__Y _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4622_ _0578_ _0579_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__nand2b_2
X_8390_ net171 _3868_ vssd1 vssd1 vccd1 vccd1 _3871_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4553_ net326 _0518_ _0521_ net329 vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__or4b_4
XFILLER_0_5_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7341_ _2995_ _3005_ net122 vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__a21oi_1
X_4484_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.drawDoneCactus vssd1
+ vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7272_ _2954_ vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6223_ _2153_ _2175_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9011_ clknet_leaf_8_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[1\]
+ net223 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8718__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4965__B _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6154_ _2098_ _2099_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__xor2_1
X_5105_ _1043_ _1057_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__and2_1
X_6085_ _1959_ _2034_ _2037_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__and3_1
X_5036_ _0987_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6987_ _0461_ _2752_ _0019_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__a21oi_1
X_5938_ _0754_ _0929_ _0931_ _0761_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__o22a_1
XANTENNA__7069__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8726_ net100 _4200_ vssd1 vssd1 vccd1 vccd1 _4204_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5869_ _1819_ _1821_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__and2b_1
X_8657_ net284 _3679_ _0640_ _2388_ vssd1 vssd1 vccd1 vccd1 _4136_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7608_ _3183_ _3196_ _3197_ vssd1 vssd1 vccd1 vccd1 _3198_ sky130_fd_sc_hd__and3_1
X_8588_ _4063_ _4066_ vssd1 vssd1 vccd1 vccd1 _4067_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_79_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7539_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[5\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[7\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[1\] vssd1
+ vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__mux4_1
XANTENNA__5317__A _1038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9209_ clknet_leaf_23_wb_clk_i _0264_ _0151_ vssd1 vssd1 vccd1 vccd1 team_08_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_1
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__7091__X _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4882__A2 _0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8073__A2 _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7820__A2 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8363__A team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9545__413 vssd1 vssd1 vccd1 vccd1 _9545__413/HI net413 sky130_fd_sc_hd__conb_1
XFILLER_0_98_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5898__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9591__455 vssd1 vssd1 vccd1 vccd1 _9591__455/HI net455 sky130_fd_sc_hd__conb_1
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8538__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7811__A2 _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7890_ _3441_ _3442_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[17\]
+ net166 vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__a2bb2o_1
X_9485__360 vssd1 vssd1 vccd1 vccd1 _9485__360/HI net360 sky130_fd_sc_hd__conb_1
X_6910_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[7\]
+ _2704_ _2706_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6841_ net528 _2658_ net271 vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__o21ai_1
X_9560_ net428 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_9_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6772_ _0465_ _2613_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8511_ _3280_ _3961_ _3990_ _3988_ _3966_ vssd1 vssd1 vccd1 vccd1 _3991_ sky130_fd_sc_hd__o32a_1
X_5723_ _1659_ _1675_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9491_ net366 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XANTENNA__8720__B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5654_ net141 _0906_ _1606_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8442_ _3330_ _3875_ vssd1 vssd1 vccd1 vccd1 _3923_ sky130_fd_sc_hd__nor2_1
X_8373_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] net289 _3471_
+ team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1 vssd1 vccd1
+ vccd1 _3856_ sky130_fd_sc_hd__o31ai_1
X_4605_ net326 _0540_ _0564_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[3\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5585_ _1481_ _1536_ _1535_ _1505_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_96_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5137__A _1087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8288__C1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8827__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7324_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[14\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[13\]
+ _2991_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4536_ net317 team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1
+ vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__xor2_4
XANTENNA_fanout203_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4467_ net307 vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__inv_2
XANTENNA__9032__RESET_B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7255_ net179 _2941_ _2943_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__and3_1
X_6206_ _1194_ _2158_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_74_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7186_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[11\] _2892_ vssd1
+ vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__nor2_1
XANTENNA_input8_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6137_ _2087_ _2089_ _2086_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_5_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _1978_ _2020_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__nand2_1
X_5019_ _0748_ _0971_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8183__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7086__X _2828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8630__B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8709_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\] _3241_ vssd1
+ vssd1 vccd1 vccd1 _4188_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8077__B team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9469__344 vssd1 vssd1 vccd1 vccd1 _9469__344/HI net344 sky130_fd_sc_hd__conb_1
XANTENNA__8805__B _3266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7156__B net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5370_ _1319_ _1321_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7040_ _0457_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\] vssd1
+ vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__or3_2
XFILLER_0_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout109 _3242_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_52_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8991_ clknet_leaf_1_wb_clk_i _0155_ net211 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7942_ _0421_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[1\] vssd1
+ vssd1 vccd1 vccd1 _3482_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6235__B _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9612_ net476 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
X_7873_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[12\]
+ _3428_ vssd1 vssd1 vccd1 vccd1 _3431_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6824_ _2648_ _2649_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout153_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6755_ net611 _2601_ net268 vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9543_ net411 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5706_ _1645_ _1657_ _1658_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__o21ai_2
XANTENNA__9284__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout320_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9474_ net349 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_66_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6686_ net270 _2553_ _2556_ _2557_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__and4_1
XANTENNA__7066__B _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8425_ net154 net94 _3903_ _3905_ vssd1 vssd1 vccd1 vccd1 _3906_ sky130_fd_sc_hd__o211a_1
X_5637_ _1539_ _1589_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_76_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9213__RESET_B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5568_ _1469_ _1520_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout206_X net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8356_ _3844_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4519_ _0484_ _0486_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__nand2_1
X_8287_ _0422_ net193 _3511_ _3780_ vssd1 vssd1 vccd1 vccd1 _3781_ sky130_fd_sc_hd__o211a_1
Xhold130 team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[1\] vssd1 vssd1
+ vccd1 vccd1 net628 sky130_fd_sc_hd__dlygate4sd3_1
X_7307_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[1\] _2975_ _2978_
+ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold152 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[2\] vssd1
+ vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold141 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _1450_ _1451_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_72_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold174 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.clk1
+ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[15\] vssd1
+ vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[9\]
+ vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__dlygate4sd3_1
X_7238_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[4\]
+ _2930_ vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__and2_1
Xhold196 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.clk1
+ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__dlygate4sd3_1
X_7169_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[4\] _2881_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6145__B _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9159__D _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8641__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7720__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6450__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4870_ _0738_ net148 _0822_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6202__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5894__B _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6540_ net572 _2457_ _2459_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[16\]
+ sky130_fd_sc_hd__a21oi_1
X_9597__461 vssd1 vssd1 vccd1 vccd1 _9597__461/HI net461 sky130_fd_sc_hd__conb_1
XFILLER_0_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6471_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[6\]
+ _2413_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_41_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5422_ net128 _1374_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__nand2_1
X_9190_ clknet_leaf_19_wb_clk_i _0259_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.clk1
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8210_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[7\]
+ _2987_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[8\]
+ vssd1 vssd1 vccd1 vccd1 _3720_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5353_ _1303_ _1305_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__nor2_1
X_8141_ _2384_ _3462_ _3665_ net238 net564 vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__o32a_1
XANTENNA__5415__A _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5284_ _1228_ _1231_ _1229_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8072_ _0704_ _3602_ vssd1 vssd1 vccd1 vccd1 _3603_ sky130_fd_sc_hd__nand2_1
XANTENNA__8726__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7023_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.tft_reset net3 vssd1
+ vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8966__B1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout270_A _2548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8974_ net311 vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7925_ net335 net333 vssd1 vssd1 vccd1 vccd1 _3466_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7856_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[7\]
+ _3416_ vssd1 vssd1 vccd1 vccd1 _3419_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6807_ _2635_ _2636_ _2637_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_65_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4999_ _0876_ _0877_ _0879_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__o21a_1
X_9526_ net401 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
X_7787_ _3372_ _3373_ _2375_ vssd1 vssd1 vccd1 vccd1 _3374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6738_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[6\]
+ _2588_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9457_ clknet_leaf_1_wb_clk_i _0395_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_cloud
+ sky130_fd_sc_hd__dfxtp_1
X_6669_ net580 _0443_ vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__nor2_2
XANTENNA__8497__A2 _3976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9388_ clknet_leaf_29_wb_clk_i _0335_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__7805__A _2972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8408_ net171 net94 _3888_ _3882_ vssd1 vssd1 vccd1 vccd1 _3889_ sky130_fd_sc_hd__a31oi_1
XANTENNA__5180__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8339_ _3576_ _3813_ _3827_ vssd1 vssd1 vccd1 vccd1 _3829_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5325__A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5060__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5235__A _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5241__Y _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8658__A1_N net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5971_ _0724_ _0929_ _1889_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__or3b_1
X_9525__400 vssd1 vssd1 vccd1 vccd1 _9525__400/HI net400 sky130_fd_sc_hd__conb_1
XFILLER_0_87_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4922_ net138 _0852_ _0815_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_75_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8281__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8690_ net119 _3608_ _4168_ vssd1 vssd1 vccd1 vccd1 _4169_ sky130_fd_sc_hd__a21o_1
X_7710_ net110 net108 vssd1 vssd1 vccd1 vccd1 _3300_ sky130_fd_sc_hd__nand2_2
XFILLER_0_87_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7641_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[7\]
+ _3229_ _3230_ vssd1 vssd1 vccd1 vccd1 _3231_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_23_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4853_ _0749_ _0803_ _0804_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7572_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.clk1
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr2\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3172_ sky130_fd_sc_hd__a21oi_1
X_4784_ _0631_ _0633_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6523_ _2447_ _2448_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[10\]
+ sky130_fd_sc_hd__nor2_1
X_9311_ clknet_leaf_0_wb_clk_i _0282_ net201 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.game.score\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9242_ clknet_leaf_20_wb_clk_i _0269_ net239 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr2\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_15_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6454_ _0419_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\]
+ net259 _2398_ _2396_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a221o_1
X_5405_ _1014_ _1357_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload50 clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5145__A _0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9173_ _0148_ _0410_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_6385_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.col net256 _2324_
+ vssd1 vssd1 vccd1 vccd1 _2336_ sky130_fd_sc_hd__or3b_2
X_5336_ _1213_ _1232_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__xnor2_1
X_8124_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\] _3647_ _3648_
+ _3649_ net278 vssd1 vssd1 vccd1 vccd1 _3651_ sky130_fd_sc_hd__a221o_1
X_5267_ net138 _1215_ _1219_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__a21o_1
X_8055_ _3587_ _3588_ _3589_ vssd1 vssd1 vccd1 vccd1 _3590_ sky130_fd_sc_hd__o21ai_1
X_7006_ _0468_ _2756_ vssd1 vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__nor2_1
X_5198_ _0856_ _1150_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8957_ _0426_ net109 _4187_ _4191_ _4185_ vssd1 vssd1 vccd1 vccd1 _4434_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_84_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7908_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[2\]
+ _0402_ _3453_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__or3b_1
XFILLER_0_39_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8888_ _3888_ _3895_ _3870_ vssd1 vssd1 vccd1 vccd1 _4366_ sky130_fd_sc_hd__a21oi_1
X_7839_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[1\] team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _3407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6431__A1_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload0 clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__inv_6
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9509_ net384 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_33_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8366__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout270 _2548_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
Xfanout292 team_08_WB.instance_to_wrap.allocation.game.cactus1size.state\[0\] vssd1
+ vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8813__B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9433__Q team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6170_ _2121_ _2122_ _1956_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5121_ _0919_ _0937_ _0935_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__o21a_2
XFILLER_0_97_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5052_ _1003_ _1004_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__nor2_1
XANTENNA__5412__B _1215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8811_ net320 net101 vssd1 vssd1 vccd1 vccd1 _4289_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4958__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8742_ _4214_ _4218_ _4215_ vssd1 vssd1 vccd1 vccd1 _4220_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_87_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5954_ _1903_ _1904_ _1906_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_62_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4905_ _0851_ _0855_ _0857_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__a21oi_1
X_5885_ net182 _0910_ _1791_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_62_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8673_ _4120_ _4133_ _4137_ _4139_ _4151_ vssd1 vssd1 vccd1 vccd1 _4152_ sky130_fd_sc_hd__o221a_1
X_4836_ _0787_ _0788_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__nand2_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7624_ _3210_ _3213_ vssd1 vssd1 vccd1 vccd1 _3214_ sky130_fd_sc_hd__nor2_2
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7555_ net548 team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4979__A _0809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4767_ _0587_ _0592_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__xnor2_1
XANTENNA__6580__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6506_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[4\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[5\]
+ _2433_ vssd1 vssd1 vccd1 vccd1 _2437_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4698_ net299 _0653_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__nand2_4
X_7486_ _3125_ _3050_ _3043_ _3116_ vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__a2bb2o_1
X_9225_ clknet_leaf_21_wb_clk_i _0049_ net240 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6437_ _0430_ _0653_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__nor2_1
X_6368_ _2318_ _2319_ _2315_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__o21ai_1
XANTENNA__8609__C1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9156_ clknet_leaf_37_wb_clk_i _0256_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.tft_dc
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5319_ _1038_ _1222_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__a21bo_1
X_8107_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[0\] net277 vssd1
+ vssd1 vccd1 vccd1 _3635_ sky130_fd_sc_hd__or2_2
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6299_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[16\]
+ _2200_ _2203_ _2251_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9087_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[17\]
+ net222 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold23 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[4\] vssd1
+ vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 _0245_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__dlygate4sd3_1
X_8038_ _3572_ _3573_ vssd1 vssd1 vccd1 vccd1 _3574_ sky130_fd_sc_hd__nor2_1
Xhold56 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[2\]
+ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.cs vssd1 vssd1
+ vccd1 vccd1 net543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold89 _0068_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_08_WB.instance_to_wrap.allocation.game.controller.color\[10\] vssd1 vssd1
+ vccd1 vccd1 net565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 team_08_WB.instance_to_wrap.allocation.game.cactusMove.cactusMovement vssd1
+ vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7060__A1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8633__B _3241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6571__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7712__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5513__A _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8824__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5670_ _1620_ _1622_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_4621_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[5\] vssd1
+ vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4552_ net320 net317 vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__nand2_1
X_7340_ net546 _2994_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8303__B2 _3527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7271_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[15\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[14\]
+ _2950_ vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__and3_1
X_4483_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__inv_2
X_6222_ _2154_ _2174_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9010_ clknet_leaf_7_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[0\]
+ net212 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__7511__C1 _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5423__A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6153_ _2103_ _2105_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_55_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5104_ _1015_ _1056_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__xnor2_1
X_6084_ _2002_ _2036_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__nor2_1
X_5035_ _0897_ _0899_ _0986_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__and3_1
XANTENNA__8734__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_69_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6986_ _2417_ _2751_ _2752_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5937_ _0772_ _0927_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__nand2_1
X_8725_ net100 _4200_ _4202_ net97 vssd1 vssd1 vccd1 vccd1 _4203_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8656_ _4133_ _4134_ vssd1 vssd1 vccd1 vccd1 _4135_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5868_ _1050_ _1820_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout236_X net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7607_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[12\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\] net176
+ _3177_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\]
+ vssd1 vssd1 vccd1 vccd1 _3197_ sky130_fd_sc_hd__a32o_1
X_5799_ _1700_ _1701_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__xor2_1
X_4819_ _0760_ _0770_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__xor2_4
XFILLER_0_44_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8587_ _0686_ _4062_ net163 vssd1 vssd1 vccd1 vccd1 _4066_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_28_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7538_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[1\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[3\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[1\] vssd1
+ vssd1 vccd1 vccd1 _3154_ sky130_fd_sc_hd__mux4_1
XANTENNA__6305__B1 _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7469_ _3107_ _3110_ net115 vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__or3b_1
X_9208_ clknet_leaf_10_wb_clk_i _0263_ net229 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr2\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__7502__C1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__4867__A0 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__8058__B1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7024__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9139_ clknet_leaf_39_wb_clk_i _0240_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5508__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8049__B1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9331__RESET_B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6840_ _2658_ _2659_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__nor2_1
X_6771_ _2611_ _2613_ _2614_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5722_ _1659_ _1673_ _1674_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__nand3_1
XANTENNA__6783__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8510_ _3981_ _3989_ _3977_ vssd1 vssd1 vccd1 vccd1 _3990_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_58_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8720__C net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9490_ net365 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_73_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5653_ _1557_ _1604_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__xor2_1
X_8441_ _3355_ _3921_ vssd1 vssd1 vccd1 vccd1 _3922_ sky130_fd_sc_hd__or2_1
X_5584_ _1505_ _1535_ _1536_ _1481_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_72_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8372_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\]
+ net289 _3471_ vssd1 vssd1 vccd1 vccd1 _3855_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4604_ net326 _0564_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5137__B _1088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4535_ net319 team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] _0503_
+ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__a21o_1
X_7323_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[12\]
+ _2990_ vssd1 vssd1 vccd1 vccd1 _2991_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__8827__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4466_ net301 vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__inv_2
X_7254_ _2942_ vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__inv_2
XANTENNA__5510__A1 _0814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6205_ net144 _0812_ _0875_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_74_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7185_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[10\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[11\]
+ _2891_ vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__and3_1
X_6136_ _2086_ _2088_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9072__RESET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _1975_ _1977_ vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout186_X net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5018_ _0969_ _0970_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ _2741_ net158 _2740_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__and3b_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8708_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\] net113 vssd1
+ vssd1 vccd1 vccd1 _4187_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8639_ _2538_ _4117_ vssd1 vssd1 vccd1 vccd1 _4118_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5047__B _0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8818__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout99_X net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5063__A _1011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6446__X _2393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8268__B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8990_ clknet_leaf_2_wb_clk_i _0154_ net211 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7941_ _0702_ _3479_ vssd1 vssd1 vccd1 vccd1 _3481_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7872_ _3428_ _3430_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[11\]
+ net165 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a2bb2o_1
X_9611_ net475 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_93_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6823_ net655 _2646_ net271 vssd1 vssd1 vccd1 vccd1 _2649_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_34_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9542_ net410 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
X_6754_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[12\]
+ _2601_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_98_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5705_ _1611_ _1612_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9473_ net348 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
X_6685_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5636_ _1537_ _1538_ _1527_ _1530_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8424_ net154 _3904_ _3323_ vssd1 vssd1 vccd1 vccd1 _3905_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_76_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout313_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4987__A _0939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5567_ _1460_ _1467_ _1468_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__and3_1
X_8355_ _3843_ _2874_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5498_ _1397_ _1398_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold142 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _0484_ _0486_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__and2_2
X_8286_ _3502_ _3509_ net196 vssd1 vssd1 vccd1 vccd1 _3780_ sky130_fd_sc_hd__a21o_1
X_7306_ _0449_ _2974_ _2979_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__o21ai_1
Xhold153 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[18\] vssd1
+ vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout101_X net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ net324 vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__inv_2
X_7237_ net179 _2929_ _2931_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__and3_1
X_7168_ net585 _2881_ _2883_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__a21oi_1
X_6119_ _1959_ _2034_ _2071_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__a21oi_1
X_7099_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[21\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[20\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[19\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[18\]
+ vssd1 vssd1 vccd1 vccd1 _2838_ sky130_fd_sc_hd__or4_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6747__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8641__B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9452__SET_B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5058__A _0825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5505__B _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5521__A _0939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6470_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[16\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[15\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[9\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_41_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5421_ _1372_ _1373_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__and2_2
X_5352_ _1011_ _0999_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8140_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\] _3664_ net137
+ vssd1 vssd1 vccd1 vccd1 _3665_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8071_ _0661_ _0703_ vssd1 vssd1 vccd1 vccd1 _3602_ sky130_fd_sc_hd__or2_1
X_5283_ _1235_ _1233_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__nand2b_1
X_7022_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[6\] team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[3\]
+ _2771_ _0459_ _0460_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__o311a_1
X_9534__490 vssd1 vssd1 vccd1 vccd1 net490 _9534__490/LO sky130_fd_sc_hd__conb_1
XANTENNA__7218__A1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoMovement
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8415__B1 _3895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8966__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8973_ net311 vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__inv_2
X_7924_ _0491_ _0549_ net193 vssd1 vssd1 vccd1 vccd1 _3465_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout263_A _0514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7855_ net159 _3417_ _3418_ net165 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__a32o_1
X_6806_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_65_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4998_ _0903_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9525_ net400 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_19_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7786_ _2373_ _2378_ vssd1 vssd1 vccd1 vccd1 _3373_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout149_X net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6737_ _2590_ _2591_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6668_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.idle
+ vssd1 vssd1 vccd1 vccd1 _2544_ sky130_fd_sc_hd__nand2b_2
X_9456_ clknet_leaf_51_wb_clk_i _0394_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_over
+ sky130_fd_sc_hd__dfxtp_1
X_5619_ net128 _1571_ _1569_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__a21o_1
X_9387_ clknet_leaf_29_wb_clk_i _0334_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__8189__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6599_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[13\] _2498_
+ _2500_ _2478_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[13\]
+ sky130_fd_sc_hd__o211a_1
X_8407_ _3314_ _3360_ vssd1 vssd1 vccd1 vccd1 _3888_ sky130_fd_sc_hd__nor2_4
XANTENNA__7093__A team_08_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5606__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8338_ _3576_ _3813_ _3827_ vssd1 vssd1 vccd1 vccd1 _3828_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7821__A team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8269_ net330 _2268_ vssd1 vssd1 vccd1 vccd1 _3764_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5059__Y _1012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7932__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7715__B net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7731__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4793__C _0744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5970_ net140 _0917_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_32_Left_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4921_ _0845_ _0873_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4852_ _0803_ _0804_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7640_ _3217_ _3227_ vssd1 vssd1 vccd1 vccd1 _3230_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4783_ _0734_ _0735_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__and2b_4
X_7571_ net257 _3171_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6522_ net658 _2445_ net156 vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9310_ clknet_leaf_0_wb_clk_i _0281_ net200 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.game.score\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9241_ clknet_leaf_20_wb_clk_i _0268_ net239 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr2\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_41_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6453_ _2383_ _2397_ vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__and2b_1
X_5404_ _1356_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload40 clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_8
XANTENNA_clkload48_A clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload51 clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__inv_6
XFILLER_0_42_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9172_ _0147_ _0409_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_8123_ net282 _0646_ vssd1 vssd1 vccd1 vccd1 _3650_ sky130_fd_sc_hd__nand2_1
X_6384_ _2331_ _2332_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.slow_clk
+ vssd1 vssd1 vccd1 vccd1 _2335_ sky130_fd_sc_hd__o21ai_4
X_5335_ _1267_ _1287_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__nand2_1
XANTENNA__8296__X _3789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5266_ _1217_ _1218_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__and2b_1
X_8054_ _3587_ _3588_ net195 vssd1 vssd1 vccd1 vccd1 _3589_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7005_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] _2756_ _2765_ vssd1
+ vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5197_ _0794_ _0798_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_50_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8956_ net287 _3214_ net119 _0427_ vssd1 vssd1 vccd1 vccd1 _4433_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_84_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7907_ _2776_ _2785_ _2840_ vssd1 vssd1 vccd1 vccd1 _3453_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8887_ _4278_ _4358_ _4364_ _4284_ vssd1 vssd1 vccd1 vccd1 _4365_ sky130_fd_sc_hd__o211a_1
XANTENNA__4505__A net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7838_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[1\] team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _3406_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9110__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7769_ net149 net133 vssd1 vssd1 vccd1 vccd1 _3359_ sky130_fd_sc_hd__nor2_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload1 clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_19_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9508_ net383 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_73_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9439_ clknet_leaf_28_wb_clk_i _0384_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__8875__B1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6350__B2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6350__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout271 _2548_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
Xfanout282 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[7\] vssd1
+ vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout293 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.init_done
+ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5120_ _1072_ _0995_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5051_ _1001_ _1002_ _0999_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_88_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8810_ _4251_ _4287_ _4256_ vssd1 vssd1 vccd1 vccd1 _4288_ sky130_fd_sc_hd__o21ai_1
X_8741_ _4214_ _4215_ vssd1 vssd1 vccd1 vccd1 _4219_ sky130_fd_sc_hd__or2_1
XANTENNA__4958__A2 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5953_ _1844_ _1905_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_62_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8149__A2 _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4904_ _0738_ _0811_ _0856_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__a21oi_1
X_5884_ _1792_ _1794_ _1793_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9097__RESET_B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8672_ _4148_ _4149_ _4150_ _4141_ vssd1 vssd1 vccd1 vccd1 _4151_ sky130_fd_sc_hd__a31o_1
X_4835_ net148 _0783_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7623_ _3206_ _3212_ _3195_ vssd1 vssd1 vccd1 vccd1 _3213_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_16_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7554_ net548 _2638_ _3015_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__mux2_1
X_4766_ _0714_ _0590_ _0591_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__mux2_2
XFILLER_0_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout226_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6505_ _2435_ _2436_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4697_ net280 _0646_ _0651_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__or3_2
X_7485_ _3084_ _3071_ vssd1 vssd1 vccd1 vccd1 _3125_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9224_ clknet_leaf_19_wb_clk_i _0265_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.clk1
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6332__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6436_ net259 _2360_ _2383_ _2325_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4995__A _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6367_ _2317_ _2304_ _2302_ _2299_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__8609__B1 _3271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9155_ clknet_leaf_37_wb_clk_i _0105_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.idle
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5318_ _1220_ _1270_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8106_ net287 _0642_ net284 vssd1 vssd1 vccd1 vccd1 _3634_ sky130_fd_sc_hd__a21o_1
X_6298_ _0447_ _2202_ _2205_ _2250_ vssd1 vssd1 vccd1 vccd1 _2251_ sky130_fd_sc_hd__a211o_1
X_9086_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[16\]
+ net222 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold13 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[5\]
+ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _1048_ _1201_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__or2_1
X_8037_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] _3561_ vssd1
+ vssd1 vccd1 vccd1 _3573_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_2_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold35 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[31\] vssd1 vssd1
+ vccd1 vccd1 net533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[6\] vssd1
+ vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 _0258_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 _0117_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7060__A2 _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8939_ _2296_ _3276_ _4414_ _2301_ _4415_ vssd1 vssd1 vccd1 vccd1 _4416_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_14_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8383__Y _3864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8824__B net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4620_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[5\] vssd1
+ vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7455__A_N _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9444__Q team_08_WB.instance_to_wrap.allocation.game.controller.v\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8303__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8839__B1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4551_ net319 net316 vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__and2_2
XFILLER_0_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7270_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[14\]
+ _2950_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__a21o_1
X_4482_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6221_ _2155_ _2173_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_38_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _2098_ _2104_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_55_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8718__C _4196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5103_ _1047_ _1054_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6083_ _1999_ _2001_ _2000_ vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__a21oi_1
X_5034_ _0897_ _0899_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9278__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout176_A _3178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9207__RESET_B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6985_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[23\]
+ _2750_ vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5936_ net167 _0931_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__nor2_1
XANTENNA__7918__X _3460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8750__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8724_ _0520_ _4197_ _4201_ vssd1 vssd1 vccd1 vccd1 _4202_ sky130_fd_sc_hd__a21o_1
X_8655_ net284 _3679_ net281 vssd1 vssd1 vccd1 vccd1 _4134_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout131_X net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5867_ _0761_ _0859_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__nand2b_1
X_7606_ _3188_ _3194_ vssd1 vssd1 vccd1 vccd1 _3196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5798_ _1750_ _1749_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__nand2b_1
X_4818_ _0760_ _0770_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8586_ net177 _4064_ vssd1 vssd1 vccd1 vccd1 _4065_ sky130_fd_sc_hd__or2_1
XANTENNA__7750__B1 _3280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7537_ net513 net507 _2545_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__mux2_1
X_4749_ _0661_ _0703_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7468_ _3067_ _3108_ vssd1 vssd1 vccd1 vccd1 _3110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9207_ clknet_leaf_19_wb_clk_i _0262_ net230 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr2\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__7372__Y _3022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6419_ _2369_ team_08_WB.instance_to_wrap.allocation.game.game.score\[2\] _2336_
+ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__mux2_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
X_7399_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[2\]
+ net308 vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__nor2_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
X_9138_ clknet_leaf_38_wb_clk_i _0239_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_9069_ clknet_leaf_9_wb_clk_i _0204_ net225 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_9510__385 vssd1 vssd1 vccd1 vccd1 _9510__385/HI net385 sky130_fd_sc_hd__conb_1
XANTENNA__6445__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7975__S net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5508__B _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8049__A1 _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8835__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9371__RESET_B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9300__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6770_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__a21o_1
X_5721_ _1645_ _1657_ _1658_ vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5652_ net141 _0906_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8440_ _3273_ _3281_ vssd1 vssd1 vccd1 vccd1 _3921_ sky130_fd_sc_hd__nand2_1
X_5583_ _1479_ _1480_ _1456_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8371_ _3854_ _3843_ _2875_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__a2bb2o_1
X_4603_ _0540_ _0563_ net256 vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_96_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4534_ _0483_ _0502_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__and2_1
XANTENNA__9321__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8288__B2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7322_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[10\]
+ _2989_ vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__or3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4465_ net303 vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__inv_2
X_7253_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[8\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[9\]
+ _2938_ vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__and3_1
XANTENNA__5510__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6204_ _1047_ _1054_ _1052_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_74_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7184_ net610 _2891_ _2893_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6135_ _2073_ _2085_ _2084_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_5_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _2018_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5017_ _0968_ _0798_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__and2b_1
XFILLER_0_68_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6968_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[17\]
+ _2738_ vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_37_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8707_ net107 _4114_ _4185_ vssd1 vssd1 vccd1 vccd1 _4186_ sky130_fd_sc_hd__and3_1
X_5919_ _1871_ _1870_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4785__B1 _0634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6899_ _2698_ _2699_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7723__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8638_ net283 net135 vssd1 vssd1 vccd1 vccd1 _4117_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8569_ net152 _4044_ _4047_ vssd1 vssd1 vccd1 vccd1 _4048_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5063__B _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_97_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8565__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7940_ net139 net137 vssd1 vssd1 vccd1 vccd1 _3480_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7871_ net160 _3429_ vssd1 vssd1 vccd1 vccd1 _3430_ sky130_fd_sc_hd__nand2_1
X_9610_ net474 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_89_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6822_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[6\]
+ _2644_ vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__and3_1
XANTENNA__6372__X _2324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9541_ net409 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
X_6753_ net272 _2600_ _2601_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__nor3_1
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9472_ net347 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
X_5704_ _1656_ _1655_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__and2b_1
X_6684_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__nand3_1
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5635_ _1585_ _1587_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8423_ net135 net112 _3302_ vssd1 vssd1 vccd1 vccd1 _3904_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5566_ _1518_ _1517_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__nand2b_1
X_8354_ _0561_ _3842_ vssd1 vssd1 vccd1 vccd1 _3843_ sky130_fd_sc_hd__or2_2
Xhold110 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[7\]
+ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__dlygate4sd3_1
X_5497_ _0745_ _0836_ _1449_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__o21ai_2
Xhold121 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ net326 team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__or2_1
X_8285_ net170 _3774_ _3778_ net297 vssd1 vssd1 vccd1 vccd1 _3779_ sky130_fd_sc_hd__o31a_1
XANTENNA__7363__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7305_ _2976_ _2978_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__nand2_1
Xhold143 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[1\] vssd1
+ vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5164__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold165 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ net326 vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__inv_2
X_7236_ _2930_ vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__inv_2
Xhold154 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[30\] vssd1
+ vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[6\]
+ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7167_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[4\] _2881_ _0523_
+ vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5247__A1 _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9222__RESET_B net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6118_ _0717_ _0926_ _0931_ net182 vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__o22a_1
X_7098_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[0\]
+ _0435_ _2776_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__or3_1
XANTENNA__8433__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4508__A _0473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6049_ _1999_ _2000_ _2001_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__and3_1
X_9581__445 vssd1 vssd1 vccd1 vccd1 _9581__445/HI net445 sky130_fd_sc_hd__conb_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5960__A2_N _1912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9475__350 vssd1 vssd1 vccd1 vccd1 _9475__350/HI net350 sky130_fd_sc_hd__conb_1
XFILLER_0_60_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9516__391 vssd1 vssd1 vccd1 vccd1 _9516__391/HI net391 sky130_fd_sc_hd__conb_1
XANTENNA__5802__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7720__C _3305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8424__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5249__A _1048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4512__A_N net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5420_ _1364_ _1369_ _1371_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__nand3_1
XFILLER_0_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5351_ _0863_ net138 _1000_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5282_ _1175_ _1234_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8070_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\] net161 _2534_
+ net299 vssd1 vssd1 vccd1 vccd1 _3601_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4662__A_N team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7021_ _0460_ _2768_ _2771_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[1\]
+ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__a31o_1
XFILLER_0_10_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8966__A2 _3276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8972_ net311 vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__inv_2
X_7923_ _0491_ _0549_ vssd1 vssd1 vccd1 vccd1 _3464_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7854_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[6\]
+ _3413_ vssd1 vssd1 vccd1 vccd1 _3418_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4615__X _0573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_A _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6805_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[9\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_65_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7785_ _2371_ _3371_ vssd1 vssd1 vccd1 vccd1 _3372_ sky130_fd_sc_hd__xnor2_1
X_4997_ _0948_ _0949_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__nand2_1
X_6736_ net682 _2588_ net268 vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__o21ai_1
X_9524_ net399 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7645__Y _3235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6667_ net279 _2543_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[8\]
+ sky130_fd_sc_hd__xnor2_1
X_9455_ clknet_leaf_0_wb_clk_i _0393_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_idle
+ sky130_fd_sc_hd__dfxtp_1
X_5618_ _1569_ _1570_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__nor2_1
X_9386_ clknet_leaf_9_wb_clk_i _0333_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6598_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[13\] _2498_
+ vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8406_ net116 net112 _3868_ net172 vssd1 vssd1 vccd1 vccd1 _3887_ sky130_fd_sc_hd__o211a_1
X_5549_ net143 _1501_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__nand2_1
XANTENNA__5606__B _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8337_ _3588_ _0570_ _3572_ vssd1 vssd1 vccd1 vccd1 _3827_ sky130_fd_sc_hd__mux2_1
X_8268_ net332 net329 vssd1 vssd1 vccd1 vccd1 _3763_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5622__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7219_ _0423_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__xnor2_1
X_8199_ _2984_ _3710_ _3713_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8406__A1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8957__A2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4701__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8099__B _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7731__B net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4682__A2 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoMovement
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7081__B1 _2823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4920_ _0871_ _0872_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__nor2_1
X_4851_ _0802_ _0786_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6187__A2 _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8581__B1 _4036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4782_ _0609_ _0630_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__xnor2_1
X_7570_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr1\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr1\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.clk1 vssd1
+ vssd1 vccd1 vccd1 _3171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6521_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[9\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[10\]
+ _2443_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9240_ clknet_leaf_19_wb_clk_i _0267_ net230 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr1\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4611__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8884__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6452_ _2362_ _2376_ _2364_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__o21ai_1
X_5403_ _1353_ _1354_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__xor2_1
Xclkload41 clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__inv_8
XFILLER_0_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9171_ _0146_ _0408_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload30 clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8122_ _0428_ _3633_ net296 vssd1 vssd1 vccd1 vccd1 _3649_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6383_ _2331_ _2332_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.slow_clk
+ vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5334_ _1269_ _1286_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__or2_2
X_5265_ _0818_ _1215_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__xnor2_1
X_8053_ _0570_ _3559_ vssd1 vssd1 vccd1 vccd1 _3588_ sky130_fd_sc_hd__xor2_1
XANTENNA__6647__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7004_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1 vssd1 vccd1 vccd1
+ _2765_ sky130_fd_sc_hd__o21ai_1
X_5196_ _0798_ _0794_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8939__A2 _3276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8955_ _4424_ _4427_ _4431_ vssd1 vssd1 vccd1 vccd1 _4432_ sky130_fd_sc_hd__or3b_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7906_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[1\]
+ _3451_ _3452_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__a21o_1
XANTENNA__7369__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout161_X net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8886_ _4360_ _4363_ _4278_ _4358_ vssd1 vssd1 vccd1 vccd1 _4364_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_84_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7837_ net159 _3404_ _3405_ net165 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7768_ net149 net135 _3301_ _3314_ vssd1 vssd1 vccd1 vccd1 _3358_ sky130_fd_sc_hd__or4_1
X_6719_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload2 clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__bufinv_16
X_9507_ net382 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
X_7699_ net153 net135 vssd1 vssd1 vccd1 vccd1 _3289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9438_ clknet_leaf_20_wb_clk_i _0383_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9369_ clknet_leaf_25_wb_clk_i _0317_ net252 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout250 net251 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_2
X_9587__451 vssd1 vssd1 vccd1 vccd1 _9587__451/HI net451 sky130_fd_sc_hd__conb_1
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
Xfanout283 net285 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
Xfanout261 _0514_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_4
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_2
XANTENNA__8663__A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7602__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5086__X _1039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8866__A1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9325__RESET_B net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8866__B2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6629__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5050_ _0999_ _1001_ _1002_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__nor3_1
XFILLER_0_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8573__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5952_ _1885_ _1886_ _1843_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__a21bo_1
XANTENNA__4606__A _0423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8740_ net334 _0405_ _4216_ _4217_ vssd1 vssd1 vccd1 vccd1 _4218_ sky130_fd_sc_hd__a31o_1
X_4903_ _0773_ _0778_ _0779_ _0784_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_62_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5883_ _1797_ _1798_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_62_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8671_ net116 _3608_ _4142_ vssd1 vssd1 vccd1 vccd1 _4150_ sky130_fd_sc_hd__or3_1
X_4834_ _0778_ _0784_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7622_ _3196_ _3211_ vssd1 vssd1 vccd1 vccd1 _3212_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4765_ _0591_ _0714_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__xnor2_4
X_7553_ net257 _3162_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7636__B net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4979__C _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6317__C1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6504_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[4\] _2433_
+ net156 vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__o21ai_1
X_9223_ clknet_leaf_17_wb_clk_i _0067_ net229 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9066__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4696_ net282 _0646_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__or2_1
X_7484_ _3073_ _3122_ _3123_ vssd1 vssd1 vccd1 vccd1 _3124_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8748__A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6435_ _2354_ _2363_ _2382_ vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__and3_1
X_6366_ net318 _2294_ net315 vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8609__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9154_ clknet_leaf_37_wb_clk_i _0255_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5317_ _1038_ _1222_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__xor2_1
X_8105_ _2385_ _0642_ vssd1 vssd1 vccd1 vccd1 _3633_ sky130_fd_sc_hd__nand2b_1
X_9085_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[15\]
+ net222 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_6297_ _0446_ _2204_ _2207_ _2249_ vssd1 vssd1 vccd1 vccd1 _2250_ sky130_fd_sc_hd__a211o_1
X_8036_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] _3561_ vssd1
+ vssd1 vccd1 vccd1 _3572_ sky130_fd_sc_hd__nor2_1
Xhold14 _0246_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _0748_ _0968_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__xnor2_1
Xhold47 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[3\]
+ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[0\] vssd1
+ vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[1\] vssd1
+ vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _1130_ _1131_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__nor2_1
XANTENNA__5900__A _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold69 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[6\]
+ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_08_WB.instance_to_wrap.allocation.game.controller.color\[8\] vssd1 vssd1
+ vccd1 vccd1 net556 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8483__A _3280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4516__A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8938_ _2301_ _4414_ net105 vssd1 vssd1 vccd1 vccd1 _4415_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8869_ net317 _3542_ vssd1 vssd1 vccd1 vccd1 _4347_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_14_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4582__A1 _0419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7833__Y _3403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8000__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4550_ net331 _0422_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4481_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[5\] vssd1
+ vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__inv_2
XANTENNA__7511__A1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8568__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6220_ _2156_ _2172_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _0723_ _0916_ _2097_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_41_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5102_ _1054_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _1959_ _2034_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7814__A2 _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5033_ _0984_ _0985_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__nand2_1
XANTENNA__5720__A _0919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6984_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[23\]
+ _2750_ vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout169_A _0685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5935_ _0813_ _0917_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8750__B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8723_ net319 _4197_ net316 vssd1 vssd1 vccd1 vccd1 _4201_ sky130_fd_sc_hd__a21oi_1
X_5866_ _1816_ _1817_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8654_ net284 net282 _3679_ vssd1 vssd1 vccd1 vccd1 _4133_ sky130_fd_sc_hd__and3_1
X_4817_ _0580_ _0597_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7605_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[10\]
+ _3190_ _3191_ _3194_ vssd1 vssd1 vccd1 vccd1 _3195_ sky130_fd_sc_hd__and4_1
X_5797_ _0743_ _1743_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_32_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7750__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8585_ _0696_ _4063_ vssd1 vssd1 vccd1 vccd1 _4064_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_79_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7536_ net563 _2546_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__xor2_1
X_4748_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\] _0656_
+ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_79_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4679_ _0429_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[2\]
+ _0635_ _0636_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7467_ net114 _3108_ vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9206_ clknet_leaf_10_wb_clk_i _0261_ net229 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr1\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6418_ _2327_ _2337_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7398_ _3041_ _3042_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__or2_2
X_9137_ clknet_leaf_39_wb_clk_i _0238_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_6349_ _2292_ _2300_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__or2_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
X_9068_ clknet_leaf_8_wb_clk_i _0203_ net223 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8463__C1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8019_ _3523_ _3555_ _3551_ net193 vssd1 vssd1 vccd1 vccd1 _3556_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_99_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8005__X _3542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8388__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8835__B _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9273__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5720_ _0919_ _1672_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5991__B1 _0744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ _0773_ _0910_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5582_ _1534_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__inv_2
X_8370_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] _3851_ vssd1
+ vssd1 vccd1 vccd1 _3854_ sky130_fd_sc_hd__xnor2_1
X_4602_ _0487_ _0496_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__xnor2_1
X_4533_ net324 net289 _0501_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__a21o_1
XANTENNA__7914__B team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8288__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7321_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[9\]
+ _2988_ vssd1 vssd1 vccd1 vccd1 _2989_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_96_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7252_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[8\]
+ _2936_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__a31o_1
X_6203_ _1036_ _1065_ _1069_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__o21ai_1
X_9492__367 vssd1 vssd1 vccd1 vccd1 _9492__367/HI net367 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_74_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7930__A team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7183_ net164 _2892_ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__nor2_1
X_6134_ _0754_ _0917_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _2015_ _2017_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_5_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _0798_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout286_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6967_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[17\]
+ _2738_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5918_ _1818_ _1825_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_37_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8706_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\] net113 vssd1
+ vssd1 vccd1 vccd1 _4185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6898_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[3\]
+ _2697_ net267 vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9081__RESET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5849_ net147 _0930_ _1800_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4513__B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8637_ net287 net127 vssd1 vssd1 vccd1 vccd1 _4116_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7723__A1 _3241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5694__A_N _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8568_ net177 _4045_ vssd1 vssd1 vccd1 vccd1 _4047_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7519_ _3040_ _3054_ net305 vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8499_ _3977_ _3978_ _3285_ vssd1 vssd1 vccd1 vccd1 _3979_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input14_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8671__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6214__A1 _1011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7478__B1 _3022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8690__A2 _3608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5270__A _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7870_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[9\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[10\] _3421_
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[11\] vssd1
+ vssd1 vccd1 vccd1 _3429_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6205__A1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6821_ _2646_ _2647_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__nor2_1
XANTENNA__7468__Y _3110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9540_ net408 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_77_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6752_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[10\]
+ _2597_ vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5703_ _1048_ _1644_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__xor2_2
XFILLER_0_72_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6683_ net267 _2549_ _2555_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__and3_1
X_9471_ net346 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_57_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5634_ _1579_ _1581_ _1585_ _1586_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_72_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7925__A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8422_ _3333_ _3355_ _3902_ vssd1 vssd1 vccd1 vccd1 _3903_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8353_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[7\] _3841_
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[6\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[5\]
+ vssd1 vssd1 vccd1 vccd1 _3842_ sky130_fd_sc_hd__and4b_1
X_5565_ _0786_ _1506_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold100 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[6\]
+ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__dlygate4sd3_1
X_7304_ _2972_ _2977_ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__nor2_1
X_5496_ _1447_ _1448_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__nand2_1
Xhold133 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ net328 team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__nor2_1
X_8284_ _3776_ _3777_ net194 vssd1 vssd1 vccd1 vccd1 _3778_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8130__A1 _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold122 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[5\]
+ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout201_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold177 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[3\]
+ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7931__Y _3472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[20\] vssd1 vssd1
+ vccd1 vccd1 net653 sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ net332 vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__inv_2
Xhold166 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[3\] vssd1 vssd1
+ vccd1 vccd1 net664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8756__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7235_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[2\]
+ _2926_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold188 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__dlygate4sd3_1
X_7166_ _0524_ _2881_ _2882_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input6_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6117_ _2068_ _2069_ vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7097_ _2834_ _2835_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[17\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__o211a_1
XANTENNA__8433__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6048_ _0715_ _0928_ _1959_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8197__A1 _3022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7999_ _3519_ _3533_ _3536_ vssd1 vssd1 vccd1 vccd1 _3537_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4758__B2 team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5707__B1 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7880__B1 _3403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5090__A _1038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7745__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9558__426 vssd1 vssd1 vccd1 vccd1 _9558__426/HI net426 sky130_fd_sc_hd__conb_1
XFILLER_0_55_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8896__C1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5265__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5350_ _0999_ _1011_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__and2b_1
XFILLER_0_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8112__A1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5281_ _1169_ _1174_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__and2_1
XANTENNA__8112__B2 team_08_WB.instance_to_wrap.allocation.game.controller.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5477__A2 _1421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7020_ _0460_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[1\] vssd1 vssd1
+ vccd1 vccd1 net62 sky130_fd_sc_hd__a21o_1
XFILLER_0_11_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4609__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8971_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[6\] vssd1 vssd1
+ vccd1 vccd1 _0401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4988__A1 _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7922_ _3457_ _3462_ _3463_ net237 net647 vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_69_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7853_ _3416_ vssd1 vssd1 vccd1 vccd1 _3417_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4996_ _0943_ _0947_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6804_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ _2634_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__or3b_1
XFILLER_0_59_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout151_A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7784_ _2368_ _2383_ _2397_ vssd1 vssd1 vccd1 vccd1 _3371_ sky130_fd_sc_hd__o21ai_1
X_6735_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[5\]
+ _2588_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__and2_1
X_9523_ net398 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
X_9454_ clknet_leaf_46_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[8\]
+ net235 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_61_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9498__373 vssd1 vssd1 vccd1 vccd1 _9498__373/HI net373 sky130_fd_sc_hd__conb_1
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6666_ _2542_ _2543_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[7\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5617_ _1555_ _1567_ _1568_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9385_ clknet_leaf_29_wb_clk_i _0332_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_6597_ _2498_ _2499_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[12\]
+ sky130_fd_sc_hd__nor2_1
X_8405_ net116 _3869_ vssd1 vssd1 vccd1 vccd1 _3886_ sky130_fd_sc_hd__nor2_1
X_5548_ _1497_ _1499_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__xnor2_1
X_8336_ _3819_ _3820_ _3826_ net239 net598 vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__o32a_1
XFILLER_0_14_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4510__C net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8267_ net330 _2268_ vssd1 vssd1 vccd1 vccd1 _3762_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5479_ _1429_ _1431_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7218_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoMovement _0433_ _0565_
+ _2914_ _2916_ vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__a221o_1
XANTENNA__7390__A _2544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8198_ _3711_ _3712_ vssd1 vssd1 vccd1 vccd1 _3713_ sky130_fd_sc_hd__nand2_1
X_7149_ _2866_ _2867_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__nor2_1
XANTENNA__8406__A2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7917__A1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4600__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8342__A1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout94 _3879_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_2
XFILLER_0_25_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4903__A1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5959__S _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4850_ _0786_ _0802_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4781_ _0731_ _0732_ _0733_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__nand3_2
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6520_ _2445_ _2446_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload20 clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload20/X sky130_fd_sc_hd__clkbuf_4
X_6451_ net292 net291 vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__nor2_1
Xclkload42 clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__inv_12
X_5402_ _1354_ _1353_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__and2b_1
XFILLER_0_70_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9170_ _0145_ _0407_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[11\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkload31 clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload31/X sky130_fd_sc_hd__clkbuf_4
X_6382_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.slow_clk
+ _2331_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__nand2_1
X_5333_ _1284_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__nand2_1
X_8121_ _0428_ _3633_ vssd1 vssd1 vccd1 vccd1 _3648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9532__407 vssd1 vssd1 vccd1 vccd1 _9532__407/HI net407 sky130_fd_sc_hd__conb_1
XFILLER_0_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5264_ _0810_ _0913_ _1214_ _0907_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__a2bb2oi_4
XFILLER_0_76_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8052_ _3572_ _3576_ vssd1 vssd1 vccd1 vccd1 _3587_ sky130_fd_sc_hd__nand2b_1
X_7003_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] _2758_ _2763_ _2764_
+ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__o22a_1
X_5195_ _1145_ _1146_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8954_ net177 _3707_ _4419_ _4420_ _4430_ vssd1 vssd1 vccd1 vccd1 _4431_ sky130_fd_sc_hd__a221o_1
XANTENNA__8472__C _3952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7905_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[1\]
+ _3451_ _0713_ vssd1 vssd1 vccd1 vccd1 _3452_ sky130_fd_sc_hd__o21ai_1
X_8885_ net101 _4243_ _4359_ net95 _4362_ vssd1 vssd1 vccd1 vccd1 _4363_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_84_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7836_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[1\] vssd1
+ vssd1 vccd1 vccd1 _3405_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout154_X net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5457__X _1410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4979_ _0809_ _0928_ _0930_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7767_ _3283_ _3341_ _3356_ _3274_ vssd1 vssd1 vccd1 vccd1 _3357_ sky130_fd_sc_hd__a22o_1
XANTENNA__4802__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6718_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[9\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__or4_1
X_9506_ net381 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7698_ net112 _3241_ vssd1 vssd1 vccd1 vccd1 _3288_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload3 clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__inv_6
XFILLER_0_62_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9437_ clknet_leaf_28_wb_clk_i _0382_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6649_ net262 _2477_ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__and2_4
XFILLER_0_21_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9368_ clknet_leaf_25_wb_clk_i _0316_ net252 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9299_ clknet_leaf_12_wb_clk_i _0119_ net217 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_8319_ _3804_ _3810_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[5\]
+ net239 vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5352__B _0999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout240 net242 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
Xfanout273 net276 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_4
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
Xfanout262 _0514_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_4
Xfanout295 team_08_WB.instance_to_wrap.allocation.game.controller.block_done vssd1
+ vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout284 net285 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_2
XANTENNA__4536__X _0505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4652__A_N team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8563__B2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8563__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6574__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7826__B1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8251__B1 _3472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5951_ _1888_ _1901_ _1902_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__nand3_1
XANTENNA__9458__Q team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_dino vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4902_ _0852_ _0854_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8670_ net126 _3681_ vssd1 vssd1 vccd1 vccd1 _4149_ sky130_fd_sc_hd__or2_1
X_5882_ _1819_ _1821_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4833_ _0769_ _0785_ _0766_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7621_ _3188_ _3194_ vssd1 vssd1 vccd1 vccd1 _3211_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4764_ _0591_ _0714_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__xor2_4
X_7552_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr2\[1\] team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr2\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.clk1 vssd1
+ vssd1 vccd1 vccd1 _3162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7483_ _3073_ _3122_ _0438_ vssd1 vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6503_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[3\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[4\]
+ _2431_ vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__and3_1
X_9222_ clknet_leaf_17_wb_clk_i _0066_ net228 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4695_ net282 _0650_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__or2_1
X_6434_ _2358_ _2377_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__or2_1
XANTENNA__8748__B team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5453__A _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6365_ _2310_ _2313_ _2314_ _2316_ vssd1 vssd1 vccd1 vccd1 _2317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8609__A2 _3284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9153_ clknet_leaf_36_wb_clk_i _0254_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_5316_ _1267_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__nand2_1
X_6296_ _0445_ _2206_ _2208_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[12\]
+ _2248_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__a221o_1
X_8104_ _3630_ _3631_ vssd1 vssd1 vccd1 vccd1 _3632_ sky130_fd_sc_hd__nand2_1
X_9084_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[14\]
+ net223 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_5247_ _1194_ _1196_ _1199_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__o21ai_1
X_8035_ _3529_ _3551_ vssd1 vssd1 vccd1 vccd1 _3571_ sky130_fd_sc_hd__and2_1
XANTENNA__9035__RESET_B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8764__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.tft_dc vssd1
+ vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _1124_ _1128_ _1129_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__and3_1
Xhold48 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[17\]
+ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[4\]
+ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5900__B _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8937_ net187 _2307_ _4413_ vssd1 vssd1 vccd1 vccd1 _4414_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_3_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4516__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8868_ _4283_ _4330_ _4279_ vssd1 vssd1 vccd1 vccd1 _4346_ sky130_fd_sc_hd__o21a_1
XANTENNA__8545__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7819_ _2788_ _2795_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _3394_ sky130_fd_sc_hd__o21ai_1
X_8799_ net97 _4266_ _4267_ net103 _4276_ vssd1 vssd1 vccd1 vccd1 _4277_ sky130_fd_sc_hd__o221a_1
XANTENNA__8004__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8010__Y _3547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7036__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8536__B2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8536__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7753__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4480_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.slow_clk
+ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6150_ _0715_ _0916_ _2083_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5101_ _1051_ _1053_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_55_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6081_ net182 _0926_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__nor2_1
X_5032_ _0981_ _0983_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6983_ _2750_ _2417_ _2749_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_0_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5934_ _1843_ _1885_ _1886_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__nand3_1
X_8722_ _4197_ _4198_ _4199_ vssd1 vssd1 vccd1 vccd1 _4200_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5865_ _1816_ _1817_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8653_ _3261_ net98 _3901_ _4131_ vssd1 vssd1 vccd1 vccd1 _4132_ sky130_fd_sc_hd__and4b_1
XFILLER_0_91_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4816_ _0766_ _0768_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__nor2_4
XFILLER_0_76_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout231_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7604_ _3193_ vssd1 vssd1 vccd1 vccd1 _3194_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5796_ _1696_ _1745_ _1746_ _1748_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout329_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8584_ _0687_ _4062_ vssd1 vssd1 vccd1 vccd1 _4063_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9287__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4747_ net139 vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7535_ _2546_ _3153_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_79_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4678_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[1\] vssd1
+ vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout117_X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7466_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_dino _3064_ _3069_
+ vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__or3_1
XANTENNA__5454__Y _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9205_ clknet_leaf_19_wb_clk_i _0260_ net229 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr1\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_7397_ _0441_ _0442_ vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6417_ _2348_ _2366_ _2367_ _2334_ vssd1 vssd1 vccd1 vccd1 _2368_ sky130_fd_sc_hd__o22a_2
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
X_6348_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[3\] _2291_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9136_ clknet_leaf_40_wb_clk_i _0237_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.frameBufferLowNibble
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6279_ _0717_ _0917_ _0921_ net182 vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__o22a_1
X_9067_ clknet_leaf_8_wb_clk_i _0202_ net224 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_76_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8018_ _3553_ _3554_ vssd1 vssd1 vccd1 vccd1 _3555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5029__B1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8454__B1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8509__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5991__A1 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6371__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5650_ _0772_ net145 vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4601_ net332 _0540_ _0562_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[1\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5581_ _1530_ _1531_ _1533_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4532_ _0484_ _0497_ _0500_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__a21oi_1
X_7320_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[8\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[7\]
+ _2987_ vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_57_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4463_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7251_ net581 _2938_ _2940_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__a21oi_1
X_6202_ net138 _1067_ _1070_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7182_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[10\] _2891_ vssd1
+ vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6133_ _2073_ _2084_ _2085_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__nor3_1
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6064_ _1883_ _2016_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5450__B _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5015_ _0744_ _0797_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6966_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[16\]
+ _2737_ _2739_ net158 vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7420__A1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_dino vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5917_ _1865_ _1868_ _1835_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7377__B _2544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8705_ _4176_ _4179_ _4182_ _4183_ vssd1 vssd1 vccd1 vccd1 _4184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6897_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[3\]
+ _2697_ vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5848_ net147 _0930_ _1800_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__nand3_1
XFILLER_0_29_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8636_ _4111_ _4114_ vssd1 vssd1 vccd1 vccd1 _4115_ sky130_fd_sc_hd__nor2_1
X_5779_ _1679_ _1681_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8489__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8567_ net152 _4044_ _4045_ net177 vssd1 vssd1 vccd1 vccd1 _4046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7518_ net307 _3055_ _3040_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7393__A _3034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8498_ _3317_ _3336_ _3897_ vssd1 vssd1 vccd1 vccd1 _3978_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7449_ net304 net309 vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9119_ clknet_leaf_28_wb_clk_i _0220_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.color\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5641__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8671__B _3608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6214__A2 _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5973__A1 _0723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8399__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5094__Y _1047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3__f_wb_clk_i_X clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__8124__C1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7478__A1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8716__A1_N net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4719__X _0674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9390__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6205__A2 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6820_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[5\]
+ _2644_ net271 vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6751_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[10\]
+ _2597_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7765__X _3355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9470_ net345 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
X_5702_ _0758_ _1646_ _1654_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_73_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6682_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__nand2_1
X_5633_ _1534_ _1584_ _1583_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7925__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8902__B2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8421_ _3279_ _3901_ vssd1 vssd1 vccd1 vccd1 _3902_ sky130_fd_sc_hd__nor2_1
X_5564_ _0847_ _1508_ _1516_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8352_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[4\] _3840_
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[2\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3841_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold101 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__dlygate4sd3_1
X_7303_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr1\[0\] team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2977_ sky130_fd_sc_hd__xor2_2
X_4515_ net326 team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9500__375 vssd1 vssd1 vccd1 vccd1 _9500__375/HI net375 sky130_fd_sc_hd__conb_1
X_5495_ _0836_ _0839_ _0745_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__mux2_1
Xhold134 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7941__A _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8283_ net327 _3764_ vssd1 vssd1 vccd1 vccd1 _3777_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold112 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[10\] vssd1 vssd1
+ vccd1 vccd1 net610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[6\] vssd1 vssd1
+ vccd1 vccd1 net621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.wr vssd1
+ vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ net291 vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__inv_2
X_7234_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[1\]
+ _2924_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__a31o_1
XANTENNA__8756__B _3542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold156 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[16\] vssd1
+ vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[7\] vssd1 vssd1
+ vccd1 vccd1 net687 sky130_fd_sc_hd__dlygate4sd3_1
X_7165_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[2\] _2877_ net664
+ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__a21oi_1
Xhold178 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[3\] vssd1 vssd1
+ vccd1 vccd1 net676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6116_ _2060_ _2062_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7096_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[15\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[14\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__or4_1
X_6047_ _0724_ _0926_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7388__A _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7998_ net324 net300 net196 _3535_ vssd1 vssd1 vccd1 vccd1 _3536_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6949_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[10\]
+ _2727_ vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4524__B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5707__A1 _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7394__Y _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8619_ _0695_ _4096_ _4097_ net169 vssd1 vssd1 vccd1 vccd1 _4098_ sky130_fd_sc_hd__o211a_1
X_9599_ net463 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_84_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5355__B _1254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8012__A team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8947__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6132__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout97_X net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5371__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6186__B _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7632__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8688__A_N net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4715__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7745__B _3241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5265__B _1215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8857__A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5280_ _1193_ _1209_ _1212_ _1213_ _1232_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8970_ net297 vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__8592__A _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4988__A2 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7921_ net298 net300 _3461_ vssd1 vssd1 vccd1 vccd1 _3463_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9645__488 vssd1 vssd1 vccd1 vccd1 _9645__488/HI net488 sky130_fd_sc_hd__conb_1
XANTENNA__7001__A team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7852_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[6\]
+ _3413_ vssd1 vssd1 vccd1 vccd1 _3416_ sky130_fd_sc_hd__and2_1
X_4995_ _0943_ _0947_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__nand2_1
X_6803_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7783_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] _2325_ _3370_ net261
+ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9522_ net397 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
X_6734_ _2588_ _2589_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9453_ clknet_leaf_46_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[7\]
+ net235 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5456__A _1217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6665_ net281 _2541_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__nand2_1
X_8404_ net112 _3865_ vssd1 vssd1 vccd1 vccd1 _3885_ sky130_fd_sc_hd__or2_1
X_5616_ _1555_ _1567_ _1568_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9384_ clknet_leaf_31_wb_clk_i _0331_ net245 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_6596_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[12\] _2497_
+ net262 vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5547_ _1497_ _1499_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__and2b_1
X_8335_ _0702_ _2278_ _3825_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _3826_ sky130_fd_sc_hd__a22o_1
XANTENNA__8767__A _0423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5478_ _1408_ _1427_ _1428_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__and3_1
X_8266_ _3759_ _3760_ vssd1 vssd1 vccd1 vccd1 _3761_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7217_ net332 _0562_ _2915_ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5191__A _1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8197_ _3022_ _3033_ _3002_ vssd1 vssd1 vccd1 vccd1 _3712_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7148_ _2859_ _2864_ _2868_ _2857_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__a31oi_1
X_7079_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[4\]
+ _2789_ _2800_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__a22o_1
XANTENNA__4806__Y _0759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9412__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6338__D1 _0684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout95 _3269_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7550__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9159__CLK _0134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4445__A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4780_ _0612_ _0629_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4451__Y _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xclkload10 clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_8
XFILLER_0_15_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6450_ net292 net656 net290 vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__o21a_1
Xclkload43 clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__inv_12
X_5401_ _1304_ _1306_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload21 clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload32 clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__clkinv_4
X_6381_ team_08_WB.instance_to_wrap.allocation.game.game.score\[3\] team_08_WB.instance_to_wrap.allocation.game.game.score\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.game.score\[4\] vssd1 vssd1 vccd1 vccd1
+ _2332_ sky130_fd_sc_hd__nor3_2
X_5332_ _1275_ _1277_ _1283_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__nand3_1
X_8120_ _3645_ _3646_ vssd1 vssd1 vccd1 vccd1 _3647_ sky130_fd_sc_hd__or2_1
XANTENNA__8097__A1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5263_ _1215_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__inv_2
X_8051_ _3472_ _3585_ net298 vssd1 vssd1 vccd1 vccd1 _3586_ sky130_fd_sc_hd__o21a_1
X_9612__476 vssd1 vssd1 vccd1 vccd1 _9612__476/HI net476 sky130_fd_sc_hd__conb_1
X_7002_ _0467_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] _2757_ vssd1
+ vssd1 vccd1 vccd1 _2764_ sky130_fd_sc_hd__a21oi_1
X_5194_ _1145_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_76_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5607__B1 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8953_ _4423_ _4429_ _4422_ vssd1 vssd1 vccd1 vccd1 _4430_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7369__C _2423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7904_ _0434_ _0403_ _3451_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__a21boi_1
X_9465__340 vssd1 vssd1 vccd1 vccd1 _9465__340/HI net340 sky130_fd_sc_hd__conb_1
X_8884_ net101 _4243_ _4247_ _4361_ _4248_ vssd1 vssd1 vccd1 vccd1 _4362_ sky130_fd_sc_hd__a221o_1
XANTENNA__8557__C1 _3280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_A _0514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7835_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[1\] vssd1
+ vssd1 vccd1 vccd1 _3404_ sky130_fd_sc_hd__or2_1
XANTENNA__8021__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8021__B2 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9505_ net380 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4978_ _0729_ _0730_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9506__381 vssd1 vssd1 vccd1 vccd1 _9506__381/HI net381 sky130_fd_sc_hd__conb_1
XFILLER_0_19_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7766_ net97 _3278_ _3355_ _3354_ vssd1 vssd1 vccd1 vccd1 _3356_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_80_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6717_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ _2576_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__or3b_1
XFILLER_0_62_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7697_ net110 net108 vssd1 vssd1 vccd1 vccd1 _3287_ sky130_fd_sc_hd__nor2_1
Xclkload4 clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_6
XFILLER_0_73_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9436_ clknet_leaf_9_wb_clk_i _0381_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6648_ net533 _2529_ _2531_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[31\]
+ sky130_fd_sc_hd__a21oi_1
X_9367_ clknet_leaf_25_wb_clk_i _0315_ net252 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4897__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8318_ net139 _2281_ _3808_ _3809_ vssd1 vssd1 vccd1 vccd1 _3810_ sky130_fd_sc_hd__o211a_1
X_6579_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[5\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[6\]
+ _2484_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__and3_1
X_9298_ clknet_leaf_12_wb_clk_i _0118_ net219 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8249_ _3744_ net255 net291 net269 vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__a2bb2o_1
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_4
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_4
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_4
Xfanout274 net276 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_2
Xfanout263 _0514_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XANTENNA__6745__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 team_08_WB.instance_to_wrap.allocation.game.controller.state\[9\] vssd1
+ vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_2
XANTENNA__8260__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout285 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[6\] vssd1
+ vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8260__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7576__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5096__A _0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7523__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8251__A1 _0552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5950_ _1901_ _1902_ _1888_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__a21o_1
X_4901_ _0851_ _0853_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__and2_1
X_5881_ _1832_ _1833_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_62_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7620_ _3204_ _3206_ _3207_ _3208_ vssd1 vssd1 vccd1 vccd1 _3210_ sky130_fd_sc_hd__and4_1
X_4832_ _0779_ _0783_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7551_ _3160_ _3161_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__nor2_1
X_4763_ _0590_ _0714_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9324__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6317__A1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4694_ _0640_ _0648_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__or2_1
X_7482_ net310 _3051_ net305 vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6502_ _2433_ _2434_ net156 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[3\]
+ sky130_fd_sc_hd__and3b_1
X_9221_ clknet_leaf_17_wb_clk_i _0065_ net229 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6433_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[2\] _2325_
+ _2359_ _2381_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6364_ net327 _2307_ _2308_ vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout107_A _3252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9152_ clknet_leaf_36_wb_clk_i _0253_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_5315_ _1263_ _1266_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6295_ _2209_ _2211_ _2247_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__or3_1
XANTENNA__7817__A1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8103_ net169 _3616_ vssd1 vssd1 vccd1 vccd1 _3631_ sky130_fd_sc_hd__nand2_1
X_9083_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[13\]
+ net222 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5246_ _1197_ _1198_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__or2_1
X_8034_ _3565_ _3569_ _3540_ vssd1 vssd1 vccd1 vccd1 _3570_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8490__A1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold38 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[21\]
+ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[7\] vssd1
+ vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[0\]
+ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _1124_ _1128_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8256__S net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold49 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[4\]
+ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8109__X _3637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9075__RESET_B net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8936_ net190 _2306_ _2307_ net187 _4412_ vssd1 vssd1 vccd1 vccd1 _4413_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8867_ _4279_ _4330_ _4332_ net96 _4344_ vssd1 vssd1 vccd1 vccd1 _4345_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7818_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\] _2793_
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\] vssd1
+ vssd1 vccd1 vccd1 _3393_ sky130_fd_sc_hd__a31oi_4
X_8798_ net103 _4267_ _4274_ _4275_ vssd1 vssd1 vccd1 vccd1 _4276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7749_ _3254_ net104 _0556_ vssd1 vssd1 vccd1 vccd1 _3339_ sky130_fd_sc_hd__or3b_2
XFILLER_0_19_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9419_ clknet_leaf_42_wb_clk_i _0364_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input37_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6475__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5097__Y _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5100_ _1012_ _1050_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__nand2_1
X_6080_ _0772_ _0916_ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_55_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5031_ _0981_ _0983_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6982_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[22\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[21\]
+ _2747_ vssd1 vssd1 vccd1 vccd1 _2750_ sky130_fd_sc_hd__and3_1
X_8721_ _0520_ _4197_ net313 vssd1 vssd1 vccd1 vccd1 _4199_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5933_ _1795_ _1837_ _1842_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__a21o_1
XANTENNA__7928__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_5864_ _1767_ _1768_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7735__B1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8652_ _4004_ _4054_ _4108_ _4130_ vssd1 vssd1 vccd1 vccd1 _4131_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4815_ _0758_ _0765_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7603_ net184 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\]
+ net176 _3192_ vssd1 vssd1 vccd1 vccd1 _3193_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8583_ net178 _4061_ vssd1 vssd1 vccd1 vccd1 _4062_ sky130_fd_sc_hd__nor2_1
X_5795_ _1696_ _1745_ _1747_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7534_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[2\]
+ _2545_ net601 vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout224_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4746_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\] _0700_ vssd1
+ vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7663__B net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4677_ net293 _0605_ _0634_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__and3_2
XFILLER_0_32_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7465_ _3102_ _3103_ _3106_ vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__a21oi_1
X_9204_ clknet_leaf_11_wb_clk_i _0025_ net219 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_7396_ net309 net308 vssd1 vssd1 vccd1 vccd1 _3041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6416_ _2366_ team_08_WB.instance_to_wrap.allocation.game.game.score\[1\] _2336_
+ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__mux2_1
XANTENNA__6847__X _2665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6347_ net315 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[6\] _2297_
+ _2298_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9135_ clknet_leaf_37_wb_clk_i net115 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ sky130_fd_sc_hd__dfxtp_4
XANTENNA__9256__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6278_ _2106_ _2230_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__nand2_1
X_9066_ clknet_leaf_8_wb_clk_i _0201_ net223 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5229_ _1181_ _1179_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__nand2b_1
X_8017_ _3528_ _3550_ vssd1 vssd1 vccd1 vccd1 _3554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8919_ net169 net136 net127 _0674_ vssd1 vssd1 vccd1 vccd1 _4396_ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8454__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7588__X _3178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5549__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4453__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5268__B _1217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4600_ _0541_ _0560_ net260 vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5580_ _1505_ _1532_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4531_ _0498_ _0499_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4462_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__inv_2
X_7250_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[8\]
+ _2938_ net179 vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__o21ai_1
X_6201_ _1078_ _1079_ _1081_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7181_ _2874_ _2890_ _2891_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__nor3_1
XFILLER_0_1_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6132_ net168 _0922_ _2072_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8445__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6063_ _0715_ net146 _0905_ _0717_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__o2bb2a_1
X_5014_ _0959_ _0966_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7939__A _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6965_ _2738_ vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7420__A2 _3064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5459__A _0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5916_ _1835_ _1868_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8704_ net150 _4178_ _4180_ _4176_ vssd1 vssd1 vccd1 vccd1 _4183_ sky130_fd_sc_hd__o211a_1
X_6896_ net274 _2696_ _2697_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__nor3_1
X_8635_ _4112_ _4113_ vssd1 vssd1 vccd1 vccd1 _4114_ sky130_fd_sc_hd__nand2_1
X_5847_ _0773_ _0929_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5778_ _1728_ _1730_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8566_ _0696_ _4043_ vssd1 vssd1 vccd1 vccd1 _4045_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8133__B1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4729_ _0680_ _0683_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__xnor2_2
X_7517_ _3040_ _3074_ _3149_ net308 vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8497_ _3974_ _3976_ _3973_ vssd1 vssd1 vccd1 vccd1 _3977_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7448_ _3043_ _3046_ vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__or2_1
XANTENNA__8684__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7379_ _3028_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9118_ clknet_leaf_19_wb_clk_i _0219_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.clk1
+ sky130_fd_sc_hd__dfxtp_1
X_9049_ clknet_leaf_35_wb_clk_i _0184_ net246 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6753__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4720__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4448__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7938__B1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6750_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[10\]
+ _2597_ _2599_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5701_ _1653_ _1652_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6681_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ net270 _2553_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__and3b_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5632_ _1534_ _1583_ _1584_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_75_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8902__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8420_ _3329_ _3353_ vssd1 vssd1 vccd1 vccd1 _3901_ sky130_fd_sc_hd__nor2_2
X_5563_ _1515_ _1514_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8351_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[1\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[3\]
+ _0517_ vssd1 vssd1 vccd1 vccd1 _3840_ sky130_fd_sc_hd__or3b_1
XFILLER_0_5_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7302_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr1\[1\] team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__xnor2_1
X_4514_ _0481_ _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5494_ _0827_ _1446_ _0828_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__o21ba_1
Xhold113 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__dlygate4sd3_1
X_8282_ net334 _3775_ vssd1 vssd1 vccd1 vccd1 _3776_ sky130_fd_sc_hd__or2_2
Xhold157 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7941__B _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold168 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[2\]
+ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__dlygate4sd3_1
X_7233_ net641 _2926_ _2928_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__o21a_1
Xhold146 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[19\] vssd1
+ vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ net292 vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__inv_2
X_7164_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[3\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[2\]
+ _2877_ vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold179 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[7\] vssd1
+ vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5461__B _1410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6115_ _2067_ _2066_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7095_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[9\]
+ _2833_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__o211a_1
X_6046_ net182 _0929_ _1960_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__or3_1
XANTENNA__4508__D _0478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_X net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7997_ _3505_ _3526_ _3534_ net297 vssd1 vssd1 vccd1 vccd1 _3535_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6948_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[10\]
+ _2727_ vssd1 vssd1 vccd1 vccd1 _2728_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7675__Y _3265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6879_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[12\]
+ _2684_ vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__and2_1
X_9598_ net462 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__5707__A2 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8618_ net162 net155 vssd1 vssd1 vccd1 vccd1 _4097_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8549_ _0432_ net106 _4006_ vssd1 vssd1 vccd1 vccd1 _4028_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8012__B _3543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9200__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6132__A2 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5652__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9482__357 vssd1 vssd1 vccd1 vccd1 _9482__357/HI net357 sky130_fd_sc_hd__conb_1
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8345__B1 _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8896__A1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7518__S _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9523__398 vssd1 vssd1 vccd1 vccd1 _9523__398/HI net398 sky130_fd_sc_hd__conb_1
XANTENNA__7745__C _3305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8857__B _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8648__A1 _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4449__Y _0423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4906__A _0634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7920_ net277 _3017_ vssd1 vssd1 vccd1 vccd1 _3462_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7851_ net159 _3414_ _3415_ net165 net691 vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6802_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4994_ _0945_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7782_ _2368_ _3369_ vssd1 vssd1 vccd1 vccd1 _3370_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6733_ net638 _2586_ net267 vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9521_ net396 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__8336__B1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5737__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6664_ net281 _2541_ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__or2_1
X_9452_ clknet_leaf_48_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[6\]
+ net225 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5615_ _1517_ _1518_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__xor2_1
X_8403_ net112 _3865_ vssd1 vssd1 vccd1 vccd1 _3884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9383_ clknet_leaf_32_wb_clk_i _0330_ net245 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6595_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[12\] _2497_
+ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__and2_1
X_5546_ _0749_ _1498_ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__nor2_1
X_8334_ net194 _3822_ _3823_ _3824_ net170 vssd1 vssd1 vccd1 vccd1 _3825_ sky130_fd_sc_hd__a311o_1
X_5477_ _1402_ _1421_ _1423_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__a21bo_1
X_8265_ _0491_ _0550_ _3492_ _3758_ vssd1 vssd1 vccd1 vccd1 _3760_ sky130_fd_sc_hd__nand4_1
XFILLER_0_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7216_ _0540_ _0562_ net332 vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8196_ net122 _3027_ vssd1 vssd1 vccd1 vccd1 _3711_ sky130_fd_sc_hd__nand2_1
XANTENNA__8783__A _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7147_ _2859_ _2873_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7078_ _2819_ _2820_ _2822_ _2818_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__o31a_1
XANTENNA__4816__A _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6029_ net182 _0860_ _1980_ _1981_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_5_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__8007__B _3542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4822__Y _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4551__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout96 _3269_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6478__A team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8396__C _3355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8802__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_X net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4726__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9564__432 vssd1 vssd1 vccd1 vccd1 _9564__432/HI net432 sky130_fd_sc_hd__conb_1
XFILLER_0_59_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5557__A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9193__RESET_B net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7772__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5400_ _1349_ _1352_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__nand2b_1
Xclkload44 clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__inv_12
Xclkload22 clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__clkinv_4
Xclkload11 clknet_leaf_47_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_8
X_6380_ team_08_WB.instance_to_wrap.allocation.game.game.score\[6\] team_08_WB.instance_to_wrap.allocation.game.game.score\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__nand2_2
Xclkload33 clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_11_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5331_ _1275_ _1277_ _1283_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9571__436 vssd1 vssd1 vccd1 vccd1 _9571__436/HI net436 sky130_fd_sc_hd__conb_1
XANTENNA__5292__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8050_ net197 _3581_ _3583_ _3584_ vssd1 vssd1 vccd1 vccd1 _3585_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7001_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] _2755_ vssd1 vssd1
+ vccd1 vccd1 _2763_ sky130_fd_sc_hd__nor2_1
X_5262_ _0907_ _1214_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__xor2_4
X_5193_ _0747_ _1091_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4907__Y _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5607__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5607__B2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8108__A _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8952_ _2537_ net119 _4428_ vssd1 vssd1 vccd1 vccd1 _4429_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7903_ _0713_ _2841_ _0434_ vssd1 vssd1 vccd1 vccd1 _3451_ sky130_fd_sc_hd__a21o_1
X_8883_ _4237_ _4287_ vssd1 vssd1 vccd1 vccd1 _4361_ sky130_fd_sc_hd__nand2b_1
XANTENNA__8557__B1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6851__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7834_ net159 net165 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__mux2_1
XANTENNA__8021__A2 _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7765_ _0555_ _3351_ vssd1 vssd1 vccd1 vccd1 _3355_ sky130_fd_sc_hd__or2_4
XFILLER_0_74_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6716_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__or4_1
X_4977_ _0729_ _0730_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__xor2_4
X_9504_ net379 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_46_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload5 clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_8
X_7696_ net106 _3261_ vssd1 vssd1 vccd1 vccd1 _3286_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9435_ clknet_leaf_29_wb_clk_i _0380_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6647_ net533 _2529_ net259 vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__o21ai_1
X_9366_ clknet_leaf_25_wb_clk_i _0314_ net250 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6578_ _2486_ _2487_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5529_ _1424_ _1426_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__or2_1
X_8317_ _2296_ net161 _2425_ _3543_ _3636_ vssd1 vssd1 vccd1 vccd1 _3809_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6099__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9297_ clknet_leaf_12_wb_clk_i _0116_ net219 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_8248_ net292 _3746_ _3745_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_2
X_8179_ _2389_ _2390_ _3696_ vssd1 vssd1 vccd1 vccd1 _3697_ sky130_fd_sc_hd__a21oi_1
Xfanout264 net266 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_2
Xfanout253 net254 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_4
Xfanout242 net254 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5930__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8245__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 net276 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_2
X_9548__416 vssd1 vssd1 vccd1 vccd1 _9548__416/HI net416 sky130_fd_sc_hd__conb_1
XANTENNA__4817__Y _0770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout297 team_08_WB.instance_to_wrap.allocation.game.controller.state\[8\] vssd1
+ vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_2
Xfanout286 net288 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_2
XANTENNA__4546__A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6480__B net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7771__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9594__458 vssd1 vssd1 vccd1 vccd1 _9594__458/HI net458 sky130_fd_sc_hd__conb_1
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5840__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7531__S team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8787__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9488__363 vssd1 vssd1 vccd1 vccd1 _9488__363/HI net363 sky130_fd_sc_hd__conb_1
XANTENNA__4456__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8251__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9374__RESET_B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5880_ _1782_ _1783_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4900_ _0846_ _0850_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4831_ _0738_ net141 vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_62_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9303__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7550_ net672 team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr2\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr2\[1\] net257 vssd1
+ vssd1 vccd1 vccd1 _3161_ sky130_fd_sc_hd__a31o_1
X_4762_ _0590_ _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4693_ _0648_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__inv_2
X_7481_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_floor team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_cactus
+ _3066_ _3068_ vssd1 vssd1 vccd1 vccd1 _3121_ sky130_fd_sc_hd__nor4_2
X_6501_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[3\] _2431_
+ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9220_ clknet_leaf_17_wb_clk_i _0064_ net227 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_6432_ net259 _2380_ vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9151_ clknet_leaf_37_wb_clk_i net508 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataDc
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6363_ net335 team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[0\] _2304_
+ _2314_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__a211o_1
X_8102_ net169 _3616_ vssd1 vssd1 vccd1 vccd1 _3630_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5314_ _1263_ _1266_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6294_ _0444_ _2210_ _2212_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[10\]
+ _2246_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__a221o_1
X_9082_ clknet_leaf_49_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[12\]
+ net222 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5245_ _1194_ _1196_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__xnor2_1
X_8033_ _0505_ _3567_ _3568_ vssd1 vssd1 vccd1 vccd1 _3569_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8490__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold28 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[7\]
+ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 _0251_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ _0992_ _0994_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__xnor2_1
Xhold39 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[3\]
+ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8432__D_N _3895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8935_ net190 _2306_ _3284_ _4411_ vssd1 vssd1 vccd1 vccd1 _4412_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5468__Y _1421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8866_ net96 _4332_ _4333_ net102 _4343_ vssd1 vssd1 vccd1 vccd1 _4344_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7817_ team_08_WB.instance_to_wrap.allocation.game.controller.block_done team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ net293 vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__mux2_1
X_8797_ _4268_ _4273_ net104 vssd1 vssd1 vccd1 vccd1 _4275_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7748_ _3270_ _3275_ vssd1 vssd1 vccd1 vccd1 _3338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7679_ _3247_ _3267_ vssd1 vssd1 vccd1 vccd1 _3269_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9418_ clknet_leaf_42_wb_clk_i _0363_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9349_ clknet_leaf_33_wb_clk_i _0297_ net247 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.wr
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7808__A2 _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8019__Y _3556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7526__S team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5030_ _0882_ _0888_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6385__B net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6981_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[21\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[20\]
+ _2744_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[22\]
+ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5932_ _1841_ _1883_ _1884_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__and3_1
X_8720_ net319 net313 net316 vssd1 vssd1 vccd1 vccd1 _4198_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5863_ _1789_ _1797_ _1798_ _1814_ _1815_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8932__B1 _3265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7735__A1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8651_ net106 _4115_ _4129_ vssd1 vssd1 vccd1 vccd1 _4130_ sky130_fd_sc_hd__and3_1
X_4814_ _0766_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__inv_2
X_5794_ _0755_ net146 _0910_ _0724_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_56_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7602_ net184 net176 _3181_ vssd1 vssd1 vccd1 vccd1 _3192_ sky130_fd_sc_hd__a21oi_1
X_8582_ _3595_ _3610_ vssd1 vssd1 vccd1 vccd1 _4061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4745_ _0692_ _0697_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7533_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[2\]
+ _2545_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9577__442 vssd1 vssd1 vccd1 vccd1 _9577__442/HI net442 sky130_fd_sc_hd__conb_1
XFILLER_0_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4676_ _0631_ _0632_ _0606_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__a21o_4
XFILLER_0_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7464_ net301 _3104_ _3105_ _3023_ vssd1 vssd1 vccd1 vccd1 _3106_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9203_ clknet_leaf_11_wb_clk_i _0024_ net220 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7395_ _3023_ _3032_ _3038_ _3040_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6415_ _2326_ _2365_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6346_ net318 _2293_ _2296_ net321 vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__o2bb2a_1
X_9134_ clknet_leaf_38_wb_clk_i _0235_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4795__S _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9065_ clknet_leaf_48_wb_clk_i _0200_ net225 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_6277_ _2103_ _2105_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__or2_1
X_8016_ _3528_ _3550_ vssd1 vssd1 vccd1 vccd1 _3553_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8463__A2 _3895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5228_ _1178_ _1180_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__nand2_1
XANTENNA__4808__B _0759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5159_ _0874_ _1111_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__or2_1
XANTENNA__8791__A _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7974__B2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7974__A1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8918_ _0657_ net109 _4394_ vssd1 vssd1 vccd1 vccd1 _4395_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8849_ _4198_ _4323_ _4326_ vssd1 vssd1 vccd1 vccd1 _4327_ sky130_fd_sc_hd__or3b_1
XANTENNA__7694__X _3284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4549__D_N net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4530_ _0423_ net289 vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4461_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.drawDoneDino vssd1 vssd1
+ vccd1 vccd1 _0433_ sky130_fd_sc_hd__inv_2
X_6200_ _1086_ _2152_ _1084_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__a21oi_1
X_7180_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[8\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[9\]
+ _2887_ vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _2034_ _2083_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__nand2_1
XANTENNA__4909__A _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6062_ _2013_ _2014_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5013_ _0964_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__nor2_1
XANTENNA__7939__B net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout167_A _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6964_ _2408_ _2734_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5459__B _1215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5915_ _1866_ _1867_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__and2_1
X_6895_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_37_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8703_ net288 net125 _4117_ _4181_ net134 vssd1 vssd1 vccd1 vccd1 _4182_ sky130_fd_sc_hd__a32o_1
X_5846_ _1797_ _1798_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__nand2_1
X_8634_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\] net109 vssd1
+ vssd1 vccd1 vccd1 _4113_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout334_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5777_ _1620_ _1729_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8565_ net163 _4039_ vssd1 vssd1 vccd1 vccd1 _4044_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4728_ _0681_ _0682_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__nor2_1
X_7516_ _3149_ _3150_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8496_ net110 net108 _3864_ _3888_ _3975_ vssd1 vssd1 vccd1 vccd1 _3976_ sky130_fd_sc_hd__a41o_1
XFILLER_0_71_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4659_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[3\] vssd1
+ vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__nand2b_1
X_7447_ _3046_ _3056_ _3089_ _3048_ vssd1 vssd1 vccd1 vccd1 _3090_ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7690__A _3265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5481__Y _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7378_ _3002_ _3027_ vssd1 vssd1 vccd1 vccd1 _3028_ sky130_fd_sc_hd__or2_2
XFILLER_0_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9117_ clknet_leaf_33_wb_clk_i _0404_ net247 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6329_ _2278_ _2280_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9048_ clknet_leaf_36_wb_clk_i _0183_ net248 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6998__A2 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5186__A1 _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8124__A1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8696__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8427__A2 _3355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9528__403 vssd1 vssd1 vccd1 vccd1 _9528__403/HI net403 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_29_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_34_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5700_ _0757_ _1646_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6680_ _2553_ vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5631_ _1530_ _1531_ _1533_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5562_ _0846_ _1508_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__xor2_1
X_8350_ net596 net241 _3839_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4513_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] net320 vssd1
+ vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__and2b_1
X_7301_ net284 net263 _0644_ _2973_ vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__nand4_4
X_8281_ net326 _3763_ vssd1 vssd1 vccd1 vccd1 _3775_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5493_ _0813_ _1445_ _0816_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__mux2_1
Xhold125 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[4\]
+ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__dlygate4sd3_1
X_7232_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[2\]
+ _2926_ net179 vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7874__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold136 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[0\] vssd1 vssd1
+ vccd1 vccd1 net645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold158 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[4\] vssd1
+ vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold169 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ _0523_ _2879_ _2880_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6114_ _2046_ _2047_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7094_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6045_ net148 _0916_ vssd1 vssd1 vccd1 vccd1 _1998_ sky130_fd_sc_hd__and2_1
XANTENNA__6854__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8051__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7996_ net325 _3505_ vssd1 vssd1 vccd1 vccd1 _3534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6947_ _2727_ net157 _2726_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__and3b_1
XFILLER_0_53_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6878_ net273 _2683_ _2684_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__nor3_1
XFILLER_0_64_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7157__A2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9597_ net461 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_91_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5829_ _0919_ _1671_ _0935_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__o21a_1
XANTENNA__4821__B _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8617_ net162 net155 vssd1 vssd1 vccd1 vccd1 _4096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4915__A1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8548_ _0697_ _4016_ _0694_ vssd1 vssd1 vccd1 vccd1 _4027_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8479_ _3300_ _3864_ vssd1 vssd1 vccd1 vccd1 _3959_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4549__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6483__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8593__B2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8593__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4603__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9638__486 vssd1 vssd1 vccd1 vccd1 _9638__486/HI net486 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_93_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9328__RESET_B net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6658__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4459__A team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7084__A1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4842__A0 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7850_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[4\]
+ _3408_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _3415_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6801_ net599 net275 vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__nor2_1
X_4993_ _0868_ _0871_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_86_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7781_ _2361_ _2383_ _2399_ _2380_ vssd1 vssd1 vccd1 vccd1 _3369_ sky130_fd_sc_hd__o31a_1
XFILLER_0_19_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9520_ net395 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6732_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[4\]
+ _2585_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9451_ clknet_leaf_46_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[5\]
+ net235 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_6663_ net283 _2539_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[6\]
+ sky130_fd_sc_hd__xor2_1
X_5614_ _1565_ _1566_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__nand2_1
X_8402_ net173 _3868_ vssd1 vssd1 vccd1 vccd1 _3883_ sky130_fd_sc_hd__nand2_1
X_9382_ clknet_leaf_33_wb_clk_i _0329_ net245 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6594_ _2497_ _2478_ _2496_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[11\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5545_ _0792_ _0859_ _0802_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__a21oi_1
X_8333_ net194 _3561_ vssd1 vssd1 vccd1 vccd1 _3824_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5476_ _1408_ _1427_ _1428_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8264_ _0491_ _0550_ _3492_ _3758_ vssd1 vssd1 vccd1 vccd1 _3759_ sky130_fd_sc_hd__a22o_1
XANTENNA__7311__A2 _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5472__B _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7215_ _0561_ _0563_ _0422_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__o21ai_1
X_8195_ net545 _2983_ vssd1 vssd1 vccd1 vccd1 _3710_ sky130_fd_sc_hd__nand2_1
X_7146_ _2864_ _2868_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7077_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[3\]
+ _2789_ _2799_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[3\]
+ _2821_ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__a221o_1
X_6028_ _1940_ _1979_ _1978_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4833__B1 _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7686__Y _3276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7979_ _0500_ _3516_ vssd1 vssd1 vccd1 vccd1 _3517_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6338__B1 _2288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4551__B net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout97 _3268_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8974__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8587__B1_N net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6577__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7529__S team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5838__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8318__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4742__A _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5557__B _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload23 clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload23/X sky130_fd_sc_hd__clkbuf_4
Xclkload12 clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_12
Xclkload34 clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_11_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5573__A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5330_ _1281_ _1282_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__nand2_1
Xclkload45 clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__inv_4
XFILLER_0_11_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5261_ _0911_ _0913_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__and2_2
XFILLER_0_50_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7000_ _0467_ _0468_ _2755_ _2762_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__a31oi_4
X_5192_ net143 _1144_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_44_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5607__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8951_ _0647_ _4189_ _4128_ vssd1 vssd1 vccd1 vccd1 _4428_ sky130_fd_sc_hd__o21ai_1
X_7902_ net665 _3450_ _2922_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_92_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8557__A1 _3355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8882_ net95 _4359_ vssd1 vssd1 vccd1 vccd1 _4360_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_84_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7833_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[2\]
+ _3393_ _3397_ vssd1 vssd1 vccd1 vccd1 _3403_ sky130_fd_sc_hd__a21oi_2
XANTENNA__5748__A _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7764_ net99 _3353_ _3330_ vssd1 vssd1 vccd1 vccd1 _3354_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6715_ net535 _2573_ _2575_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__a21oi_1
X_4976_ _0731_ _0732_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout247_A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9503_ net378 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
X_7695_ net97 _3278_ _3284_ _3283_ vssd1 vssd1 vccd1 vccd1 _3285_ sky130_fd_sc_hd__o31ai_2
X_9434_ clknet_leaf_29_wb_clk_i _0379_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload6 clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_6_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6646_ _2529_ _2530_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[30\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9365_ clknet_leaf_26_wb_clk_i _0313_ net250 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_6577_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[5\] _2484_ net262
+ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__o21ai_1
X_5528_ _1456_ _1479_ _1480_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8316_ net170 _3807_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _3808_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9296_ clknet_leaf_12_wb_clk_i _0115_ net219 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5459_ _0867_ _1215_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__xnor2_1
X_8247_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.state\[0\] _3743_
+ net291 vssd1 vssd1 vccd1 vccd1 _3746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout232 net254 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
Xfanout221 net232 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
X_8178_ net282 _2390_ _2387_ vssd1 vssd1 vccd1 vccd1 _3696_ sky130_fd_sc_hd__o21ai_1
Xfanout210 net212 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_1
Xfanout254 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.reset
+ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_4
Xfanout243 net253 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_4
X_7129_ net184 _2851_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__a21oi_1
Xfanout276 _2547_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_2
Xfanout298 team_08_WB.instance_to_wrap.allocation.game.controller.state\[8\] vssd1
+ vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_2
Xfanout287 net288 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_2
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8548__A1 _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7771__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8969__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5393__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5840__B _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8787__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4830_ _0738_ net141 vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__and2_2
XFILLER_0_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4761_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[0\] vssd1
+ vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__and2b_4
XFILLER_0_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4692_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[4\] _0647_ vssd1
+ vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__or2_2
X_7480_ net521 net114 _3110_ _3120_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__o22a_1
X_6500_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[3\] _2431_
+ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6431_ net255 _2380_ _2325_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6362_ _2310_ _2312_ _2313_ vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__or3b_1
XFILLER_0_11_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9150_ clknet_leaf_41_wb_clk_i net515 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5313_ _1265_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__inv_2
X_8101_ _3614_ _3627_ _3628_ _0431_ vssd1 vssd1 vccd1 vccd1 _3629_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6293_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[10\]
+ _2212_ _2214_ _2245_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_41_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9081_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[11\]
+ net224 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_5244_ _0819_ _0862_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__nor2_1
X_8032_ _0505_ _3567_ net199 vssd1 vssd1 vccd1 vccd1 _3568_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5175_ _1127_ _1125_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__nand2b_1
Xhold18 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[2\] vssd1
+ vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 _0244_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8490__A3 _3864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8778__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6789__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6862__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9011__Q team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8934_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[0\]
+ _4410_ net192 vssd1 vssd1 vccd1 vccd1 _4411_ sky130_fd_sc_hd__a22o_1
X_8865_ net102 _4333_ _4342_ vssd1 vssd1 vccd1 vccd1 _4343_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7816_ net293 net574 net575 _3392_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5197__B _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8796_ _4268_ _4273_ vssd1 vssd1 vccd1 vccd1 _4274_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout152_X net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4959_ _0739_ _0911_ _0907_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8789__A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7747_ _3317_ _3336_ _3304_ vssd1 vssd1 vccd1 vccd1 _3337_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9084__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7678_ _3247_ _3267_ vssd1 vssd1 vccd1 vccd1 _3268_ sky130_fd_sc_hd__xor2_2
XFILLER_0_85_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9013__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6629_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[24\] _2518_
+ net260 vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__o21ai_1
X_9417_ clknet_leaf_42_wb_clk_i _0362_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9348_ clknet_leaf_46_wb_clk_i _0296_ net235 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[5\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9279_ clknet_leaf_5_wb_clk_i net555 net204 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7744__A2 _0425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9602__466 vssd1 vssd1 vccd1 vccd1 _9602__466/HI net466 sky130_fd_sc_hd__conb_1
XFILLER_0_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6704__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9393__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7417__D1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7968__C1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6980_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[21\]
+ _2747_ _2748_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_0_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7778__A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5931_ _1838_ _1840_ _1839_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5862_ _1789_ _1799_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7735__A2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8650_ _2536_ _4116_ _4127_ _4128_ vssd1 vssd1 vccd1 vccd1 _4129_ sky130_fd_sc_hd__a211oi_1
X_4813_ _0758_ _0765_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__and2_2
X_5793_ _0761_ _0905_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7601_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[11\]
+ net153 vssd1 vssd1 vccd1 vccd1 _3191_ sky130_fd_sc_hd__xnor2_2
X_8581_ _4055_ _4056_ _4059_ _4036_ vssd1 vssd1 vccd1 vccd1 _4060_ sky130_fd_sc_hd__o31a_1
XFILLER_0_84_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4744_ _0698_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7532_ net507 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[8\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet vssd1 vssd1
+ vccd1 vccd1 _0252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8402__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8145__C1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9202_ clknet_leaf_11_wb_clk_i _0023_ net218 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_4675_ _0606_ _0632_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7463_ _0437_ net309 _0442_ vssd1 vssd1 vccd1 vccd1 _3105_ sky130_fd_sc_hd__a21o_1
X_7394_ _3026_ _3037_ vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout112_A _3234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6414_ team_08_WB.instance_to_wrap.allocation.game.game.score\[0\] team_08_WB.instance_to_wrap.allocation.game.game.score\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__nor2_1
X_6345_ net315 _2294_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9133_ clknet_leaf_41_wb_clk_i _0234_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_6276_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[3\]
+ _2228_ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__nor2_1
X_9064_ clknet_leaf_47_wb_clk_i _0199_ net225 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_5227_ _1167_ _1175_ _1177_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__or3_1
X_8015_ _3528_ _3550_ vssd1 vssd1 vccd1 vccd1 _3552_ sky130_fd_sc_hd__nor2_1
X_5158_ _0845_ _0873_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__nor2_1
X_5089_ _1039_ _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__xor2_1
XANTENNA__8136__X _3662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7688__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7974__A2 _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8917_ _0432_ net107 _4007_ vssd1 vssd1 vccd1 vccd1 _4394_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4824__B _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5001__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8848_ _4227_ _4228_ _4319_ _4325_ vssd1 vssd1 vccd1 vccd1 _4326_ sky130_fd_sc_hd__or4_1
X_8779_ _3313_ _3860_ vssd1 vssd1 vccd1 vccd1 _4257_ sky130_fd_sc_hd__nor2_1
XANTENNA__4840__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5936__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5671__A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8982__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6007__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4460_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\] vssd1 vssd1
+ vccd1 vccd1 _0432_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9537__493 vssd1 vssd1 vccd1 vccd1 net493 _9537__493/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_74_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6130_ _0717_ _0921_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4909__B _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6061_ _2011_ _2012_ _1998_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__a21oi_1
XANTENNA__6456__A2 _2325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5012_ _0767_ _0963_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6963_ _2737_ net158 _2736_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__and3b_1
XFILLER_0_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5914_ _0755_ _0859_ _1014_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6894_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__a21oi_1
X_8702_ _0640_ _2385_ vssd1 vssd1 vccd1 vccd1 _4181_ sky130_fd_sc_hd__nand2_1
X_5845_ _1749_ _1750_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__xnor2_2
XANTENNA__8905__A1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8633_ _0426_ _3241_ vssd1 vssd1 vccd1 vccd1 _4112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5756__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5776_ _0742_ _1619_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout327_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8564_ net163 _4039_ vssd1 vssd1 vccd1 vccd1 _4043_ sky130_fd_sc_hd__and2_1
X_4727_ net282 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__nor2_1
X_7515_ net309 _3040_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__or2_1
X_8495_ net116 _3300_ _3359_ _3870_ vssd1 vssd1 vccd1 vccd1 _3975_ sky130_fd_sc_hd__a31o_1
X_4658_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[3\] vssd1
+ vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7446_ _0440_ _3072_ vssd1 vssd1 vccd1 vccd1 _3089_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7690__B net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9116_ clknet_leaf_33_wb_clk_i _0403_ net247 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_7377_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[2\] _2544_
+ _3026_ vssd1 vssd1 vccd1 vccd1 _3027_ sky130_fd_sc_hd__or3b_1
X_4589_ net191 _0405_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4819__B _0770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6328_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[5\] _2273_ vssd1
+ vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__and2_1
XANTENNA__8436__A3 _3916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6259_ _2032_ _2119_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__xnor2_1
X_9047_ clknet_leaf_36_wb_clk_i _0182_ net248 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7689__Y _3279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4835__A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4554__B _0522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5186__A2 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8977__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4584__A_N net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6944__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9608__472 vssd1 vssd1 vccd1 vccd1 _9608__472/HI net472 sky130_fd_sc_hd__conb_1
XFILLER_0_98_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8348__C1 _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5630_ _1553_ _1582_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5561_ _1509_ _1510_ _1513_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5492_ _0813_ _0860_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4512_ net319 team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__and2b_1
X_8280_ _3772_ _3773_ vssd1 vssd1 vccd1 vccd1 _3774_ sky130_fd_sc_hd__nor2_1
X_7300_ net283 net262 _0644_ _2973_ vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__and4_4
XANTENNA__7791__A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[5\]
+ vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__dlygate4sd3_1
X_7231_ _2926_ _2927_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__nor2_1
Xhold148 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7162_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[2\] _2877_ vssd1
+ vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7093_ team_08_WB.EN_VAL_REG net264 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__or2_1
XFILLER_0_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6113_ _0772_ _0916_ _2044_ _2043_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6044_ _1984_ _1985_ _1980_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__o21bai_1
XANTENNA__6854__B _2665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_A _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8051__A1 _3472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7995_ net300 _3531_ _3532_ net193 vssd1 vssd1 vccd1 vccd1 _3533_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6870__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6946_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[9\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[8\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[7\]
+ _2404_ vssd1 vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__and4_1
XANTENNA__7966__A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5486__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6877_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[10\]
+ _2680_ vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9596_ net460 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5828_ _1778_ _1780_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8616_ net178 _4090_ vssd1 vssd1 vccd1 vccd1 _4095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4915__A2 _0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5759_ _1661_ _1709_ _1711_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__a21oi_1
XANTENNA__7972__Y _3511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8547_ _4015_ _4024_ _4025_ vssd1 vssd1 vccd1 vccd1 _4026_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8478_ _3956_ _3957_ _3330_ vssd1 vssd1 vccd1 vccd1 _3958_ sky130_fd_sc_hd__a21oi_1
XANTENNA__7865__B2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7429_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[2\]
+ _3072_ _3071_ vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_9_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4549__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8409__A3 _3888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8290__A1 _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8037__A team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9280__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8042__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5396__A _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6356__A1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6356__B2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8502__C1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9368__RESET_B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7084__A2 _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8033__A1 _0505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6800_ net519 _2630_ _2632_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__a21oi_1
X_4992_ _0942_ _0944_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_86_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7780_ _3176_ _3368_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6731_ _2586_ _2587_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9327__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6347__A1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6662_ net286 net283 _2532_ _2536_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__and4_1
X_9450_ clknet_leaf_45_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[4\]
+ net237 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5613_ _1087_ _1554_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__xor2_1
X_9381_ clknet_leaf_32_wb_clk_i _0328_ net247 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_8401_ net174 _3869_ vssd1 vssd1 vccd1 vccd1 _3882_ sky130_fd_sc_hd__nor2_1
X_8332_ _0505_ _3821_ vssd1 vssd1 vccd1 vccd1 _3823_ sky130_fd_sc_hd__nand2_1
X_6593_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[10\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[11\]
+ _2493_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5544_ _1449_ _1496_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6849__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5475_ _1363_ _1380_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__xnor2_4
X_8263_ _0494_ _3490_ vssd1 vssd1 vccd1 vccd1 _3758_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8194_ net576 _0456_ _2532_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__a21o_1
X_7214_ net334 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9014__Q team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7145_ _2861_ _2871_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5086__A1 _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7076_ team_08_WB.instance_to_wrap.allocation.game.controller.color\[11\] _2796_
+ _2800_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__a22o_1
X_6027_ _1940_ _1978_ _1979_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout182_X net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7696__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7978_ _0488_ _3484_ _3501_ _3515_ vssd1 vssd1 vccd1 vccd1 _3516_ sky130_fd_sc_hd__a211o_1
XANTENNA__5928__B _1867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6929_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[0\]
+ net554 _2717_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_25_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6338__A1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout98 _3268_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_2
X_9579_ net443 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_91_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout95_X net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6015__A _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8819__A2_N net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5854__A _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload24 clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_6
Xclkload13 clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_11_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload35 clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload46 clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__inv_12
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5260_ _1210_ _1212_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5191_ _1142_ _1143_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__nor2_1
XANTENNA__7057__A2 _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8254__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8079__B1_N team_08_WB.instance_to_wrap.allocation.game.controller.state\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8950_ _3864_ _4115_ _4128_ _4426_ vssd1 vssd1 vccd1 vccd1 _4427_ sky130_fd_sc_hd__and4_1
X_7901_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.state\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.state\[1\] vssd1
+ vssd1 vccd1 vccd1 _3450_ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_8881_ _3816_ _4232_ _4358_ vssd1 vssd1 vccd1 vccd1 _4359_ sky130_fd_sc_hd__o21a_1
XANTENNA__8557__A2 _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7832_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[2\]
+ _3393_ _3395_ vssd1 vssd1 vccd1 vccd1 _3402_ sky130_fd_sc_hd__a21o_1
XANTENNA__8405__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4975_ _0731_ _0732_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__xor2_4
XANTENNA__4652__B team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7763_ net105 _3352_ vssd1 vssd1 vccd1 vccd1 _3353_ sky130_fd_sc_hd__nor2_1
X_6714_ net535 _2573_ net268 vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__o21ai_1
X_9502_ net377 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9433_ clknet_leaf_47_wb_clk_i _0378_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_7694_ net192 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3284_ sky130_fd_sc_hd__or2_4
Xclkload7 clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_6
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6645_ net652 _2528_ net259 vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__o21ai_1
X_9364_ clknet_leaf_26_wb_clk_i _0312_ net250 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6576_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[5\] _2484_ vssd1
+ vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5527_ _1472_ _1474_ _1478_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_9295_ clknet_leaf_12_wb_clk_i _0114_ net217 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_8315_ _3544_ _3806_ net193 vssd1 vssd1 vccd1 vccd1 _3807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9219__RESET_B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8246_ net255 net269 _3744_ vssd1 vssd1 vccd1 vccd1 _3745_ sky130_fd_sc_hd__a21oi_1
X_9472__347 vssd1 vssd1 vccd1 vccd1 _9472__347/HI net347 sky130_fd_sc_hd__conb_1
X_5458_ _0867_ _1215_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__nand2_1
XANTENNA__4645__A_N team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5389_ _1292_ _1341_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout211 net212 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_4
X_8177_ _0691_ _3642_ _0692_ vssd1 vssd1 vccd1 vccd1 _3695_ sky130_fd_sc_hd__a21bo_1
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_4
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_4
Xfanout233 net234 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_4
Xfanout244 net253 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
X_7128_ _2852_ _2858_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__or2_1
Xfanout266 net88 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_2
X_9513__388 vssd1 vssd1 vccd1 vccd1 _9513__388/HI net388 sky130_fd_sc_hd__conb_1
X_7059_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[1\] _0436_
+ _2777_ _2775_ vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__a41o_1
Xfanout277 _0637_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
Xfanout299 team_08_WB.instance_to_wrap.allocation.game.controller.state\[2\] vssd1
+ vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_4
Xfanout288 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[5\] vssd1
+ vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_2
XANTENNA__5004__A _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8985__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8787__A2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4760_ _0713_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4691_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__and2_2
XFILLER_0_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6430_ _2344_ _2379_ vssd1 vssd1 vccd1 vccd1 _2380_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6361_ net333 _2311_ vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5312_ _1210_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8100_ _0686_ _3614_ vssd1 vssd1 vccd1 vccd1 _3628_ sky130_fd_sc_hd__nor2_1
X_6292_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[9\]
+ _2213_ _2216_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[8\]
+ _2244_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__o221a_1
X_9080_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[10\]
+ net222 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8475__A1 _3305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5243_ _1151_ _1195_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__or2_2
X_8031_ _3518_ _3566_ _0481_ vssd1 vssd1 vccd1 vccd1 _3567_ sky130_fd_sc_hd__a21o_1
X_5174_ _1124_ _1126_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__nand2_1
XANTENNA__7304__A _2972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[3\] vssd1
+ vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8778__A2 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7023__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8933_ _0405_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[0\] team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _4410_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8864_ _4334_ _4340_ _4341_ vssd1 vssd1 vccd1 vccd1 _4342_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7815_ net293 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _3392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8795_ net186 _4270_ _4272_ vssd1 vssd1 vccd1 vccd1 _4273_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4958_ net145 _0909_ _0809_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout145_X net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7746_ _3315_ _3335_ vssd1 vssd1 vccd1 vccd1 _3336_ sky130_fd_sc_hd__nand2_1
X_4889_ _0834_ _0840_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7677_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[5\]
+ net106 _3263_ vssd1 vssd1 vccd1 vccd1 _3267_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6628_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[24\] _2518_
+ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__and2_1
X_9416_ clknet_leaf_43_wb_clk_i _0361_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9347_ clknet_leaf_46_wb_clk_i _0295_ net233 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_9554__422 vssd1 vssd1 vccd1 vccd1 _9554__422/HI net422 sky130_fd_sc_hd__conb_1
XFILLER_0_30_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6559_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[3\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[2\]
+ _2472_ _2473_ vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__or4_1
X_9278_ clknet_leaf_5_wb_clk_i _0106_ net214 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6477__B1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8229_ _3027_ _3712_ vssd1 vssd1 vccd1 vccd1 _3733_ sky130_fd_sc_hd__or2_1
XANTENNA__7214__A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_1__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8045__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4573__A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8154__B1 _3608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4748__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5930_ _0718_ net146 _1882_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5861_ _0919_ _1813_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8932__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7600_ _3188_ _3189_ vssd1 vssd1 vccd1 vccd1 _3190_ sky130_fd_sc_hd__nor2_1
XANTENNA__7735__A3 _3261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4812_ _0762_ _0764_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__xnor2_4
X_5792_ net168 net145 vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8580_ _4038_ _4051_ _4057_ _4058_ vssd1 vssd1 vccd1 vccd1 _4059_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4743_ _0688_ _0696_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7531_ net514 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet vssd1 vssd1
+ vccd1 vccd1 _0251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7462_ net302 net305 _0441_ _3045_ vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9201_ clknet_leaf_15_wb_clk_i _0022_ net217 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_4674_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[7\] vssd1
+ vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__nand2b_1
X_6413_ _2354_ _2363_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__nand2_1
X_7393_ _3034_ _3039_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6344_ _2293_ _2295_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9132_ clknet_leaf_41_wb_clk_i _0233_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout105_A _3271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6275_ _2108_ _2227_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__nand2_1
X_9063_ clknet_leaf_33_wb_clk_i _0198_ net247 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_5226_ net123 _1170_ _1172_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__o21ai_1
X_8014_ _3523_ _3550_ vssd1 vssd1 vccd1 vccd1 _3551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5157_ _1095_ _1109_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__and2_1
X_9584__448 vssd1 vssd1 vccd1 vccd1 _9584__448/HI net448 sky130_fd_sc_hd__conb_1
X_5088_ _0863_ _0875_ _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__o21bai_2
XANTENNA__7688__B net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6631__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8916_ _4389_ _4390_ _4392_ vssd1 vssd1 vccd1 vccd1 _4393_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8847_ _4292_ _4324_ vssd1 vssd1 vccd1 vccd1 _4325_ sky130_fd_sc_hd__nand2_1
XANTENNA__4680__X _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8778_ net313 _0520_ _4232_ _4255_ vssd1 vssd1 vccd1 vccd1 _4256_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8923__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4840__B net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5936__B _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7729_ _3294_ _3307_ vssd1 vssd1 vccd1 vccd1 _3319_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6698__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9478__353 vssd1 vssd1 vccd1 vccd1 _9478__353/HI net353 sky130_fd_sc_hd__conb_1
XFILLER_0_34_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9519__394 vssd1 vssd1 vccd1 vccd1 _9519__394/HI net394 sky130_fd_sc_hd__conb_1
XFILLER_0_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input35_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6007__B _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8678__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8678__B2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6060_ _1998_ _2011_ _2012_ vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__and3_1
X_5011_ _0767_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7301__B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6613__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6962_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[15\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[14\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[13\]
+ _2733_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__and4_1
X_5913_ _1863_ _1864_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__xnor2_1
X_6893_ net270 _2692_ _2694_ _2695_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_0__f_wb_clk_i_X clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_8701_ _4179_ vssd1 vssd1 vccd1 vccd1 _4180_ sky130_fd_sc_hd__inv_2
X_5844_ _1790_ _1796_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8632_ _4109_ _4110_ vssd1 vssd1 vccd1 vccd1 _4111_ sky130_fd_sc_hd__nor2_1
XANTENNA__5756__B _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8563_ net127 _3619_ _4041_ net136 vssd1 vssd1 vccd1 vccd1 _4042_ sky130_fd_sc_hd__o22a_1
X_5775_ _1726_ _1727_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__and2_1
X_7514_ net310 _3040_ vssd1 vssd1 vccd1 vccd1 _3149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4726_ net282 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout222_A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8494_ net171 net116 _3318_ _3343_ _3346_ vssd1 vssd1 vccd1 vccd1 _3974_ sky130_fd_sc_hd__a41o_1
X_4657_ _0613_ _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__nand2b_2
XANTENNA__9017__Q team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7445_ net523 net115 _3070_ _3088_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7376_ net302 net301 _3025_ _3023_ vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4588_ _0419_ _0553_ _0420_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[0\]
+ sky130_fd_sc_hd__o21a_1
X_9115_ clknet_leaf_46_wb_clk_i _0218_ net234 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_6327_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[5\] _2273_ vssd1
+ vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout108_X net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9069__SET_B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6258_ _0444_ _2210_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9046_ clknet_leaf_37_wb_clk_i _0181_ net248 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6189_ _1394_ _2141_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__and2b_1
X_5209_ _1160_ _1161_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9233__CLK clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8109__B1 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7580__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4585__X _0551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4745__B _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Left_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8899__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5560_ _1511_ _1512_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__nand2b_1
X_4511_ team_08_WB.EN_VAL_REG net38 _0480_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__mux2_1
X_5491_ _1405_ _1443_ vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6688__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7791__B team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5592__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[0\]
+ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold116 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__dlygate4sd3_1
X_7230_ net648 _2924_ net181 vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8520__B1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold127 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.clk1
+ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[0\]
+ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[2\] vssd1 vssd1
+ vccd1 vccd1 net636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7161_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[2\] _2877_ vssd1
+ vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6112_ _2054_ _2063_ _2064_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__nand3_1
X_7092_ _2825_ _2831_ _2832_ _2775_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__o31a_1
XFILLER_0_42_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6043_ _1994_ _1995_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7994_ _0485_ _3521_ _3522_ _3530_ vssd1 vssd1 vccd1 vccd1 _3532_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_53_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout172_A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6945_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[9\]
+ _2725_ vssd1 vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__or2_1
XANTENNA__8414__Y _3895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6876_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[10\]
+ _2680_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9595_ net459 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
X_5827_ _1726_ _1732_ _1779_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8615_ net162 net169 _4093_ vssd1 vssd1 vccd1 vccd1 _4094_ sky130_fd_sc_hd__and3_1
X_5758_ net141 _0928_ _0931_ net140 vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout225_X net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8546_ net118 _3674_ vssd1 vssd1 vccd1 vccd1 _4025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_62_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4709_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[4\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_20_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8477_ net186 _3284_ _3921_ net189 vssd1 vssd1 vccd1 vccd1 _3957_ sky130_fd_sc_hd__or4b_1
X_5689_ _1640_ _1641_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__nand2_1
X_7428_ net310 _0442_ vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7359_ net606 _2974_ _3013_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__o21a_1
XANTENNA__4549__C net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6825__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9029_ clknet_leaf_53_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[11\]
+ net200 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__7222__A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8053__A _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5619__A1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4991_ net128 _0941_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_86_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6730_ net679 _2585_ net267 vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4491__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7792__A1 _2368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6347__A2 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6661_ _2539_ _2540_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5612_ _0826_ _1556_ _1564_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9380_ clknet_leaf_31_wb_clk_i _0327_ net244 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6592_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[9\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[10\]
+ _2492_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[11\] vssd1
+ vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__a31o_1
X_8400_ net175 net151 vssd1 vssd1 vccd1 vccd1 _3881_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5543_ _1447_ _1448_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8331_ _0505_ _3821_ vssd1 vssd1 vccd1 vccd1 _3822_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__6849__C _2665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5474_ _1424_ _1426_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__nand2_1
XANTENNA__6211__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8262_ net139 _2267_ vssd1 vssd1 vccd1 vccd1 _3757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7026__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8193_ _3597_ _3705_ _3709_ net244 net595 vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__o32a_1
X_7213_ net329 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7144_ net184 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[11\]
+ _2850_ _2872_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__a31o_1
XANTENNA__4666__A team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7075_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[3\]
+ _2792_ _2809_ team_08_WB.instance_to_wrap.allocation.game.controller.color\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__a22o_1
X_6026_ _1937_ _1938_ _1939_ _1887_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__a22oi_1
XANTENNA__7480__B1 _3110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7977__A _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9078__RESET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7696__B _3261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7977_ _0422_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 _3515_ sky130_fd_sc_hd__nor2_1
XANTENNA__7783__B2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7783__A1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5794__B1 _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6928_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[0\]
+ net554 net158 vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4597__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6859_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[4\]
+ _2670_ _2672_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout99 _3266_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_4
XFILLER_0_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9578_ team_08_WB.instance_to_wrap.allocation.game.collides vssd1 vssd1 vccd1 vccd1
+ net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8529_ _3261_ _4004_ _4007_ vssd1 vssd1 vccd1 vccd1 _4008_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_92_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5849__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5959__X _1912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5200__A _0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4588__A1 _0419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6015__B _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8723__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5854__B _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6332__A1_N net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload25 clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload14 clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload47 clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__inv_8
XFILLER_0_3_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload36 clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_23_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5190_ _1141_ _1140_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__and2b_1
X_7900_ _3449_ _3447_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[20\]
+ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__mux2_1
X_8880_ net320 _4232_ net316 vssd1 vssd1 vccd1 vccd1 _4358_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7831_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\]
+ _3395_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__and2_1
X_4974_ _0926_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__inv_2
XANTENNA__6206__A _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7762_ net191 _3351_ vssd1 vssd1 vccd1 vccd1 _3352_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6713_ _2573_ _2574_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9501_ net376 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XANTENNA__7517__A1 _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_7693_ _0556_ net97 _3278_ net100 vssd1 vssd1 vccd1 vccd1 _3283_ sky130_fd_sc_hd__o31a_1
X_9432_ clknet_leaf_29_wb_clk_i _0377_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6644_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[30\] _2528_
+ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload8 clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_6
XFILLER_0_34_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout135_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8421__A _3279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9363_ clknet_leaf_26_wb_clk_i _0311_ net250 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6575_ _2484_ _2485_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5483__C _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5526_ _1472_ _1474_ _1478_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_70_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9294_ clknet_leaf_13_wb_clk_i _0113_ net217 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_8314_ _0483_ _3805_ vssd1 vssd1 vccd1 vccd1 _3806_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5457_ _1366_ _1409_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__and2_2
XFILLER_0_30_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8245_ _2331_ _3742_ _3743_ net259 vssd1 vssd1 vccd1 vccd1 _3744_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5388_ _1281_ _1284_ _1291_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__nand3_1
Xfanout212 net232 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_2
Xfanout223 net231 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_4
X_8176_ _3693_ _3694_ net685 net244 vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout201 net206 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_4
Xfanout234 net236 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
Xfanout245 net248 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_4
Xfanout256 _0515_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_2
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7127_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\]
+ _2853_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__nor2_1
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
Xfanout289 team_08_WB.instance_to_wrap.allocation.game.controller.v\[4\] vssd1 vssd1
+ vccd1 vccd1 net289 sky130_fd_sc_hd__buf_2
X_7058_ _2775_ _2786_ _2802_ _2805_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__o22a_1
Xfanout278 _0637_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_2
X_6009_ net167 _0926_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5020__A _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8331__A _0505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7444__B1 _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7995__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8065__X _3597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5758__B1 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8172__B2 _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4690_ _0640_ _0643_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6360_ net335 team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[0\] _2311_
+ net333 vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5311_ _1193_ _1209_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6291_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[8\]
+ _2216_ _2243_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__a21oi_1
X_8030_ _0482_ _0498_ vssd1 vssd1 vccd1 vccd1 _3566_ sky130_fd_sc_hd__nor2_1
XANTENNA__6486__A1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5242_ _0856_ _1150_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__nor2_1
X_5173_ _1113_ _1121_ _1123_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__or3_1
Xinput1 gpio_in[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
X_8932_ _2294_ net98 _3265_ vssd1 vssd1 vccd1 vccd1 _4409_ sky130_fd_sc_hd__a21oi_1
X_8863_ _4334_ _4340_ _3271_ vssd1 vssd1 vccd1 vccd1 _4341_ sky130_fd_sc_hd__a21o_1
XANTENNA__5478__C _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7814_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[5\] _2975_ _3387_
+ _3390_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__a22o_1
XANTENNA__8935__B1 _3284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8794_ net185 _4270_ _4271_ vssd1 vssd1 vccd1 vccd1 _4272_ sky130_fd_sc_hd__a21bo_1
X_4957_ _0736_ _0737_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7745_ net110 _3241_ _3305_ vssd1 vssd1 vccd1 vccd1 _3335_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4888_ _0834_ _0840_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7676_ _3257_ _3264_ _3259_ vssd1 vssd1 vccd1 vccd1 _3266_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9415_ clknet_leaf_43_wb_clk_i _0360_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_6627_ _2518_ net260 _2517_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[23\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__7990__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9346_ clknet_leaf_46_wb_clk_i _0294_ net235 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_6558_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5509_ _0814_ net145 _1461_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__and3_1
X_9277_ clknet_leaf_18_wb_clk_i _0276_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.clk1
+ sky130_fd_sc_hd__dfxtp_1
X_6489_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[6\] team_08_WB.instance_to_wrap.allocation.game.controller.state\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__or2_4
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8228_ _2992_ _3731_ net121 vssd1 vssd1 vccd1 vccd1 _3732_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7989__X _3527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8159_ net286 _2388_ vssd1 vssd1 vccd1 vccd1 _3679_ sky130_fd_sc_hd__or2_1
XANTENNA__9093__RESET_B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5015__A _0744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9022__RESET_B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8326__A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4860__Y _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8154__B2 _2393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7665__B1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6963__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6308__X _2261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5860_ _1810_ _1811_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7584__A1_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4811_ net168 _0756_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5791_ _0743_ _1743_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4770__Y _0723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4742_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__inv_2
X_7530_ net505 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet vssd1 vssd1
+ vccd1 vccd1 _0250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4673_ _0608_ _0630_ _0607_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_32_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7461_ net302 _3099_ _3101_ _0438_ vssd1 vssd1 vccd1 vccd1 _3103_ sky130_fd_sc_hd__o31a_1
XFILLER_0_16_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9200_ clknet_leaf_16_wb_clk_i _0034_ net217 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_6412_ _2362_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7392_ _3032_ _3037_ net500 vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4939__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6343_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[5\] _2292_ vssd1
+ vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__nand2_1
X_9131_ clknet_leaf_41_wb_clk_i _0232_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_6274_ _2106_ _2107_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__nand2_1
X_9062_ clknet_leaf_33_wb_clk_i _0197_ net247 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_5225_ _1167_ _1175_ _1177_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__o21ai_1
X_8013_ _3548_ _3549_ vssd1 vssd1 vccd1 vccd1 _3550_ sky130_fd_sc_hd__or2_1
XANTENNA__4658__B team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5156_ _1104_ _1107_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7959__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5087_ _0850_ _0875_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__and2b_1
X_8915_ _4008_ _4386_ _4391_ vssd1 vssd1 vccd1 vccd1 _4392_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8846_ _4293_ _4295_ vssd1 vssd1 vccd1 vccd1 _4324_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _1907_ _1940_ _1941_ vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__nand3_1
X_8777_ _4237_ _4251_ _4254_ _4249_ vssd1 vssd1 vccd1 vccd1 _4255_ sky130_fd_sc_hd__o22a_1
X_7728_ net112 net109 _3305_ vssd1 vssd1 vccd1 vccd1 _3318_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7659_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[7\]
+ _3227_ net110 _3226_ vssd1 vssd1 vccd1 vccd1 _3249_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9329_ clknet_leaf_0_wb_clk_i _0012_ net200 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5122__A1 _0919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8608__X _4087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input28_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8375__B2 team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8678__A2 _3622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5010_ _0961_ _0962_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__or2_1
XANTENNA__8850__A2 _3888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4765__Y _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6961_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[14\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[13\]
+ _2733_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__a31o_1
X_8700_ net176 _4175_ _4178_ net150 vssd1 vssd1 vccd1 vccd1 _4179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5912_ _1863_ _1864_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__and2b_1
X_6892_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5843_ _1792_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8631_ _2534_ net113 vssd1 vssd1 vccd1 vccd1 _4110_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8562_ _4039_ _4040_ vssd1 vssd1 vccd1 vccd1 _4041_ sky130_fd_sc_hd__nor2_1
X_5774_ _1675_ _1725_ _1724_ _1708_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__a211o_1
X_7513_ _3023_ _3032_ _3038_ _3066_ _3148_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__a41o_1
XFILLER_0_12_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4725_ _0678_ _0679_ _0676_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__o21a_1
X_8493_ _3866_ _3904_ _3881_ _3366_ vssd1 vssd1 vccd1 vccd1 _3973_ sky130_fd_sc_hd__o211a_1
XANTENNA__7877__B1 _3403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4656_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[4\] vssd1
+ vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7444_ _3083_ _3087_ _3023_ vssd1 vssd1 vccd1 vccd1 _3088_ sky130_fd_sc_hd__a21oi_1
X_4587_ net334 _0546_ _0552_ _0540_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7375_ net307 net304 vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9114_ clknet_leaf_46_wb_clk_i _0217_ net234 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6326_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[5\] _2273_ vssd1
+ vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6257_ _1996_ _2120_ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4956__X _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9045_ clknet_leaf_37_wb_clk_i net553 net248 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_6188_ _1391_ _1393_ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__or2_1
X_5208_ _1155_ _1157_ _1159_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7699__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5139_ _0749_ _0805_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8054__B1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8829_ net317 net95 _4306_ vssd1 vssd1 vccd1 vccd1 _4307_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8348__A1 _3511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5264__A1_N _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9196__RESET_B net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4510_ net39 net37 net40 _0479_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__and4_1
X_5490_ _0748_ _1404_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[0\]
+ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7160_ net164 _2877_ _2878_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold128 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[5\] vssd1
+ vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6111_ _2051_ _2053_ _2052_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__a21o_1
X_7091_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[7\]
+ _2789_ _2800_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6042_ _1992_ _1993_ vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__nor2_1
XANTENNA__8587__A1 _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7993_ _3523_ _3530_ vssd1 vssd1 vccd1 vccd1 _3531_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout165_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6944_ _2725_ net158 _2724_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__and3b_1
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_92_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6875_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[10\]
+ _2680_ _2682_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8614_ _0696_ _3178_ vssd1 vssd1 vccd1 vccd1 _4093_ sky130_fd_sc_hd__xnor2_1
X_9594_ net458 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_92_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5826_ _1726_ _1733_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout332_A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5757_ _0813_ _0926_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8545_ net127 _3685_ _4023_ vssd1 vssd1 vccd1 vccd1 _4024_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4708_ _0656_ _0660_ _0658_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout120_X net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8476_ _3273_ _3281_ _3351_ _3279_ vssd1 vssd1 vccd1 vccd1 _3956_ sky130_fd_sc_hd__a31o_1
X_5688_ _1638_ _1639_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7427_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[2\]
+ _0441_ vssd1 vssd1 vccd1 vccd1 _3071_ sky130_fd_sc_hd__nand2_2
XANTENNA__8511__A1 _3280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4639_ _0582_ _0596_ _0581_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_9_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7358_ _2975_ _3011_ _3014_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_9_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5007__B _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6309_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[2\]
+ _0635_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__nand2_1
X_7289_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[21\]
+ _2964_ net181 vssd1 vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9028_ clknet_leaf_53_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[10\]
+ net207 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5023__A _0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8578__A1 _3241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5958__A _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4846__A_N _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6029__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9401__Q team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8569__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5868__A _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4990_ _0915_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_86_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6660_ net286 _2532_ _2538_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__o21ai_1
X_5611_ _1563_ _1562_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6591_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[10\] _2493_
+ _2495_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5542_ _1494_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8330_ _3566_ _3792_ _0481_ vssd1 vssd1 vccd1 vccd1 _3821_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5473_ _1408_ _1425_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8261_ _3755_ _3756_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[1\]
+ net235 vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7212_ net313 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8192_ _0654_ _3706_ _3708_ _3704_ vssd1 vssd1 vccd1 vccd1 _3709_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7143_ _2862_ _2869_ _2871_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7074_ _2811_ _2814_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__nand2b_1
XANTENNA__4666__B team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6025_ _1975_ _1977_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7977__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout168_X net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7976_ net325 _2426_ net277 vssd1 vssd1 vccd1 vccd1 _3514_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7783__A2 _2325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5794__B2 _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6927_ net600 _0019_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__nor2_1
XANTENNA__4597__A2 team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9646_ net264 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6858_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[4\]
+ _2670_ net273 vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9047__RESET_B net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9577_ net442 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_92_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5809_ _1759_ _1760_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__xor2_1
X_6789_ net637 _2624_ net270 vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__o21ai_1
XANTENNA__7057__X _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8528_ _4005_ _4006_ vssd1 vssd1 vccd1 vccd1 _4007_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8459_ _3867_ _3923_ _3932_ _3939_ vssd1 vssd1 vccd1 vccd1 _3940_ sky130_fd_sc_hd__a31oi_1
XANTENNA__5849__A2 _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8248__A0 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8799__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8799__B2 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5482__B1 _1434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input10_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7774__A2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8723__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload26 clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_4
XTAP_TAPCELL_ROW_11_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload15 clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload48 clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload37 clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8239__A _3034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7830_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[3\]
+ _3400_ _3401_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__a22o_1
XANTENNA__8411__B1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4973_ _0729_ _0925_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__or2_4
X_7761_ net188 net185 vssd1 vssd1 vccd1 vccd1 _3351_ sky130_fd_sc_hd__or2_1
X_6712_ net623 _2572_ net268 vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7692_ net100 net95 vssd1 vssd1 vccd1 vccd1 _3282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9500_ net375 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_50_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9431_ clknet_leaf_1_wb_clk_i _0376_ net211 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6643_ _2528_ net260 _2527_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[29\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload9 clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_8
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8421__B _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_A _0939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9362_ clknet_leaf_26_wb_clk_i _0310_ net250 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6574_ net659 _2482_ net263 vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5525_ _1476_ _1477_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__and2_1
X_9293_ clknet_leaf_13_wb_clk_i _0112_ net218 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_8313_ _0498_ _3792_ vssd1 vssd1 vccd1 vccd1 _3805_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_48_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5456_ _1217_ _1365_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8244_ team_08_WB.instance_to_wrap.allocation.game.game.score\[6\] team_08_WB.instance_to_wrap.allocation.game.game.score\[5\]
+ _2326_ _2332_ vssd1 vssd1 vccd1 vccd1 _3743_ sky130_fd_sc_hd__nand4_1
XFILLER_0_30_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5387_ _1337_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__nand2_1
Xfanout213 net216 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4677__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8175_ _0701_ _3687_ _3691_ net244 vssd1 vssd1 vccd1 vccd1 _3694_ sky130_fd_sc_hd__o211a_1
Xfanout202 net206 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_4
Xfanout224 net231 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_4
Xfanout246 net248 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_4
X_7126_ _2854_ _2856_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__nand2_1
Xfanout268 _2548_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_2
X_7057_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[0\]
+ _2800_ _2803_ _2804_ vssd1 vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__a211o_1
XANTENNA_input2_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout279 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[8\] vssd1
+ vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6008_ _0724_ _0929_ _1960_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__or3_1
XANTENNA__9119__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9299__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9228__RESET_B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7756__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7959_ net297 _3489_ _3497_ _3498_ vssd1 vssd1 vccd1 vccd1 _3499_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8612__A _0674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9629_ net266 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_42_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5971__A _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8944__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5758__B2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5310_ _1251_ _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__nor2_1
X_6290_ _2218_ _2240_ _2241_ _2242_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5241_ _0758_ _0785_ _1045_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__a21oi_4
XANTENNA__8880__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4497__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5172_ net123 _1116_ _1118_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_20_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput2 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_8931_ _2280_ _3329_ _4372_ _4378_ _4407_ vssd1 vssd1 vccd1 vccd1 _4408_ sky130_fd_sc_hd__o221a_1
X_8862_ _4227_ _4228_ _4338_ _4339_ _4336_ vssd1 vssd1 vccd1 vccd1 _4340_ sky130_fd_sc_hd__o32a_1
XANTENNA__8935__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7813_ net689 _2974_ _3389_ _3391_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__o211a_1
X_8793_ _4230_ _4218_ _4219_ vssd1 vssd1 vccd1 vccd1 _4271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7744_ net188 _0425_ _0555_ _3333_ _3332_ vssd1 vssd1 vccd1 vccd1 _3334_ sky130_fd_sc_hd__o41ai_2
XANTENNA__8432__A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ _0736_ _0737_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__xor2_4
XFILLER_0_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout245_A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4887_ net143 _0839_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__xnor2_1
X_7675_ _3257_ _3264_ _3259_ vssd1 vssd1 vccd1 vccd1 _3265_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_85_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9414_ clknet_leaf_43_wb_clk_i _0359_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_6626_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[23\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[22\]
+ _2514_ vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__and3_1
XANTENNA__7990__B _3527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9345_ clknet_leaf_47_wb_clk_i _0293_ net224 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6557_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[5\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[6\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__or4b_1
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5791__A _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5508_ net140 _0910_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9276_ clknet_leaf_20_wb_clk_i _0275_ net241 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr2\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_6488_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[6\] team_08_WB.instance_to_wrap.allocation.game.controller.state\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__nor2_2
XFILLER_0_30_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5439_ net129 _1344_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__or2_1
X_8227_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[13\]
+ _2991_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[14\]
+ vssd1 vssd1 vccd1 vccd1 _3731_ sky130_fd_sc_hd__o21ai_1
X_8158_ _2321_ _3677_ vssd1 vssd1 vccd1 vccd1 _3678_ sky130_fd_sc_hd__and2_1
XANTENNA_input5_X net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7109_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[6\] _2842_
+ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__and3_1
X_8089_ _0706_ net178 vssd1 vssd1 vccd1 vccd1 _3618_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_2_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6346__A1_N net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5206__A _1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9434__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7421__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7778__D _3367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9462__337 vssd1 vssd1 vccd1 vccd1 _9462__337/HI net337 sky130_fd_sc_hd__conb_1
XFILLER_0_75_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4810_ _0740_ _0756_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__nor2_1
XANTENNA__6928__B1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5790_ _1697_ _1698_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4741_ _0694_ _0695_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__and2_4
XFILLER_0_28_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4672_ _0611_ _0629_ _0610_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9503__378 vssd1 vssd1 vccd1 vccd1 _9503__378/HI net378 sky130_fd_sc_hd__conb_1
X_7460_ net302 _3101_ _3099_ vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6411_ _2344_ _2350_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7391_ _3037_ vssd1 vssd1 vccd1 vccd1 _3038_ sky130_fd_sc_hd__inv_2
X_9130_ clknet_leaf_41_wb_clk_i _0231_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6342_ _2293_ vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__inv_2
X_6273_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[4\]
+ _2225_ vssd1 vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9061_ clknet_leaf_33_wb_clk_i _0196_ net247 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8853__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5224_ _1121_ _1176_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__nor2_1
X_8012_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] _3543_ vssd1
+ vssd1 vccd1 vccd1 _3549_ sky130_fd_sc_hd__and2_1
X_5155_ _1104_ _1107_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout195_A _3460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5086_ _0826_ _1010_ _1009_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__a21o_2
XFILLER_0_79_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8914_ _0689_ net118 _4385_ vssd1 vssd1 vccd1 vccd1 _4391_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8845_ _4300_ _4319_ _4322_ _4315_ vssd1 vssd1 vccd1 vccd1 _4323_ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5988_ _1903_ _1904_ _1906_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout248_X net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8776_ _4241_ _4253_ _4240_ vssd1 vssd1 vccd1 vccd1 _4254_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4939_ net143 _0839_ _0890_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__and3_1
X_7727_ net171 _3313_ _3315_ _3316_ vssd1 vssd1 vccd1 vccd1 _3317_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7658_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[5\]
+ _3238_ _3247_ vssd1 vssd1 vccd1 vccd1 _3248_ sky130_fd_sc_hd__and3_1
X_6609_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[17\] _2505_
+ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7589_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[16\]
+ _2855_ _3177_ vssd1 vssd1 vccd1 vccd1 _3179_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_63_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9328_ clknet_leaf_30_wb_clk_i _0011_ net238 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9259_ clknet_leaf_10_wb_clk_i _0077_ net227 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4584__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5696__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8800__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8850__A3 _3895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4872__A1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8249__A2_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6960_ _0462_ _2734_ _2735_ net158 vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9544__412 vssd1 vssd1 vccd1 vccd1 _9544__412/HI net412 sky130_fd_sc_hd__conb_1
XFILLER_0_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5911_ _1814_ _1815_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6891_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5842_ _1792_ _1793_ _1794_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__nand3_1
X_8630_ _2533_ net111 vssd1 vssd1 vccd1 vccd1 _4109_ sky130_fd_sc_hd__nor2_1
X_5773_ _1708_ _1724_ _1725_ _1675_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8561_ net169 _3618_ vssd1 vssd1 vccd1 vccd1 _4040_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4724_ _0672_ _0673_ _0670_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__o21a_2
XFILLER_0_29_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7512_ _0134_ _3147_ vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__nor2_1
X_8492_ _3966_ _3968_ _3971_ _3283_ vssd1 vssd1 vccd1 vccd1 _3972_ sky130_fd_sc_hd__o211a_1
X_4655_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[4\] vssd1
+ vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7443_ net310 net308 _3024_ _3077_ _3086_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__o311a_1
XFILLER_0_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4586_ _0551_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__inv_2
X_7374_ net303 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout110_A _3235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9590__454 vssd1 vssd1 vccd1 vccd1 _9590__454/HI net454 sky130_fd_sc_hd__conb_1
X_9113_ clknet_leaf_46_wb_clk_i _0216_ net234 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_6325_ net328 _2271_ _2275_ net325 _2272_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__o221a_1
XANTENNA__9314__Q team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9044_ clknet_leaf_35_wb_clk_i _0179_ net246 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6256_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[12\]
+ _2208_ vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6187_ _1442_ _2138_ _1440_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__a21o_1
X_5207_ _1155_ _1157_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_4_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4685__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5138_ _1089_ _1090_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7996__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5069_ _0997_ _1020_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8828_ _4289_ _4303_ _4305_ vssd1 vssd1 vccd1 vccd1 _4306_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8759_ _4220_ _4230_ _4236_ vssd1 vssd1 vccd1 vccd1 _4237_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7583__A1_N net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input40_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4882__X _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7556__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6969__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold107 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[3\]
+ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[12\] vssd1
+ vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.internalSck
+ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__dlygate4sd3_1
X_6110_ _2060_ _2062_ vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__nor2_1
X_9615__479 vssd1 vssd1 vccd1 vccd1 _9615__479/HI net479 sky130_fd_sc_hd__conb_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7090_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[7\]
+ _2792_ _2799_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__a22o_1
XANTENNA__8284__A1 _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6041_ _1992_ _1993_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_47_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_7992_ _3528_ _3529_ vssd1 vssd1 vccd1 vccd1 _3530_ sky130_fd_sc_hd__and2_1
X_9468__343 vssd1 vssd1 vccd1 vccd1 _9468__343/HI net343 sky130_fd_sc_hd__conb_1
X_6943_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[8\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[7\]
+ _2404_ vssd1 vssd1 vccd1 vccd1 _2725_ sky130_fd_sc_hd__and3_1
XANTENNA__5400__Y _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6874_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[10\]
+ _2680_ net273 vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5825_ _1772_ _1775_ _1776_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9509__384 vssd1 vssd1 vccd1 vccd1 _9509__384/HI net384 sky130_fd_sc_hd__conb_1
XFILLER_0_14_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8613_ _0685_ net136 vssd1 vssd1 vccd1 vccd1 _4092_ sky130_fd_sc_hd__xnor2_1
X_9593_ net457 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
XANTENNA__5022__A1 _0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5756_ net141 _0930_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout325_A team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8544_ net136 _4014_ _4021_ _4022_ vssd1 vssd1 vccd1 vccd1 _4023_ sky130_fd_sc_hd__a211o_1
X_5687_ _1639_ _1638_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__nand2b_1
X_4707_ _0656_ _0660_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8475_ _3305_ _3309_ _3886_ _3953_ vssd1 vssd1 vccd1 vccd1 _3955_ sky130_fd_sc_hd__a31o_1
X_4638_ _0593_ _0594_ _0584_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__a21o_2
XFILLER_0_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7426_ net534 net114 _3063_ _3070_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout113_X net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4569_ _0504_ _0505_ _0537_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o21ai_1
X_7357_ net569 _2975_ vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6308_ _2151_ _2178_ _2260_ _2176_ _2177_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__a2111o_4
XTAP_TAPCELL_ROW_90_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7288_ net180 _2963_ _2965_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__and3_1
X_6239_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[20\]
+ _2191_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9027_ clknet_leaf_53_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[9\]
+ net200 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8027__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5958__B _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7002__A2 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6029__B _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6045__A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5610_ _0825_ _1556_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6590_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[10\] _2493_
+ net258 vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5541_ _1491_ _1492_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8260_ net139 _2264_ _2276_ _2311_ net161 vssd1 vssd1 vccd1 vccd1 _3756_ sky130_fd_sc_hd__o32a_1
XFILLER_0_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5472_ _1405_ _1407_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__nand2_1
X_7211_ _0424_ _2909_ _2910_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8191_ _2391_ _3707_ net296 vssd1 vssd1 vccd1 vccd1 _3708_ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7142_ _2862_ _2863_ _2869_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__a21oi_1
X_7073_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[1\]
+ _2777_ _2817_ _2775_ vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6024_ _1885_ _1976_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__nor2_1
XANTENNA__7610__Y _3200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout275_A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7975_ net669 _3513_ net242 vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6926_ net530 _2714_ _2716_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8717__C1 _4087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9645_ net488 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
X_6857_ _0466_ _2668_ _2671_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9039__Q team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoMovement
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9576_ net441 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_91_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5808_ _1760_ _1759_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6788_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[9\]
+ _2624_ vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5739_ _1689_ _1690_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8527_ _0657_ _3241_ vssd1 vssd1 vccd1 vccd1 _4006_ sky130_fd_sc_hd__nand2_1
X_9596__460 vssd1 vssd1 vccd1 vccd1 _9596__460/HI net460 sky130_fd_sc_hd__conb_1
XFILLER_0_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8458_ net154 net94 _3905_ _3332_ vssd1 vssd1 vccd1 vccd1 _3939_ sky130_fd_sc_hd__o211a_1
XANTENNA__8496__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7409_ _0441_ _3051_ vssd1 vssd1 vccd1 vccd1 _3054_ sky130_fd_sc_hd__nor2_1
X_8389_ net175 _3869_ vssd1 vssd1 vccd1 vccd1 _3870_ sky130_fd_sc_hd__nand2_2
XANTENNA__6991__A_N team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4873__A _0825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6417__X _2368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6431__B1 _2325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7774__A3 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_11_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload27 clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_51_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload49 clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload38 clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__inv_8
XFILLER_0_24_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7424__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8411__A1 _0425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4972_ _0625_ _0727_ _0728_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__o21ba_1
X_7760_ _3334_ _3337_ _3341_ _3349_ _3328_ vssd1 vssd1 vccd1 vccd1 _3350_ sky130_fd_sc_hd__a221o_1
XANTENNA__4984__B1 _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6711_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[12\]
+ _2572_ vssd1 vssd1 vccd1 vccd1 _2573_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8175__B1 _3691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7691_ net99 net97 vssd1 vssd1 vccd1 vccd1 _3281_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9430_ clknet_leaf_2_wb_clk_i _0375_ net204 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_6642_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[29\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[28\]
+ _2524_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__and3_1
X_9361_ clknet_leaf_26_wb_clk_i _0309_ net251 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__7922__B1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8312_ net198 _3801_ _3802_ _3803_ vssd1 vssd1 vccd1 vccd1 _3804_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6573_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[3\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[4\]
+ _2481_ vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5524_ _1450_ _1451_ _1475_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9292_ clknet_leaf_14_wb_clk_i _0111_ net215 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5455_ _1405_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8243_ team_08_WB.instance_to_wrap.allocation.game.game.score\[2\] team_08_WB.instance_to_wrap.allocation.game.game.score\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.game.score\[4\] team_08_WB.instance_to_wrap.allocation.game.game.score\[3\]
+ vssd1 vssd1 vccd1 vccd1 _3742_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8174_ _0709_ _3692_ net137 vssd1 vssd1 vccd1 vccd1 _3693_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5386_ _1327_ _1330_ _1337_ _1338_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__o211ai_2
Xfanout214 net216 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4677__B _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout203 net206 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
X_7125_ _2851_ _2855_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__nand2_1
Xfanout225 net231 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
Xfanout247 net248 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_4
Xfanout236 net254 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
XANTENNA__9322__Q team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8717__X _4196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4964__Y _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7056_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[0\]
+ _2792_ _2796_ team_08_WB.instance_to_wrap.allocation.game.controller.color\[8\]
+ _2801_ vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__a221o_1
Xfanout269 _2548_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_4
Xfanout258 _0515_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_4
XANTENNA__8650__A1 _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6007_ _0718_ _0930_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7958_ net330 _2426_ net277 vssd1 vssd1 vccd1 vccd1 _3498_ sky130_fd_sc_hd__a21o_1
X_7889_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[17\]
+ _3439_ net160 vssd1 vssd1 vccd1 vccd1 _3442_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6909_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[7\]
+ _2704_ net272 vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8612__B _3214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9628_ net266 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_42_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9559_ net427 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_0_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8469__A1 _3279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _1145_ _1192_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__and2_1
XANTENNA__7154__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8880__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5171_ _1113_ _1121_ _1123_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8930_ _4400_ _4403_ _4404_ _4405_ _4393_ vssd1 vssd1 vccd1 vccd1 _4407_ sky130_fd_sc_hd__o41a_2
XFILLER_0_78_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput3 gpio_in[6] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_4
X_8861_ _4325_ _4337_ _4338_ _4297_ vssd1 vssd1 vccd1 vccd1 _4339_ sky130_fd_sc_hd__o22ai_1
X_7812_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[3\] _2975_ _3388_
+ _3390_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__a211o_1
X_8792_ _4260_ _4269_ vssd1 vssd1 vccd1 vccd1 _4270_ sky130_fd_sc_hd__nor2_1
XANTENNA__8713__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4960__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4955_ _0734_ _0735_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7743_ net105 net101 _3282_ vssd1 vssd1 vccd1 vccd1 _3333_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8148__B1 _3597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8432__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4886_ _0837_ _0838_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout140_A _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7674_ _3247_ _3263_ vssd1 vssd1 vccd1 vccd1 _3264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9413_ clknet_leaf_46_wb_clk_i _0401_ net233 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.drawDoneCactus
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__9317__Q team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6625_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[21\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[22\]
+ _2513_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[23\] vssd1
+ vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4959__Y _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9344_ clknet_leaf_47_wb_clk_i _0292_ net235 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6556_ _2467_ _2468_ _2469_ _2470_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__or4_1
X_5507_ _1216_ _1458_ _0856_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__a21bo_1
X_9275_ clknet_leaf_28_wb_clk_i _0274_ net241 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6487_ _2423_ _2424_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8226_ net121 _3730_ _3035_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5685__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5438_ _1339_ _1387_ _1388_ _1390_ net129 vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5369_ _1316_ _1318_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__a21oi_1
XANTENNA__6882__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8157_ net287 _0648_ vssd1 vssd1 vccd1 vccd1 _3677_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8088_ _3616_ vssd1 vssd1 vccd1 vccd1 _3617_ sky130_fd_sc_hd__inv_2
X_7108_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[5\]
+ _2842_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7039_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\] vssd1
+ vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_22_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8926__A2 _3200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9561__429 vssd1 vssd1 vccd1 vccd1 _9561__429/HI net429 sky130_fd_sc_hd__conb_1
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4870__B net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7665__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7702__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7421__B _3022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8533__A _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8917__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6053__A _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4740_ net280 _0693_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__or2_1
XANTENNA__6988__A team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4671_ _0614_ _0628_ _0613_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7390_ _2544_ _3002_ vssd1 vssd1 vccd1 vccd1 _3037_ sky130_fd_sc_hd__or2_1
X_6410_ _2360_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6341_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[5\] _2292_ vssd1
+ vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__or2_2
XFILLER_0_84_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6272_ _2110_ _2224_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__nand2_1
X_9060_ clknet_leaf_33_wb_clk_i _0195_ net245 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8853__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5223_ _1115_ _1120_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__and2_1
XANTENNA__4795__X _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6864__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8011_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] _3543_ vssd1
+ vssd1 vccd1 vccd1 _3548_ sky130_fd_sc_hd__nor2_1
X_5154_ _1089_ _1106_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5085_ _0820_ _0867_ _1001_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__a21o_2
XANTENNA_fanout188_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8913_ _4379_ _4383_ _4381_ _4380_ vssd1 vssd1 vccd1 vccd1 _4390_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4971__A _0809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8844_ _4312_ _4321_ _4318_ vssd1 vssd1 vccd1 vccd1 _4322_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5987_ _1887_ _1937_ _1938_ _1939_ vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8775_ _4244_ _4247_ _4252_ vssd1 vssd1 vccd1 vccd1 _4253_ sky130_fd_sc_hd__o21ai_1
X_4938_ net143 _0839_ _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout143_X net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7726_ net174 _3312_ vssd1 vssd1 vccd1 vccd1 _3316_ sky130_fd_sc_hd__nor2_1
X_4869_ _0762_ _0774_ _0821_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7657_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[6\]
+ _3240_ _3243_ vssd1 vssd1 vccd1 vccd1 _3247_ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6608_ _2505_ _2506_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[16\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7588_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[16\]
+ _2855_ _3177_ vssd1 vssd1 vccd1 vccd1 _3178_ sky130_fd_sc_hd__o21a_2
XFILLER_0_16_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9327_ clknet_leaf_29_wb_clk_i _0010_ net233 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6539_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[16\] _2457_
+ _2428_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9258_ clknet_leaf_19_wb_clk_i _0271_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.clk1
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5658__A1 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9189_ clknet_leaf_11_wb_clk_i _0039_ net219 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_8209_ net121 _3719_ _3036_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4865__B _0809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9283__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9212__RESET_B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8800__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7151__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6990__B team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5910_ _1836_ _1843_ _1844_ _1862_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__o31a_1
XANTENNA__4791__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6890_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ net270 _2692_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__and3b_1
XFILLER_0_75_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5841_ _0718_ _0909_ _1745_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5772_ _1659_ _1674_ _1673_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8560_ net169 _3618_ vssd1 vssd1 vccd1 vccd1 _4039_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4723_ _0676_ _0677_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__nand2_4
XFILLER_0_29_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7511_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\] _3032_
+ _3038_ _3023_ vssd1 vssd1 vccd1 vccd1 _3147_ sky130_fd_sc_hd__o211a_1
X_8491_ _3295_ _3299_ _3970_ _3311_ vssd1 vssd1 vccd1 vccd1 _3971_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7442_ _3084_ _3085_ _3049_ vssd1 vssd1 vccd1 vccd1 _3086_ sky130_fd_sc_hd__a21o_1
X_4654_ _0610_ _0611_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4585_ _0549_ _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7373_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\] _3021_
+ vssd1 vssd1 vccd1 vccd1 _3023_ sky130_fd_sc_hd__nand2_4
X_6324_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[0\] team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__nor2_1
X_9112_ clknet_leaf_46_wb_clk_i _0215_ net234 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout103_A _3276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6255_ _2121_ _2122_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__xnor2_1
X_9043_ clknet_leaf_35_wb_clk_i _0178_ net246 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6657__S _2532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5206_ _1142_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4966__A _0809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6186_ _1442_ _2138_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5137_ _1087_ _1088_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5068_ _0997_ _1020_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5797__A _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8173__A _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8827_ net317 net96 _4304_ vssd1 vssd1 vccd1 vccd1 _4305_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8758_ _3775_ _4212_ _0425_ vssd1 vssd1 vccd1 vccd1 _4236_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8762__B1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7709_ net153 net126 vssd1 vssd1 vccd1 vccd1 _3299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8689_ _4110_ _4143_ _4166_ _4167_ vssd1 vssd1 vccd1 vccd1 _4168_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7868__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5352__A_N _1011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9567__435 vssd1 vssd1 vccd1 vccd1 _9567__435/HI net435 sky130_fd_sc_hd__conb_1
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5500__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8811__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9574__439 vssd1 vssd1 vccd1 vccd1 _9574__439/HI net439 sky130_fd_sc_hd__conb_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[6\] vssd1
+ vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8520__A3 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold119 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.clk1
+ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8808__A1 _3976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6040_ _1951_ _1952_ vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_13_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7991_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[4\] _3527_ vssd1
+ vssd1 vccd1 vccd1 _3529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6942_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[6\]
+ _2403_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_6873_ _2680_ _2681_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5824_ _1775_ _1776_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_33_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8744__B1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_22_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8612_ _0674_ _3214_ vssd1 vssd1 vccd1 vccd1 _4091_ sky130_fd_sc_hd__xnor2_1
X_9592_ net456 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5755_ _1707_ _1706_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8543_ net152 _4018_ _4020_ vssd1 vssd1 vccd1 vccd1 _4022_ sky130_fd_sc_hd__o21ai_1
X_5686_ net131 _1592_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout318_A team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4706_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[2\] _0647_
+ _0659_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_20_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8474_ _3953_ vssd1 vssd1 vccd1 vccd1 _3954_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4637_ _0584_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__nand2b_2
X_7425_ _3068_ _3069_ net114 _3067_ vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__o211ai_4
XANTENNA__4533__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4568_ _0535_ _0536_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7356_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[4\] _3012_
+ _2974_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Left_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout106_X net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4499_ net16 net5 net30 net27 vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__or4_1
X_6307_ _2147_ _2181_ _2259_ _2180_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_90_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7287_ _2964_ vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__inv_2
XANTENNA__4696__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6238_ _2132_ _2134_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_90_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9026_ clknet_leaf_53_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[8\]
+ net200 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_6169_ _1954_ _1955_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_40_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8806__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7710__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5540_ _1491_ _1492_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5471_ _1420_ _1422_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6996__A team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7210_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[19\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[20\]
+ _2906_ net164 vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8190_ net279 _2387_ vssd1 vssd1 vccd1 vccd1 _3707_ sky130_fd_sc_hd__xor2_2
XFILLER_0_50_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7141_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[11\]
+ _2870_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__xor2_1
XANTENNA__5405__A _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7072_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[2\] vssd1
+ vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__nand2_1
X_6023_ _1841_ _1884_ _1883_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8435__B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7974_ net328 _2426_ _3507_ net297 _3512_ vssd1 vssd1 vccd1 vccd1 _3513_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout170_A _3472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5140__A _0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout268_A _2548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6925_ net530 _2714_ net267 vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9644_ net265 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6856_ net273 _2670_ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8193__A1 _3597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9575_ net440 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_5807_ _1710_ _1712_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__xnor2_1
X_6787_ net274 _2623_ _2624_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__nor3_1
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5738_ _1690_ _1689_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout223_X net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8526_ _0656_ net109 vssd1 vssd1 vccd1 vccd1 _4005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5669_ _1575_ _1621_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__nor2_1
X_8457_ _3330_ _3935_ _3936_ _3937_ vssd1 vssd1 vccd1 vccd1 _3938_ sky130_fd_sc_hd__or4b_1
XANTENNA__8496__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7408_ _3052_ _3048_ _3047_ vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__or3b_1
XFILLER_0_20_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8388_ net126 _3359_ vssd1 vssd1 vccd1 vccd1 _3869_ sky130_fd_sc_hd__nand2_2
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9056__RESET_B net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7514__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7339_ _2983_ _3004_ net121 vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9009_ clknet_leaf_6_wb_clk_i _0173_ net204 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5969__B _1912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5050__A _0999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8184__A1 _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload17 clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_11_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload28 clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_11_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload39 clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__inv_8
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7998__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6958__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4971_ _0809_ _0922_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4984__A1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6710_ net272 _2571_ _2572_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__nor3_1
X_7690_ _3265_ net98 vssd1 vssd1 vccd1 vccd1 _3280_ sky130_fd_sc_hd__nand2_4
XFILLER_0_58_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6641_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[27\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[28\]
+ _2523_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[29\] vssd1
+ vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9360_ clknet_leaf_26_wb_clk_i _0308_ net249 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8311_ net198 _3800_ _3540_ vssd1 vssd1 vccd1 vccd1 _3803_ sky130_fd_sc_hd__o21ai_1
X_6572_ _2482_ _2483_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[3\]
+ sky130_fd_sc_hd__nor2_1
X_5523_ _1450_ _1451_ _1475_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__nand3_1
X_9291_ clknet_leaf_14_wb_clk_i _0110_ net214 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5454_ _1358_ _1406_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__nand2_2
XFILLER_0_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8242_ _3034_ _3741_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5385_ _1287_ _1336_ _1335_ _1315_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__a211o_1
X_8173_ _0686_ _0707_ vssd1 vssd1 vccd1 vccd1 _3692_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4677__C _0634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout204 net206 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7124_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[15\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\] net184
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\] vssd1
+ vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__and4_2
Xfanout226 net228 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_4
Xfanout215 net216 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4974__A _0926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7055_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[0\]
+ _2789_ _2799_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[0\]
+ _2798_ vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__a221o_1
Xfanout248 net253 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
Xfanout259 net261 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_4
X_6006_ _0717_ _0931_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_31_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8938__B1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout173_X net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7957_ net330 net197 _3496_ net300 vssd1 vssd1 vccd1 vccd1 _3497_ sky130_fd_sc_hd__o211a_1
X_7888_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[17\]
+ _3439_ vssd1 vssd1 vccd1 vccd1 _3441_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6908_ _2704_ _2705_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8181__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9627_ net266 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6839_ net657 _2657_ net271 vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9558_ net426 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XANTENNA__9237__RESET_B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9489_ net364 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
X_8509_ net117 _3288_ _3883_ vssd1 vssd1 vccd1 vccd1 _3989_ sky130_fd_sc_hd__a21oi_2
XANTENNA__4868__B _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4884__A _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5170_ _0951_ _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nor2_1
XANTENNA__4794__A _0719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 wb_rst_i vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_1
XANTENNA__5402__B _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8860_ _4324_ _4336_ _4337_ vssd1 vssd1 vccd1 vccd1 _4338_ sky130_fd_sc_hd__or3_1
X_7811_ net597 _2974_ _3391_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__o21a_1
X_8791_ _0422_ _3486_ vssd1 vssd1 vccd1 vccd1 _4269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4954_ _0810_ _0905_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__nor2_4
XFILLER_0_47_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7742_ net95 net104 _3331_ _3330_ vssd1 vssd1 vccd1 vccd1 _3332_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_74_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4885_ _0835_ _0836_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__nor2_1
X_9412_ clknet_leaf_8_wb_clk_i _0400_ net223 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.drawDoneDino
+ sky130_fd_sc_hd__dfrtp_1
X_7673_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[4\]
+ _3254_ _3261_ vssd1 vssd1 vccd1 vccd1 _3263_ sky130_fd_sc_hd__and3_2
XFILLER_0_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6624_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[22\] _2514_
+ _2516_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[22\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout133_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9343_ clknet_leaf_47_wb_clk_i _0291_ net235 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6555_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[29\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[28\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[31\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[30\]
+ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__or4_1
XANTENNA__9330__RESET_B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5506_ _1215_ _1458_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__and2b_1
X_9274_ clknet_leaf_20_wb_clk_i _0273_ net239 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr1\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_15_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6486_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[6\] team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ net294 vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__mux2_1
XANTENNA__6331__A0 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8225_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[13\]
+ _2991_ vssd1 vssd1 vccd1 vccd1 _3730_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_5_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5437_ _1387_ _1389_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__xnor2_2
X_5368_ _1271_ _1320_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8156_ _3597_ _3675_ _3676_ net243 net591 vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__o32a_1
X_5299_ _1039_ _1047_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8087_ net178 _0706_ vssd1 vssd1 vccd1 vccd1 _3616_ sky130_fd_sc_hd__nand2b_1
X_7107_ _2842_ _2843_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7038_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[2\] _2777_
+ _2785_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_52_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8989_ clknet_leaf_7_wb_clk_i _0153_ net205 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7079__X _2823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9071__RESET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5046__Y _0999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7702__B net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6053__B _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6988__B team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7889__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4670_ _0617_ _0627_ _0616_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6340_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[4\] team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[3\]
+ _2291_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6271_ _2108_ _2109_ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5222_ _1169_ _1174_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nor2_1
X_8010_ _3538_ _3539_ _3546_ vssd1 vssd1 vccd1 vccd1 _3547_ sky130_fd_sc_hd__a21oi_2
X_5153_ _0866_ _1105_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__nor2_1
XANTENNA__8066__A0 _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7612__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8708__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5413__A _1217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5084_ _0748_ _0971_ _1017_ _1019_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__a31o_1
X_8912_ _4385_ _4388_ vssd1 vssd1 vccd1 vccd1 _4389_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4971__B _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8369__B2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8843_ net320 _4302_ _4320_ vssd1 vssd1 vccd1 vccd1 _4321_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5986_ _1843_ _1886_ _1885_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__a21o_1
X_8774_ net103 _4243_ vssd1 vssd1 vccd1 vccd1 _4252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4937_ _0747_ _0769_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9328__Q team_08_WB.instance_to_wrap.allocation.game.controller.state\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7725_ _3307_ _3314_ vssd1 vssd1 vccd1 vccd1 _3315_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_96_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4868_ _0762_ _0773_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7656_ _3237_ _3244_ vssd1 vssd1 vccd1 vccd1 _3246_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout136_X net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6607_ net654 _2503_ _2478_ vssd1 vssd1 vccd1 vccd1 _2506_ sky130_fd_sc_hd__o21ai_1
XANTENNA__8541__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8541__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4799_ _0593_ _0595_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__xnor2_4
X_9326_ clknet_leaf_30_wb_clk_i _0009_ net237 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7587_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[16\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[15\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\] vssd1
+ vssd1 vccd1 vccd1 _3177_ sky130_fd_sc_hd__nand4_4
XFILLER_0_63_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6538_ _2457_ _2458_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[15\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9257_ clknet_leaf_15_wb_clk_i _0095_ net214 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_6469_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[19\]
+ _2405_ _2411_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[22\]
+ vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9188_ clknet_leaf_11_wb_clk_i _0038_ net220 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8208_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[7\]
+ _2987_ vssd1 vssd1 vccd1 vccd1 _3719_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8057__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8139_ net299 _3454_ vssd1 vssd1 vccd1 vccd1 _3664_ sky130_fd_sc_hd__nor2_1
XANTENNA__8618__B net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8634__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6791__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7638__A3 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4857__B1 _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8048__B1 _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8599__B2 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4791__B _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5840_ net167 _0905_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9624__482 vssd1 vssd1 vccd1 vccd1 _9624__482/HI net482 sky130_fd_sc_hd__conb_1
X_5771_ _1722_ _1723_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4722_ net284 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7510_ net518 _3146_ net115 vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8490_ net112 net108 _3864_ _3969_ vssd1 vssd1 vccd1 vccd1 _3970_ sky130_fd_sc_hd__a31o_1
XFILLER_0_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7441_ net310 _0442_ _3045_ net306 _3051_ vssd1 vssd1 vccd1 vccd1 _3085_ sky130_fd_sc_hd__o221a_1
Xinput40 wbs_we_i vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
XFILLER_0_86_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4653_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[5\] vssd1
+ vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__nand2b_1
XANTENNA__8602__A1_N net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4584_ net334 team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] vssd1
+ vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__nand2b_2
X_7372_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[2\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8287__B1 _3511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6323_ _2273_ _2274_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__or2_1
XANTENNA__8719__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9111_ clknet_leaf_46_wb_clk_i _0214_ net234 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[2\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7629__A3 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6254_ _0445_ _2206_ vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__nor2_1
X_9042_ clknet_leaf_35_wb_clk_i _0177_ net246 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5205_ _0863_ _1103_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6185_ _1495_ _2137_ _1493_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout298_A team_08_WB.instance_to_wrap.allocation.game.controller.state\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5136_ _1087_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5067_ _1008_ _1018_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout253_X net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8826_ net320 net101 vssd1 vssd1 vccd1 vccd1 _4304_ sky130_fd_sc_hd__nand2_1
X_5969_ _1910_ _1912_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__xnor2_1
X_8757_ _0520_ _4232_ vssd1 vssd1 vccd1 vccd1 _4235_ sky130_fd_sc_hd__nand2_1
XANTENNA__6702__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7708_ _3286_ _3287_ _3289_ _3293_ _3297_ vssd1 vssd1 vccd1 vccd1 _3298_ sky130_fd_sc_hd__a41o_1
XFILLER_0_35_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8688_ net107 _4113_ vssd1 vssd1 vccd1 vccd1 _4167_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_90_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7639_ _3204_ _3228_ vssd1 vssd1 vccd1 vccd1 _3229_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_95_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9309_ clknet_leaf_1_wb_clk_i _0280_ net207 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.game.score\[3\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_101_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input26_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7005__A1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8811__B net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5319__A1 _1038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold109 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[1\]
+ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7990_ net289 _3527_ vssd1 vssd1 vccd1 vccd1 _3528_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6941_ net604 _2404_ _2723_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6872_ net688 _2679_ net269 vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9591_ net455 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
X_5823_ _1728_ _1730_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__xor2_1
XANTENNA__6755__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8611_ _0703_ _3610_ vssd1 vssd1 vccd1 vccd1 _4090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8542_ net177 _4019_ vssd1 vssd1 vccd1 vccd1 _4021_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5754_ _1655_ _1656_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__xor2_1
X_5685_ net131 _1637_ _1636_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4705_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[2\] _0647_
+ _0659_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_20_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8473_ net117 _3301_ _3883_ vssd1 vssd1 vccd1 vccd1 _3953_ sky130_fd_sc_hd__a21o_1
X_4636_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[3\] vssd1
+ vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_44_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7424_ net312 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_floor team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_cactus
+ _3021_ vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__or4_2
XANTENNA__4533__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7355_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[2\] _2974_
+ _3012_ _3013_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__o22a_1
XANTENNA__7624__Y _3214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6306_ _2144_ _2184_ _2258_ _2182_ _2183_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4567_ _0504_ _0505_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4498_ net32 net31 net34 net33 vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__or4_1
X_7286_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[20\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[19\]
+ _2960_ vssd1 vssd1 vccd1 vccd1 _2964_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6237_ _1551_ _2135_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_90_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9025_ clknet_leaf_53_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[7\]
+ net200 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6168_ _1995_ _2120_ _1994_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5119_ _0817_ _1071_ _1035_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6099_ net142 _0916_ _1974_ _1973_ vssd1 vssd1 vccd1 vccd1 _2052_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8471__X _3952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8809_ _4219_ _4229_ _4230_ vssd1 vssd1 vccd1 vccd1 _4287_ sky130_fd_sc_hd__or3b_1
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8631__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6432__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5048__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5990__B _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4887__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8816__A_N net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8806__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7710__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8094__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7777__A2 _3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9580__444 vssd1 vssd1 vccd1 vccd1 _9580__444/HI net444 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_86_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5470_ _1422_ _1420_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6996__B team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5712__A1 _0809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4797__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7140_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[10\]
+ _2848_ _2850_ _2868_ vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__a22o_1
X_7071_ _2813_ _2816_ _2779_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__o21a_1
XFILLER_0_10_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5476__B1 _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9515__390 vssd1 vssd1 vccd1 vccd1 _9515__390/HI net390 sky130_fd_sc_hd__conb_1
X_6022_ _1958_ _1974_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__xnor2_1
XANTENNA__9355__RESET_B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7973_ net327 net197 _3510_ _3511_ vssd1 vssd1 vccd1 vccd1 _3512_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6924_ _2714_ _2715_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout163_A _0684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9643_ net265 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6855_ _0466_ _2668_ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9574_ net439 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_92_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5806_ _1757_ _1758_ _1756_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__a21o_1
X_6786_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[8\]
+ _2620_ vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout330_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5737_ net131 _1637_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8525_ _4002_ _4003_ vssd1 vssd1 vccd1 vccd1 _4004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8456_ net172 _3884_ _3888_ _3889_ vssd1 vssd1 vccd1 vccd1 _3937_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_92_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5668_ _0747_ _1574_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4978__Y _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7407_ net304 _3050_ _3049_ vssd1 vssd1 vccd1 vccd1 _3052_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8496__A3 _3864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5599_ net143 _1501_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__or2_1
X_4619_ _0575_ _0576_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_5_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8387_ net124 _3360_ vssd1 vssd1 vccd1 vccd1 _3868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7338_ net542 _2982_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7269_ net573 _2950_ _2952_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__a21oi_1
X_9008_ clknet_leaf_6_wb_clk_i _0172_ net204 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__9096__RESET_B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6427__A _2368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9605__469 vssd1 vssd1 vccd1 vccd1 _9605__469/HI net469 sky130_fd_sc_hd__conb_1
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload18 clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinv_8
Xclkload29 clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_11_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7695__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__7424__C team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_cactus vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9437__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7998__A2 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4970_ _0810_ _0921_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4984__A2 _0926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6640_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[28\] _2524_
+ _2526_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[28\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6571_ net676 _2481_ net263 vssd1 vssd1 vccd1 vccd1 _2483_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5522_ _0940_ _1419_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__xnor2_1
X_8310_ team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[4\] _3776_ net322
+ vssd1 vssd1 vccd1 vccd1 _3802_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9290_ clknet_leaf_14_wb_clk_i _0109_ net213 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5453_ _1014_ _1357_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__or2_1
X_8241_ _2998_ _3740_ net122 vssd1 vssd1 vccd1 vccd1 _3741_ sky130_fd_sc_hd__a21o_1
X_5384_ _1315_ _1335_ _1336_ _1287_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__o211ai_2
X_8172_ _2394_ _3689_ _3690_ _3688_ _0654_ vssd1 vssd1 vccd1 vccd1 _3691_ sky130_fd_sc_hd__o32a_1
Xfanout205 net206 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_2
XFILLER_0_1_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7123_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[15\]
+ _2852_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__or2_1
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_4
Xfanout216 net232 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_2
Xfanout238 net254 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
XANTENNA__8727__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout249 net251 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
X_7054_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\]
+ _2788_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[8\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[3\] vssd1
+ vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__and4bb_1
X_6005_ net142 _0916_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5621__B1 _1088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout166_X net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7956_ net197 _3495_ vssd1 vssd1 vccd1 vccd1 _3496_ sky130_fd_sc_hd__nand2_1
X_7887_ _3439_ _3440_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[16\]
+ net166 vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__a2bb2o_1
X_6907_ net662 _2702_ net267 vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8166__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9626_ net266 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
X_6838_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[12\]
+ _2657_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9557_ net425 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6769_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__nand3_1
XFILLER_0_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8508_ _3898_ _3987_ _3327_ vssd1 vssd1 vccd1 vccd1 _3988_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9488_ net363 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_66_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6710__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8439_ net151 _3324_ _3334_ net94 vssd1 vssd1 vccd1 vccd1 _3920_ sky130_fd_sc_hd__nand4_1
XFILLER_0_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9570__498 vssd1 vssd1 vccd1 vccd1 net498 _9570__498/LO sky130_fd_sc_hd__conb_1
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5061__A _1012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8372__A team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7716__A _3305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4794__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_1
X_9586__450 vssd1 vssd1 vccd1 vccd1 _9586__450/HI net450 sky130_fd_sc_hd__conb_1
X_7810_ _3387_ _3390_ vssd1 vssd1 vccd1 vccd1 _3391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8790_ net324 _4260_ vssd1 vssd1 vccd1 vccd1 _4268_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8282__A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4953_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7741_ net191 net188 net185 vssd1 vssd1 vccd1 vccd1 _3331_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7672_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[4\]
+ _3261_ vssd1 vssd1 vccd1 vccd1 _3262_ sky130_fd_sc_hd__nand2_1
X_4884_ _0835_ _0836_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__and2_2
XFILLER_0_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9411_ clknet_leaf_46_wb_clk_i _0358_ net233 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.cactusMovement
+ sky130_fd_sc_hd__dfrtp_1
X_6623_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[22\] _2514_
+ net255 vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9342_ clknet_leaf_4_wb_clk_i net558 net205 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.det
+ sky130_fd_sc_hd__dfrtp_1
X_6554_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[25\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[24\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[27\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[26\]
+ vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout126_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5505_ _0811_ _0909_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9273_ clknet_leaf_28_wb_clk_i _0272_ net241 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr1\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_6485_ _0431_ _0700_ vssd1 vssd1 vccd1 vccd1 _2423_ sky130_fd_sc_hd__nor2_1
X_5436_ _1339_ _1388_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__nand2_1
XANTENNA__5146__A _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8224_ _3727_ _3729_ _3711_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9370__RESET_B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5367_ _1220_ _1270_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__or2_1
XANTENNA__7361__A _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8155_ _0689_ net137 _3674_ net139 vssd1 vssd1 vccd1 vccd1 _3676_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_11_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5298_ _1202_ _1250_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8086_ _0657_ _0660_ net183 _2286_ vssd1 vssd1 vccd1 vccd1 _3615_ sky130_fd_sc_hd__a31o_1
X_7106_ net185 _0557_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_87_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7037_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[1\] vssd1
+ vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_52_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8904__B _3178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8988_ net4 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7939_ _0654_ net137 vssd1 vssd1 vccd1 vccd1 _3479_ sky130_fd_sc_hd__nand2_2
XFILLER_0_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9609_ net473 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_80_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4879__B _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4895__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8367__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7586__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6010__B1 _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8087__A_N net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9434__Q team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6270_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[5\]
+ _2222_ vssd1 vssd1 vccd1 vccd1 _2223_ sky130_fd_sc_hd__and2_1
X_5221_ _1172_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__nand2_1
XANTENNA__8277__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7181__A _2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5152_ _0862_ _0865_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8066__A1 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5083_ _1024_ _1025_ _1021_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8911_ _0689_ net118 _4029_ _4386_ _4387_ vssd1 vssd1 vccd1 vccd1 _4388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8842_ _0423_ net320 net105 net103 vssd1 vssd1 vccd1 vccd1 _4320_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8773_ _4244_ _4250_ _4247_ _4241_ vssd1 vssd1 vccd1 vccd1 _4251_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5985_ _1935_ _1936_ _1923_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__a21o_1
X_7724_ net126 net120 vssd1 vssd1 vccd1 vccd1 _3314_ sky130_fd_sc_hd__or2_2
X_4936_ _0882_ _0888_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout243_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4867_ _0813_ _0819_ _0816_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7655_ _3237_ _3244_ vssd1 vssd1 vccd1 vccd1 _3245_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_31_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6606_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[15\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[16\]
+ _2502_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7586_ net290 team_08_WB.instance_to_wrap.allocation.game.game.score\[6\] net259
+ _2344_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout129_X net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4798_ _0750_ net144 _0741_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__or3b_2
X_9325_ clknet_leaf_29_wb_clk_i _0008_ net237 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4699__B _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6537_ net660 _2455_ _2429_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4986__Y _0939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9256_ clknet_leaf_15_wb_clk_i _0094_ net213 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_6468_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[16\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[15\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[14\]
+ _2410_ _2406_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__a41o_1
XFILLER_0_101_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5419_ _1364_ _1369_ _1371_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__a21o_1
X_9187_ clknet_leaf_11_wb_clk_i _0037_ net220 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_8207_ _3029_ _3033_ _3718_ _3002_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6399_ _2335_ _2340_ _2349_ _2347_ _2346_ vssd1 vssd1 vccd1 vccd1 _2350_ sky130_fd_sc_hd__a32oi_4
XANTENNA__5604__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8057__A1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8138_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[8\]
+ net243 _3656_ _3663_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input3_X net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8069_ _3597_ _3599_ _3600_ net243 net560 vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__o32a_1
XANTENNA__8634__B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4507__X _0478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7568__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6345__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5770_ _1706_ _1707_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4721_ net284 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6080__A _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4652_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[5\] vssd1
+ vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7176__A _2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7440_ net306 _3045_ vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput30 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4583_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] net334 vssd1
+ vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__nand2b_1
X_9110_ clknet_leaf_29_wb_clk_i _0213_ net233 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7371_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[2\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8287__A1 _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6322_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[3\] _2265_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__a21oi_1
X_9551__419 vssd1 vssd1 vccd1 vccd1 _9551__419/HI net419 sky130_fd_sc_hd__conb_1
X_6253_ _1921_ _2123_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9041_ clknet_leaf_34_wb_clk_i _0176_ net246 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5204_ _0862_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__nand2_1
X_6184_ _1551_ _2135_ _1548_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__a21bo_1
XANTENNA__5143__B _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5135_ _0769_ _0785_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__xor2_4
XANTENNA_fanout193_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8735__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5066_ _1008_ _1018_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9339__Q team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8825_ _4300_ _4301_ _4302_ vssd1 vssd1 vccd1 vccd1 _4303_ sky130_fd_sc_hd__o21ba_1
X_5968_ _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8756_ net317 _3542_ vssd1 vssd1 vccd1 vccd1 _4234_ sky130_fd_sc_hd__nand2_1
X_4919_ _0858_ _0866_ _0870_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__nor3_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7707_ _3290_ _3296_ net172 vssd1 vssd1 vccd1 vccd1 _3297_ sky130_fd_sc_hd__o21a_1
X_5899_ _1803_ _1850_ _1851_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8687_ _4111_ _4112_ _4145_ vssd1 vssd1 vccd1 vccd1 _4166_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7638_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[8\]
+ _3217_ net117 _3216_ vssd1 vssd1 vccd1 vccd1 _3228_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7569_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr1\[0\] net541 _3170_
+ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9320__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9308_ clknet_leaf_1_wb_clk_i _0279_ net208 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.game.score\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_9239_ clknet_leaf_19_wb_clk_i _0266_ net239 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr1\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9491__366 vssd1 vssd1 vccd1 vccd1 _9491__366/HI net366 sky130_fd_sc_hd__conb_1
XFILLER_0_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7025__S net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8645__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8450__A1 _3916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8380__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5509__A _0814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8505__A2 _3976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7724__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6940_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[7\]
+ _2404_ net157 vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__o21ai_1
XANTENNA__8274__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6871_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[9\]
+ _2679_ vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__and2_1
XANTENNA__9159__Q team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9590_ net454 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
X_5822_ _1773_ _1774_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8610_ net102 _3280_ _4088_ vssd1 vssd1 vccd1 vccd1 _4089_ sky130_fd_sc_hd__or3b_1
X_5753_ _1012_ _1694_ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_57_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8541_ net152 _4018_ _4019_ net177 vssd1 vssd1 vccd1 vccd1 _4020_ sky130_fd_sc_hd__a22oi_1
X_4704_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\] vssd1 vssd1 vccd1
+ vccd1 _0659_ sky130_fd_sc_hd__a21oi_2
X_5684_ _1633_ _1635_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8472_ net208 _2396_ _3952_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4635_ _0586_ _0592_ _0585_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__a21o_2
XFILLER_0_44_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7423_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_dino _3064_ vssd1
+ vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_25_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout206_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4566_ _0523_ _0534_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__nand2_1
X_7354_ _3009_ _3010_ _2975_ vssd1 vssd1 vccd1 vccd1 _3013_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6305_ _2139_ _2188_ _2257_ _2185_ _2187_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8449__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7285_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[19\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[18\]
+ _2958_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[20\]
+ vssd1 vssd1 vccd1 vccd1 _2963_ sky130_fd_sc_hd__a31o_1
X_9024_ clknet_leaf_53_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[6\]
+ net201 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4497_ net312 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__inv_2
X_6236_ _1494_ _2137_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_90_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6167_ _2032_ _2119_ _2031_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5118_ _1029_ _1066_ _1070_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6098_ _2024_ _2050_ _2049_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__or3b_1
X_5049_ net138 _1000_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_49_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7809__A _2972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8808_ _3976_ _4280_ _4282_ _4285_ _4259_ vssd1 vssd1 vccd1 vccd1 _4286_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_45_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8739_ net332 net191 vssd1 vssd1 vccd1 vccd1 _4217_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5239__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5712__A2 _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4797__B net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7070_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[2\]
+ _2799_ _2810_ _2815_ vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6021_ _1971_ _1972_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6425__B1 _2325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7972_ _0463_ _3472_ vssd1 vssd1 vccd1 vccd1 _3511_ sky130_fd_sc_hd__nor2_2
X_6923_ net642 _2713_ net267 vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__o21ai_1
X_9642_ net264 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6854_ net269 _2665_ _2668_ _2669_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9573_ net438 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5805_ _1709_ _1755_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6785_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[7\]
+ _2620_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__a21oi_1
X_5736_ net131 _1688_ _1687_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8524_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\] net106
+ vssd1 vssd1 vccd1 vccd1 _4003_ sky130_fd_sc_hd__and2_1
X_5667_ _1619_ net143 vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__and2b_1
X_9557__425 vssd1 vssd1 vccd1 vccd1 _9557__425/HI net425 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_40_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8455_ _3302_ net94 _3359_ net171 vssd1 vssd1 vccd1 vccd1 _3936_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_92_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4618_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[6\] vssd1
+ vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7406_ net307 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout111_X net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8496__A4 _3888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5598_ _1550_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout209_X net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8386_ net154 _3862_ _3866_ _3863_ vssd1 vssd1 vccd1 vccd1 _3867_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4549_ net333 net324 net313 net334 vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__or4b_1
X_7337_ _2982_ _3003_ net121 vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7268_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[14\]
+ _2950_ net180 vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5467__A1 _0939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6219_ _2170_ _2171_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__xnor2_1
X_9007_ clknet_leaf_5_wb_clk_i _0171_ net205 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7199_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[15\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[16\]
+ _2900_ vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9065__RESET_B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5059__A _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload19 clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload19/X sky130_fd_sc_hd__clkbuf_4
X_9497__372 vssd1 vssd1 vccd1 vccd1 _9497__372/HI net372 sky130_fd_sc_hd__conb_1
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8089__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8817__B net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5522__A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9437__Q team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6570_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[3\] _2481_ vssd1
+ vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__and2_1
X_5521_ _0939_ _1473_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8240_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[19\]
+ _2996_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[20\]
+ vssd1 vssd1 vccd1 vccd1 _3740_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5452_ _0748_ _1404_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7615__C net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5383_ _1269_ _1286_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8171_ net287 _2388_ net285 vssd1 vssd1 vccd1 vccd1 _3690_ sky130_fd_sc_hd__a21oi_1
XANTENNA__7912__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8096__C1 _3597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7122_ net184 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\]
+ _2851_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__and3_1
Xfanout228 net231 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
Xfanout217 net221 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_4
X_7053_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\]
+ _2781_ _2787_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2801_ sky130_fd_sc_hd__nor4b_1
Xfanout206 net232 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
X_6004_ _1942_ _1945_ _1944_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__a21o_1
Xfanout239 net242 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout273_A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5621__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7955_ _3493_ _3494_ vssd1 vssd1 vccd1 vccd1 _3495_ sky130_fd_sc_hd__nand2_1
X_7886_ _0448_ _3438_ net160 vssd1 vssd1 vccd1 vccd1 _3440_ sky130_fd_sc_hd__a21bo_1
X_6906_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[6\]
+ _2700_ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9625_ net265 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
X_6837_ net275 _2656_ _2657_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__nor3_1
XANTENNA__8020__C1 _3556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9556_ net424 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_9_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6768_ net586 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ _2612_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_8507_ _3293_ _3959_ _3297_ vssd1 vssd1 vccd1 vccd1 _3987_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_28_Left_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5719_ _0934_ _1671_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__nor2_1
X_6699_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[7\]
+ _2563_ _2565_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__o21a_1
X_9487_ net362 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_66_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8874__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7677__A2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8438_ _3908_ _3918_ vssd1 vssd1 vccd1 vccd1 _3919_ sky130_fd_sc_hd__nor2_1
X_8369_ _3853_ _3843_ _2875_ net289 vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__7822__A team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9531__406 vssd1 vssd1 vccd1 vccd1 _9531__406/HI net406 sky130_fd_sc_hd__conb_1
XANTENNA__6637__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8637__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9246__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5612__A1 _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8372__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4899__Y _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8865__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7732__A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4794__C _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_1
XFILLER_0_87_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4952_ _0734_ _0904_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__nand2_4
XFILLER_0_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7740_ _3280_ _3329_ vssd1 vssd1 vccd1 vccd1 _3330_ sky130_fd_sc_hd__and2_2
XFILLER_0_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4883_ _0751_ _0756_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7671_ _3259_ _3260_ vssd1 vssd1 vccd1 vccd1 _3261_ sky130_fd_sc_hd__or2_4
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9410_ clknet_leaf_31_wb_clk_i _0357_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_6622_ _2514_ _2515_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[21\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__8305__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9341_ clknet_leaf_3_wb_clk_i net499 net202 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.button
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6553_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[19\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[18\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[17\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[16\]
+ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__or4bb_1
XANTENNA__7626__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5504_ _1217_ _1412_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__xor2_1
X_9272_ clknet_leaf_10_wb_clk_i _0081_ net228 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_6484_ net294 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoMovement net590
+ _2422_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a31o_1
X_5435_ _1337_ _1338_ _1327_ _1330_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8223_ _2991_ _3728_ net122 vssd1 vssd1 vccd1 vccd1 _3729_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout119_A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5366_ _1316_ _1318_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__nand2_1
XANTENNA__7361__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8154_ _0654_ _2537_ _3608_ _2393_ vssd1 vssd1 vccd1 vccd1 _3675_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_10_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5297_ _1048_ _1201_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__nand2_1
X_8085_ _0656_ _0661_ _0689_ _2285_ vssd1 vssd1 vccd1 vccd1 _3614_ sky130_fd_sc_hd__or4_2
XFILLER_0_10_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7105_ net185 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[4\]
+ _0557_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_87_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7036_ net3 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.tft_sdi
+ _2779_ _2784_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8987_ net312 vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7938_ _3473_ _3474_ _3478_ net225 net607 vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__o32a_1
XFILLER_0_33_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9608_ net472 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_77_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7869_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[11\] _3424_
+ vssd1 vssd1 vccd1 vccd1 _3428_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9539_ net495 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_80_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5056__B _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6858__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4895__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7035__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8383__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7586__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6010__A1 _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6010__B2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5220_ _0943_ _1171_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5151_ _0862_ _1102_ _1101_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5082_ _0953_ _0956_ _1033_ _1034_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7813__A2 _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8910_ _0689_ net118 net111 _0663_ vssd1 vssd1 vccd1 vccd1 _4387_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8841_ _4312_ _4315_ _4316_ _4318_ vssd1 vssd1 vccd1 vccd1 _4319_ sky130_fd_sc_hd__or4b_1
XFILLER_0_17_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8772_ _4240_ _4248_ _4249_ vssd1 vssd1 vccd1 vccd1 _4250_ sky130_fd_sc_hd__or3_1
X_5984_ _1923_ _1935_ _1936_ vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__nand3_1
X_7723_ _3241_ _3286_ net112 vssd1 vssd1 vccd1 vccd1 _3313_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4935_ _0837_ _0887_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__xor2_1
X_4866_ net144 _0813_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout236_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7654_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[6\]
+ _3238_ net108 vssd1 vssd1 vccd1 vccd1 _3244_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4797_ _0718_ net168 vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6605_ net683 _2502_ _2504_ _2478_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[15\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7585_ net290 team_08_WB.instance_to_wrap.allocation.game.game.score\[5\] net259
+ _2350_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9324_ clknet_leaf_29_wb_clk_i _0007_ net233 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8829__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6536_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[14\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[15\]
+ _2453_ vssd1 vssd1 vccd1 vccd1 _2457_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4996__A _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9255_ clknet_leaf_15_wb_clk_i _0093_ net215 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_6467_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[9\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[8\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[7\]
+ _2409_ vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5418_ _1318_ _1370_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__nand2_1
X_9186_ clknet_leaf_11_wb_clk_i _0036_ net218 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_8206_ _2987_ _3717_ vssd1 vssd1 vccd1 vccd1 _3718_ sky130_fd_sc_hd__nand2_1
X_6398_ team_08_WB.instance_to_wrap.allocation.game.game.score\[5\] _2339_ vssd1 vssd1
+ vccd1 vccd1 _2349_ sky130_fd_sc_hd__nand2_1
X_5349_ _1300_ _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__and2b_1
XANTENNA__5604__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8057__A2 _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8137_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\] _3653_ _3654_
+ _3662_ vssd1 vssd1 vccd1 vccd1 _3663_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8068_ _0656_ _0702_ _2419_ _3596_ vssd1 vssd1 vccd1 vccd1 _3600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5620__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7019_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\] _2773_
+ _0459_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6451__A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5801__Y _1754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6185__X _2138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6361__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4720_ _0669_ net178 vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__nand2_2
XFILLER_0_86_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4651_ _0607_ _0608_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__nand2b_1
XANTENNA__9445__Q team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput20 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7370_ team_08_WB.instance_to_wrap.allocation.game.controller.color\[11\] net238
+ _3018_ _3020_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__o22a_1
X_4582_ _0419_ _0548_ _0420_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[2\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6321_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[3\] team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[4\]
+ _2265_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6252_ _0446_ _2204_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9040_ clknet_leaf_34_wb_clk_i _0175_ net246 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6183_ _1551_ _2135_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__nand2_1
X_5203_ _1152_ _1154_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__xnor2_1
X_5134_ _0824_ _0839_ _0837_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__a21o_2
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7920__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5065_ _0972_ _1017_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout186_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_2__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8824_ net324 net104 vssd1 vssd1 vccd1 vccd1 _4302_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5967_ _1919_ _1918_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8755_ _3542_ _3763_ vssd1 vssd1 vccd1 vccd1 _4233_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4918_ _0858_ _0866_ _0870_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout141_X net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8686_ net125 _3622_ _4157_ _4164_ vssd1 vssd1 vccd1 vccd1 _4165_ sky130_fd_sc_hd__o211a_1
X_7706_ net124 net117 vssd1 vssd1 vccd1 vccd1 _3296_ sky130_fd_sc_hd__nor2_1
X_5898_ net142 _0927_ _1801_ _1802_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7637_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[8\]
+ net117 vssd1 vssd1 vccd1 vccd1 _3227_ sky130_fd_sc_hd__xor2_2
XFILLER_0_90_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4849_ _0794_ _0801_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__xor2_2
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7568_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr1\[0\] _3169_ net257
+ vssd1 vssd1 vccd1 vccd1 _3170_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7373__Y _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6519_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[9\] _2443_
+ _2429_ vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__o21ai_1
X_7499_ net522 net114 _3121_ _3137_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__o22a_1
X_9307_ clknet_leaf_1_wb_clk_i _0278_ net211 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.game.score\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9238_ clknet_leaf_18_wb_clk_i _0053_ net240 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout99_A _3266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9169_ _0144_ _0406_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8645__B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6213__A1 _1038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5509__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9239__SET_B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4527__A1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8910__B1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9442__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7724__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5244__B _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7740__A _3280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6204__A1 _1047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6870_ net273 _2678_ _2679_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__nor3_1
XFILLER_0_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5821_ _0749_ _1139_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_33_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5752_ _1704_ _1703_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_60_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4604__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7187__A _2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8540_ _0696_ _4016_ vssd1 vssd1 vccd1 vccd1 _4019_ sky130_fd_sc_hd__xor2_1
XFILLER_0_72_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4703_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\] _0656_ vssd1
+ vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__nand2_2
X_5683_ _1633_ _1635_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8471_ _3942_ _3951_ _3950_ vssd1 vssd1 vccd1 vccd1 _3952_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4634_ _0589_ _0591_ _0588_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7422_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_floor _3065_ _3066_
+ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__or3_2
X_4565_ _0526_ _0529_ _0531_ _0533_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__and4_1
X_7353_ _3009_ _3010_ vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6304_ _2136_ _2190_ _2192_ _2256_ _2189_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout101_A _3277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4496_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1 vssd1 vccd1
+ vccd1 _0468_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7284_ net584 _2960_ _2962_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9023_ clknet_leaf_53_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[5\]
+ net200 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_6235_ _1442_ _2138_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_90_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _2058_ _2118_ _2057_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5117_ _1027_ _1030_ _1067_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__o211a_1
X_6097_ _1982_ _2023_ _2022_ vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__a21oi_1
X_5048_ net138 _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8481__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8807_ _4264_ _4284_ _4278_ vssd1 vssd1 vccd1 vccd1 _4285_ sky130_fd_sc_hd__a21o_1
X_6999_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] _0467_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] vssd1 vssd1 vccd1 vccd1
+ _2762_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8738_ net332 net191 vssd1 vssd1 vccd1 vccd1 _4216_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_97_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8669_ _4109_ _4146_ _4147_ vssd1 vssd1 vccd1 vccd1 _4148_ sky130_fd_sc_hd__or3_1
XFILLER_0_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5345__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input31_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8959__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5239__B _1144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6370__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8566__A _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6020_ _1972_ _1971_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6086__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6425__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7971_ _3503_ _3509_ vssd1 vssd1 vccd1 vccd1 _3510_ sky130_fd_sc_hd__nand2_1
X_6922_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[12\]
+ _2713_ vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__and2_1
XANTENNA__8178__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9641_ net266 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6853_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5804_ _0791_ _0926_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9572_ net437 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6784_ net678 _2620_ _2622_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout149_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5735_ _1685_ _1686_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8523_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\] net106
+ vssd1 vssd1 vccd1 vccd1 _4002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5666_ net147 _0859_ _1141_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_40_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8454_ net104 _3331_ net95 vssd1 vssd1 vccd1 vccd1 _3935_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_92_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4617_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[6\] vssd1
+ vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7405_ _0439_ _0442_ vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__nor2_1
X_5597_ _1548_ _1549_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__nand2_1
XANTENNA__5165__A _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8385_ _3865_ vssd1 vssd1 vccd1 vccd1 _3866_ sky130_fd_sc_hd__inv_2
X_4548_ _0513_ _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__nand2_1
X_7336_ net539 net501 vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout104_X net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4479_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[1\] vssd1 vssd1
+ vccd1 vccd1 _0451_ sky130_fd_sc_hd__inv_2
X_7267_ net179 _2949_ _2951_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__and3_1
XANTENNA__7651__Y _3241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6218_ _1037_ _1060_ _1063_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__a21boi_1
X_9006_ clknet_leaf_5_wb_clk_i _0170_ net205 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__7380__A team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7198_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[15\] _2900_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[16\]
+ vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__a21oi_1
X_6149_ _2100_ _2101_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9034__RESET_B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7695__A3 _3284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5803__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4984__A4 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5520_ _1470_ _1471_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5451_ _1402_ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5382_ _1332_ _1334_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__nor2_1
X_8170_ net287 net284 _2388_ vssd1 vssd1 vccd1 vccd1 _3689_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6809__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7121_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[12\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\]
+ _2851_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__and4_1
XANTENNA__5713__A _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout229 net230 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
Xfanout218 net221 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
X_7052_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\]
+ _2780_ _2781_ vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__nor3_4
Xfanout207 net210 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_4
X_6003_ _1955_ _1954_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7954_ _0494_ _3491_ vssd1 vssd1 vccd1 vccd1 _3494_ sky130_fd_sc_hd__nand2b_1
XANTENNA__5621__A2 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6905_ _2702_ _2703_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7885_ _0448_ _3438_ vssd1 vssd1 vccd1 vccd1 _3439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9624_ net482 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
X_6836_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[10\]
+ _2653_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8020__B1 _3472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8571__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6767_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ _2611_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__o21ai_1
X_9555_ net423 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
X_5718_ _0937_ _1670_ _1669_ _0933_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8506_ _3963_ _3982_ _3985_ _3341_ _3979_ vssd1 vssd1 vccd1 vccd1 _3986_ sky130_fd_sc_hd__a221o_1
X_9486_ net361 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
X_6698_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[7\]
+ _2563_ net276 vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5649_ _1601_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold109_A team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8874__A2 _3543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7662__X _3252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8437_ net172 _3912_ _3915_ _3917_ vssd1 vssd1 vccd1 vccd1 _3918_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8368_ _3851_ _3852_ vssd1 vssd1 vccd1 vccd1 _3853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7319_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[6\]
+ _2986_ vssd1 vssd1 vccd1 vccd1 _2987_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_57_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8299_ _3501_ _3508_ _3515_ _0500_ vssd1 vssd1 vccd1 vccd1 _3792_ sky130_fd_sc_hd__o31ai_2
XANTENNA__6438__B net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9611__475 vssd1 vssd1 vccd1 vccd1 _9611__475/HI net475 sky130_fd_sc_hd__conb_1
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8653__B net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9286__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8372__C net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9505__380 vssd1 vssd1 vccd1 vccd1 _9505__380/HI net380 sky130_fd_sc_hd__conb_1
XFILLER_0_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5300__A1 _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_1
XFILLER_0_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4951_ _0731_ _0732_ _0733_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__a21o_1
XANTENNA__9448__Q team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4882_ net168 _0746_ _0743_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__a21o_4
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7670_ _3246_ _3251_ _3248_ vssd1 vssd1 vccd1 vccd1 _3260_ sky130_fd_sc_hd__mux2_1
X_6621_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[21\] _2513_
+ net260 vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_15_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5708__A _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9340_ clknet_leaf_3_wb_clk_i net2 net202 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.sync0
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6552_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[21\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[20\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[23\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[22\]
+ vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5503_ _1454_ _1455_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__nor2_1
XANTENNA__5119__A1 _0817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9271_ clknet_leaf_10_wb_clk_i _0080_ net226 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_6483_ net294 net298 vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__and2b_1
XANTENNA__7659__A3 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5434_ _1381_ _1383_ _1386_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__a21o_1
X_8222_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[12\]
+ _2990_ vssd1 vssd1 vccd1 vccd1 _3728_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8153_ _3672_ _3673_ vssd1 vssd1 vccd1 vccd1 _3674_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5365_ _1220_ _1317_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7104_ _0713_ _2840_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5296_ _1243_ _1245_ _1246_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__a21oi_1
X_8084_ _3607_ _3613_ net668 net244 vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_10_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7035_ _2782_ _2783_ net293 vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4758__A2_N net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8754__A _0423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8986_ net311 vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7937_ net333 net197 _3477_ net300 vssd1 vssd1 vccd1 vccd1 _3478_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7868_ net686 net166 _3427_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9607_ net471 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6819_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[5\]
+ _2644_ vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8544__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7799_ _3378_ _3384_ _2380_ vssd1 vssd1 vccd1 vccd1 _3385_ sky130_fd_sc_hd__mux2_1
X_9538_ net494 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9469_ net344 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_59_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8383__B _3261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7743__A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5263__A _1215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5150_ _1101_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5081_ _0996_ _1032_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8840_ net100 _4314_ _4317_ vssd1 vssd1 vccd1 vccd1 _4318_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5983_ _1898_ _1934_ _1933_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_56_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8771_ net100 _4238_ vssd1 vssd1 vccd1 vccd1 _4249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4934_ _0884_ _0886_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__nor2_1
X_7722_ _3289_ _3299_ vssd1 vssd1 vccd1 vccd1 _3312_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_19_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7637__B net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4865_ _0738_ _0809_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__nand2_4
XFILLER_0_75_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7653_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[6\]
+ net108 vssd1 vssd1 vccd1 vccd1 _3243_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout131_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4796_ _0743_ _0748_ _0745_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout229_A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6604_ _2503_ vssd1 vssd1 vccd1 vccd1 _2504_ sky130_fd_sc_hd__inv_2
X_7584_ net255 _2354_ net290 team_08_WB.instance_to_wrap.allocation.game.game.score\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_9323_ clknet_leaf_29_wb_clk_i _0006_ net237 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8829__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6535_ _2455_ _2456_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[14\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9254_ clknet_leaf_15_wb_clk_i _0092_ net216 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_65_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6466_ _0462_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[11\]
+ _2407_ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8205_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[6\]
+ _2986_ vssd1 vssd1 vccd1 vccd1 _3717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5417_ _1220_ _1317_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__or2_1
X_9185_ clknet_leaf_11_wb_clk_i _0048_ net219 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_6397_ team_08_WB.instance_to_wrap.allocation.game.game.score\[6\] team_08_WB.instance_to_wrap.allocation.game.game.score\[5\]
+ _2326_ _2335_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__a31o_1
X_5348_ _1297_ _1299_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8136_ net299 _3657_ _3658_ _3661_ vssd1 vssd1 vccd1 vccd1 _3662_ sky130_fd_sc_hd__a31o_1
X_8067_ _3598_ vssd1 vssd1 vccd1 vccd1 _3599_ sky130_fd_sc_hd__inv_2
X_5279_ _1228_ _1231_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__xor2_1
XANTENNA__5276__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7018_ _0453_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[2\]
+ _2768_ vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4517__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7973__C1 _3511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_8969_ net278 _4443_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_92_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4650_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[6\] vssd1
+ vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__nand2b_1
Xinput10 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_1
Xinput21 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput32 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
X_4581_ _0495_ _0541_ _0545_ _0547_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6320_ net330 _2267_ _2271_ net327 _2270_ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5264__Y _1217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6251_ _1879_ _2124_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6182_ _2132_ _2134_ _1596_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__a21bo_1
X_5202_ _1154_ _1152_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5133_ _1084_ _1085_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5721__A _1645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5064_ _1015_ _1016_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8823_ _0423_ net105 vssd1 vssd1 vccd1 vccd1 _4301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5966_ _1873_ _1874_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8754_ _0423_ _4212_ vssd1 vssd1 vccd1 vccd1 _4232_ sky130_fd_sc_hd__nor2_2
X_4917_ _0868_ _0869_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5897_ _1847_ _1849_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7367__B net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7705_ net175 _3289_ vssd1 vssd1 vccd1 vccd1 _3295_ sky130_fd_sc_hd__nor2_1
X_8685_ net133 _4156_ _4161_ _4163_ vssd1 vssd1 vccd1 vccd1 _4164_ sky130_fd_sc_hd__o211a_1
X_4848_ _0799_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7636_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[8\]
+ net117 vssd1 vssd1 vccd1 vccd1 _3226_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7567_ net540 team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr1\[1\] vssd1
+ vssd1 vccd1 vccd1 _3169_ sky130_fd_sc_hd__nand2_1
X_4779_ _0615_ _0628_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__xnor2_4
X_9306_ clknet_leaf_2_wb_clk_i _0277_ net204 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.game.score\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6518_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[9\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[8\]
+ _2441_ vssd1 vssd1 vccd1 vccd1 _2445_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7498_ _3135_ _3136_ net114 vssd1 vssd1 vccd1 vccd1 _3137_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9237_ clknet_leaf_21_wb_clk_i _0052_ net239 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_6449_ _2384_ _2395_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9168_ _0143_ _0418_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_12_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8119_ net162 _3630_ vssd1 vssd1 vccd1 vccd1 _3646_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9099_ clknet_leaf_52_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[29\]
+ net207 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5350__B _1011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6749__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7740__B _3329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8426__B1 _3280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8852__A _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7739__Y _3329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7937__C1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5820_ _1770_ _1771_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_33_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5751_ _1012_ _1694_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8470_ _3878_ _3893_ _3906_ _3919_ _3354_ vssd1 vssd1 vccd1 vccd1 _3951_ sky130_fd_sc_hd__o41a_1
X_4702_ _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__inv_2
X_5682_ _1587_ _1634_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8901__A1 _3271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7421_ net312 _3022_ vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4633_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[1\] vssd1
+ vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__xnor2_4
X_4564_ _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__inv_2
X_7352_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\] _3011_
+ _2974_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__mux2_1
X_6303_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[20\]
+ _2191_ _2194_ _2255_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__a211o_1
X_7283_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[19\]
+ _2960_ net180 vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6234_ _2143_ _2186_ vssd1 vssd1 vccd1 vccd1 _2187_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4495_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] vssd1 vssd1 vccd1
+ vccd1 _0467_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7931__A _0522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9022_ clknet_leaf_53_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[4\]
+ net201 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6165_ _2054_ _2063_ _2064_ _2117_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout296_A team_08_WB.instance_to_wrap.allocation.game.controller.state\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5116_ _1068_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__inv_2
X_6096_ _2021_ _2048_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5047_ _0820_ _0867_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_34_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_49_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6998_ _0467_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] _2758_ _2761_
+ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__a31oi_1
X_8806_ net313 net99 vssd1 vssd1 vccd1 vccd1 _4284_ sky130_fd_sc_hd__nand2_1
X_5949_ _1855_ _1900_ _1899_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_66_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8737_ net188 _3486_ _3763_ vssd1 vssd1 vccd1 vccd1 _4215_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8668_ _4110_ _4112_ vssd1 vssd1 vccd1 vccd1 _4147_ sky130_fd_sc_hd__nor2_1
XANTENNA__5706__A1 _1645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4801__Y _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7619_ _3204_ _3208_ vssd1 vssd1 vccd1 vccd1 _3209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8599_ net111 _4076_ _4077_ net116 vssd1 vssd1 vccd1 vccd1 _4078_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_90_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4530__A _0423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8496__X _3976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input24_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9541__409 vssd1 vssd1 vccd1 vccd1 _9541__409/HI net409 sky130_fd_sc_hd__conb_1
XFILLER_0_86_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7395__B1 _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8344__C1 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5271__A _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6086__B _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7970_ _0487_ _3500_ _3493_ vssd1 vssd1 vccd1 vccd1 _3509_ sky130_fd_sc_hd__mux2_1
X_6921_ net272 _2712_ _2713_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__nor3_1
XFILLER_0_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9640_ net487 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
X_6852_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7386__B1 _3034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9571_ net436 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
X_9481__356 vssd1 vssd1 vccd1 vccd1 _9481__356/HI net356 sky130_fd_sc_hd__conb_1
X_5803_ net141 _0930_ _1755_ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6783_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[7\]
+ _2620_ net274 vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_44_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8522_ _3340_ _4000_ vssd1 vssd1 vccd1 vccd1 _4001_ sky130_fd_sc_hd__and2_2
X_5734_ _1685_ _1686_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5665_ net128 _1617_ _1616_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__a21bo_1
X_9522__397 vssd1 vssd1 vccd1 vccd1 _9522__397/HI net397 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_40_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8453_ _3872_ _3933_ _3891_ vssd1 vssd1 vccd1 vccd1 _3934_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4616_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[7\] vssd1
+ vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_40_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7404_ _0437_ net301 vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__nand2_1
X_8384_ _3241_ _3864_ vssd1 vssd1 vccd1 vccd1 _3865_ sky130_fd_sc_hd__nand2_2
XFILLER_0_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5596_ _1543_ _1545_ _1547_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_92_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7335_ net501 net121 vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__nor2_1
XANTENNA__9333__RESET_B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4500__D net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4547_ net292 _0420_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.button
+ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__and3_1
XANTENNA__8757__A _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6113__A1 _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4478_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[0\] vssd1 vssd1
+ vccd1 vccd1 _0450_ sky130_fd_sc_hd__inv_2
X_7266_ _2950_ vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6217_ _2168_ _2169_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__xnor2_1
X_9005_ clknet_leaf_4_wb_clk_i _0169_ net203 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_7197_ net594 _2900_ _2901_ net164 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__a211oi_1
X_6148_ _2090_ _2091_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__xor2_1
X_6079_ _2029_ _2030_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4525__A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9074__RESET_B net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7571__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5803__B _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7368__B1 _2423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5450_ _1399_ _1401_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5556__A_N net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5381_ _1315_ _1333_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6649__X _2532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7120_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[11\] _2848_
+ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__and3_1
Xfanout219 net221 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_4
X_7051_ _2790_ _2794_ vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__nor2_2
XFILLER_0_10_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout208 net210 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dlymetal6s2s_1
X_6002_ _1916_ _1917_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7953_ _3491_ _3492_ vssd1 vssd1 vccd1 vccd1 _3493_ sky130_fd_sc_hd__or2_1
X_9563__431 vssd1 vssd1 vccd1 vccd1 _9563__431/HI net431 sky130_fd_sc_hd__conb_1
X_6904_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[5\]
+ _2700_ net267 vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__o21ai_1
X_7884_ _3403_ _3437_ _3438_ _3402_ net663 vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8020__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout259_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9623_ net264 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
X_6835_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[10\]
+ _2653_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9554_ net422 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
X_6766_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ _2611_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__and2b_1
X_5717_ _0927_ _0928_ _0930_ _0922_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__o31a_1
X_8505_ _3872_ _3976_ _3984_ _3905_ _3983_ vssd1 vssd1 vccd1 vccd1 _3985_ sky130_fd_sc_hd__a221o_1
X_9485_ net360 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6697_ _2563_ _2564_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5648_ _1559_ _1561_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8436_ _3865_ _3869_ _3916_ net174 vssd1 vssd1 vccd1 vccd1 _3917_ sky130_fd_sc_hd__o31a_1
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5579_ _1502_ _1504_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8367_ net289 _3471_ vssd1 vssd1 vccd1 vccd1 _3852_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4896__B2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8298_ net196 _3790_ _3788_ net170 vssd1 vssd1 vccd1 vccd1 _3791_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7318_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[5\]
+ _2985_ vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7249_ _2938_ _2939_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8653__C _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8154__A1_N _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8950__A _3864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6325__B2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6325__A1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5300__A2 _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_0__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9547__415 vssd1 vssd1 vccd1 vccd1 _9547__415/HI net415 sky130_fd_sc_hd__conb_1
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4950_ _0901_ _0902_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4811__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4881_ _0832_ _0833_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6620_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[21\] _2513_
+ vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_15_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6551_ net529 _2464_ _2466_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[20\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5502_ _1444_ _1453_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4612__B _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9270_ clknet_leaf_10_wb_clk_i _0079_ net226 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6482_ net295 net296 _2420_ _2421_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__a211o_1
X_9593__457 vssd1 vssd1 vccd1 vccd1 _9593__457/HI net457 sky130_fd_sc_hd__conb_1
X_5433_ _1385_ _1384_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8221_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[2\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ net122 vssd1 vssd1 vccd1 vccd1 _3727_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5724__A _0939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5364_ _0998_ _1222_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8069__A1 _3597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8100__A _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8152_ _0662_ net183 vssd1 vssd1 vccd1 vccd1 _3673_ sky130_fd_sc_hd__and2_1
XANTENNA__7816__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7103_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.state\[1\]
+ _2841_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5295_ _1247_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8083_ _0430_ _3608_ _3609_ _3612_ net238 vssd1 vssd1 vccd1 vccd1 _3613_ sky130_fd_sc_hd__o2111a_1
X_7034_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\]
+ _0457_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\] vssd1
+ vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_87_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9487__362 vssd1 vssd1 vccd1 vccd1 _9487__362/HI net362 sky130_fd_sc_hd__conb_1
XFILLER_0_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8985_ net312 vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7936_ net197 _3475_ vssd1 vssd1 vccd1 vccd1 _3477_ sky130_fd_sc_hd__nand2_1
XANTENNA__8770__A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7867_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[10\]
+ _3424_ _3426_ vssd1 vssd1 vccd1 vccd1 _3427_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9606_ net470 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
XANTENNA__4803__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6818_ _2644_ _2645_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7798_ _2361_ _3381_ _3383_ _2363_ _2358_ vssd1 vssd1 vccd1 vccd1 _3384_ sky130_fd_sc_hd__o32a_1
X_9537_ net493 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_73_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6749_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[10\]
+ _2597_ net273 vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9323__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9468_ net343 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8929__B _3265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8419_ _3344_ _3898_ _3899_ _3896_ vssd1 vssd1 vccd1 vccd1 _3900_ sky130_fd_sc_hd__a31o_1
X_9399_ clknet_leaf_31_wb_clk_i _0346_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8664__B _3608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5046__A1 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7743__B net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8855__A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5080_ _0996_ _1032_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8066__S team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9459__Q team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_cactus vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5982_ _1898_ _1933_ _1934_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__nand3_1
X_8770_ net105 _4246_ vssd1 vssd1 vccd1 vccd1 _4248_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8590__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4933_ _0850_ _0883_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__and2_1
X_7721_ _3304_ _3310_ _3298_ vssd1 vssd1 vccd1 vccd1 _3311_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4864_ net144 _0810_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__nor2_1
XANTENNA__8931__C1 _4407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7652_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[6\]
+ _3230_ _3238_ _3240_ vssd1 vssd1 vccd1 vccd1 _3242_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4795_ _0724_ _0740_ _0747_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__mux2_4
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6603_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[15\] _2502_
+ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__and2_1
X_7583_ net260 _2358_ _0420_ team_08_WB.instance_to_wrap.allocation.game.game.score\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_28_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9322_ clknet_leaf_31_wb_clk_i _0005_ net244 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_31_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6534_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[14\] _2453_
+ net156 vssd1 vssd1 vccd1 vccd1 _2456_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout124_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9253_ clknet_leaf_15_wb_clk_i _0104_ net216 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_6465_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[16\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[15\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__nand3_1
XANTENNA__7653__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5416_ _1368_ _1367_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8204_ _3031_ _3716_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9184_ clknet_leaf_11_wb_clk_i _0047_ net226 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6396_ team_08_WB.instance_to_wrap.allocation.game.game.score\[6\] team_08_WB.instance_to_wrap.allocation.game.game.score\[5\]
+ _2326_ _2335_ vssd1 vssd1 vccd1 vccd1 _2347_ sky130_fd_sc_hd__a31oi_4
X_5347_ _1245_ _1297_ _1298_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_54_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8135_ net296 _3659_ _3660_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[0\]
+ _3597_ vssd1 vssd1 vccd1 vccd1 _3661_ sky130_fd_sc_hd__a311o_1
XFILLER_0_11_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5278_ _1229_ _1230_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__nor2_1
X_8066_ _0654_ net161 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _3598_ sky130_fd_sc_hd__mux2_1
XANTENNA__8462__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7017_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[1\] team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\]
+ _2772_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__or3_1
XANTENNA__4517__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8968_ _4442_ _4444_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7919_ net335 _0552_ net197 vssd1 vssd1 vccd1 vccd1 _3461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8899_ net187 _2271_ _4375_ vssd1 vssd1 vccd1 vccd1 _4376_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8005__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9576__441 vssd1 vssd1 vccd1 vccd1 _9576__441/HI net441 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_78_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5364__A _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8150__B1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5267__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5539__A _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput22 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_2
Xinput11 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4580_ net329 _0546_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__nand2_1
XANTENNA__4730__X _0685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput33 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5274__A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8141__B1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6250_ _0447_ _2202_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6181_ _1596_ _2133_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__and2_1
X_5201_ _1098_ _1153_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8585__A _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5132_ _1073_ _1077_ _1083_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__nor3_1
XFILLER_0_23_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5063_ _1011_ _1014_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8822_ net326 _0425_ _4299_ vssd1 vssd1 vccd1 vccd1 _4300_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7000__Y net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5965_ _1916_ _1917_ _1915_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8753_ _4211_ _4219_ _4229_ _4230_ _4225_ vssd1 vssd1 vccd1 vccd1 _4231_ sky130_fd_sc_hd__o41ai_1
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4916_ _0803_ _0861_ _0867_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__nor3_1
X_5896_ net147 _0927_ _1847_ _1848_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__nand4_1
XANTENNA_fanout241_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7704_ net174 _3292_ vssd1 vssd1 vccd1 vccd1 _3294_ sky130_fd_sc_hd__or2_1
X_8684_ net149 _4160_ _4162_ vssd1 vssd1 vccd1 vccd1 _4163_ sky130_fd_sc_hd__o21ba_1
X_9599__463 vssd1 vssd1 vccd1 vccd1 _9599__463/HI net463 sky130_fd_sc_hd__conb_1
X_4847_ _0797_ _0798_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7635_ net119 vssd1 vssd1 vccd1 vccd1 _3225_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4778_ _0729_ _0730_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__and2_4
X_7566_ net540 _2693_ _3015_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8479__B _3864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9305_ clknet_leaf_1_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.collides
+ net209 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.col
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_95_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6517_ _2443_ _2444_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[8\]
+ sky130_fd_sc_hd__nor2_1
X_7497_ net301 _3100_ _3133_ _3101_ _3059_ vssd1 vssd1 vccd1 vccd1 _3136_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9236_ clknet_leaf_21_wb_clk_i _0051_ net239 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4664__A_N team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6448_ _2393_ net299 net295 vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9167_ _0142_ _0417_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_12_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6379_ team_08_WB.instance_to_wrap.allocation.game.game.score\[5\] team_08_WB.instance_to_wrap.allocation.game.game.score\[4\]
+ _2328_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8118_ net162 _3630_ vssd1 vssd1 vccd1 vccd1 _3645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9098_ clknet_leaf_53_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[28\]
+ net200 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_8049_ _0570_ _3567_ _3582_ net195 vssd1 vssd1 vccd1 vccd1 _3584_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8006__Y _3543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8426__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5750_ _0835_ _1695_ _1702_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_33_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5681_ _1585_ _1586_ _1579_ _1581_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4701_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__xor2_4
XFILLER_0_17_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4632_ _0589_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__inv_2
X_7420_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_dino _3064_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_cactus
+ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_72_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4563_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[19\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[20\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[18\] vssd1 vssd1 vccd1
+ vccd1 _0532_ sky130_fd_sc_hd__or3b_1
X_7351_ _3010_ _3009_ vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6302_ _2195_ _2197_ _2198_ _2254_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__or4b_1
X_4494_ net633 vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__inv_2
X_7282_ _2960_ _2961_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6233_ _2140_ _2142_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9021_ clknet_leaf_0_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[3\]
+ net201 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6164_ _2065_ _2115_ _2116_ vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__and3_1
X_5115_ _1029_ _1066_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__nor2_1
X_6095_ _2046_ _2047_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout191_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5046_ _0743_ _0797_ _0969_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__a21oi_2
XANTENNA__9192__RESET_B net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout289_A team_08_WB.instance_to_wrap.allocation.game.controller.v\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9527__402 vssd1 vssd1 vccd1 vccd1 _9527__402/HI net402 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_49_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8107__X _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6563__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6997_ _2758_ _2760_ _0467_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8805_ net313 _3266_ vssd1 vssd1 vccd1 vccd1 _4283_ sky130_fd_sc_hd__and2_1
X_5948_ _1855_ _1899_ _1900_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_66_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8736_ _3486_ _3763_ net188 vssd1 vssd1 vccd1 vccd1 _4214_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5879_ _1828_ _1831_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__nor2_1
XANTENNA__5907__A _0919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8667_ _4142_ _4145_ vssd1 vssd1 vccd1 vccd1 _4146_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7618_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[9\]
+ _3191_ vssd1 vssd1 vccd1 vccd1 _3208_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8598_ net183 _4075_ _4061_ vssd1 vssd1 vccd1 vccd1 _4077_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7549_ net617 team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr2\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr2\[0\] vssd1 vssd1 vccd1
+ vccd1 _3160_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4530__B net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7681__X _3271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9219_ clknet_leaf_17_wb_clk_i _0076_ net230 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8959__A2 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input17_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7919__A0 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7395__A1 _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5089__A _1039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8344__B1 _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8895__B2 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5095__Y _1048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8647__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7083__B1 _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6920_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[10\]
+ _2709_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6851_ net269 _2661_ _2667_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4615__B team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7386__A1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9570_ net498 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
X_5802_ net147 _0928_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6782_ _2620_ _2621_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8521_ _0555_ _3339_ _3999_ vssd1 vssd1 vccd1 vccd1 _4000_ sky130_fd_sc_hd__o21ai_1
X_5733_ _1630_ _1631_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5664_ _1614_ _1615_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_40_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8452_ net175 _3884_ _3888_ _3931_ vssd1 vssd1 vccd1 vccd1 _3933_ sky130_fd_sc_hd__a31o_1
X_5595_ _1543_ _1545_ _1547_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__o21ai_1
X_4615_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[8\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[8\] vssd1
+ vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__and2b_2
X_7403_ _0439_ _0441_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__nor2_1
X_8383_ net107 _3261_ vssd1 vssd1 vccd1 vccd1 _3864_ sky130_fd_sc_hd__nor2_2
XFILLER_0_25_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4546_ net292 _0420_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__nand2_2
X_7334_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[22\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[23\]
+ _2999_ vssd1 vssd1 vccd1 vccd1 _3002_ sky130_fd_sc_hd__or3_2
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout204_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4477_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[0\] vssd1 vssd1
+ vccd1 vccd1 _0449_ sky130_fd_sc_hd__inv_2
X_7265_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[12\]
+ _2946_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__and3_1
XANTENNA__9373__RESET_B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6216_ _2164_ _2167_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__xnor2_1
X_7196_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[15\] _2900_ vssd1
+ vssd1 vccd1 vccd1 _2901_ sky130_fd_sc_hd__nor2_1
X_9004_ clknet_leaf_4_wb_clk_i _0168_ net203 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input9_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6147_ _2098_ _2099_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__and2b_1
XANTENNA__9302__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6078_ _2029_ _2030_ vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__nand2_1
X_5029_ _0837_ _0887_ _0861_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7676__X _3266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8719_ net324 _3775_ vssd1 vssd1 vccd1 vccd1 _4197_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_81_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8877__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5372__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4716__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6650__B _2532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4451__A team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5380_ _1312_ _1314_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8096__A2 _3622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7481__B team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_cactus vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7050_ _2797_ vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_4
X_6001_ _1948_ _1950_ _1953_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7952_ _0494_ _3490_ vssd1 vssd1 vccd1 vccd1 _3492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6903_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[5\]
+ _2700_ vssd1 vssd1 vccd1 vccd1 _2702_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_9622_ net265 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
X_7883_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[15\]
+ _3435_ vssd1 vssd1 vccd1 vccd1 _3438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8556__B1 _4001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6834_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[10\]
+ _2653_ _2655_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__o21a_1
XANTENNA__8020__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout154_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9553_ net421 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
X_6765_ net274 _2610_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9484_ net359 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
X_5716_ _0923_ _1668_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout321_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8504_ net154 _3959_ vssd1 vssd1 vccd1 vccd1 _3984_ sky130_fd_sc_hd__or2_1
X_6696_ net619 _2562_ net267 vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8435_ _3225_ net112 vssd1 vssd1 vccd1 vccd1 _3916_ sky130_fd_sc_hd__nand2_2
X_5647_ _1562_ _1563_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5578_ _1525_ _1529_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__nand2_1
X_8366_ net289 _3471_ vssd1 vssd1 vccd1 vccd1 _3851_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4896__A2 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4529_ _0423_ net289 vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__nor2_1
X_8297_ net324 _3776_ vssd1 vssd1 vccd1 vccd1 _3790_ sky130_fd_sc_hd__xnor2_1
X_7317_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[4\]
+ _2984_ vssd1 vssd1 vccd1 vccd1 _2985_ sky130_fd_sc_hd__or2_1
XANTENNA__5192__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7248_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[7\]
+ _2936_ net179 vssd1 vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__o21ai_1
X_7179_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[8\] _2887_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2890_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4536__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9295__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4880_ _0807_ _0831_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_15_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4452__Y _0425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5277__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6550_ net529 _2464_ net156 vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5501_ _1405_ _1443_ _1453_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6481_ net280 net296 _2391_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__and3_1
XANTENNA__7513__A1 _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7492__A _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5432_ _1381_ _1383_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__xnor2_2
X_8220_ _3035_ _3726_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__nand2_1
X_5363_ _0998_ _1222_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_39_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8151_ _0662_ net183 vssd1 vssd1 vccd1 vccd1 _3672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7102_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[1\] team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[2\]
+ _2776_ _2840_ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__a311o_1
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5294_ _1243_ _1245_ _1246_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__and3_1
XANTENNA__9275__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8082_ _0705_ _3611_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3612_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4908__X _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7033_ _2780_ _2781_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[3\]
+ _0458_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_93_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5053__A_N _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout271_A _2548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8984_ net312 vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7935_ _3475_ vssd1 vssd1 vccd1 vccd1 _3476_ sky130_fd_sc_hd__inv_2
X_7866_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[10\]
+ _3424_ net160 vssd1 vssd1 vccd1 vccd1 _3426_ sky130_fd_sc_hd__o21ai_1
X_9605_ net469 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6817_ net629 _2642_ net271 vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9536_ net492 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XANTENNA__4803__B net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7797_ _2358_ _2373_ _3382_ _2350_ vssd1 vssd1 vccd1 vccd1 _3383_ sky130_fd_sc_hd__o211a_1
X_6748_ _2597_ _2598_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__nor2_1
XANTENNA__6960__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9467_ net342 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6679_ _2549_ _2550_ _2551_ _2552_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__or4_2
XFILLER_0_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9398_ clknet_leaf_31_wb_clk_i _0345_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_8418_ _3290_ _3880_ vssd1 vssd1 vccd1 vccd1 _3899_ sky130_fd_sc_hd__or2_1
XANTENNA__9390__Q team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8349_ _0702_ _2279_ _3833_ net298 _3838_ vssd1 vssd1 vccd1 vccd1 _3839_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_76_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7807__A2 _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5650__A _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6481__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4553__X _0522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5097__A _1048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8871__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5981_ _1895_ _1897_ _1896_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4932_ _0884_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__inv_2
XANTENNA__4796__A1 _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7720_ net135 _3303_ _3305_ _3309_ vssd1 vssd1 vccd1 vccd1 _3310_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7651_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[6\]
+ _3230_ _3238_ _3240_ vssd1 vssd1 vccd1 vccd1 _3241_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4863_ _0783_ _0793_ _0808_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6602_ _2502_ net262 _2501_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[14\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_28_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9601__465 vssd1 vssd1 vccd1 vccd1 _9601__465/HI net465 sky130_fd_sc_hd__conb_1
XFILLER_0_90_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4794_ _0719_ net144 _0743_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__or3_4
XFILLER_0_6_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7582_ net291 team_08_WB.instance_to_wrap.allocation.game.game.score\[2\] net259
+ _2371_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9321_ clknet_leaf_29_wb_clk_i _0000_ net237 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_31_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6533_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[13\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[14\]
+ _2451_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__and3_1
X_9252_ clknet_leaf_15_wb_clk_i _0103_ net215 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_6464_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[12\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5415_ _0959_ _1222_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8203_ _2986_ _3715_ net121 vssd1 vssd1 vccd1 vccd1 _3716_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout117_A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9183_ clknet_leaf_10_wb_clk_i _0046_ net226 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_28_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_6395_ _2330_ _2345_ vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5346_ _1245_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8134_ net280 _0642_ _2386_ vssd1 vssd1 vccd1 vccd1 _3660_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5277_ net123 _1205_ _1207_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__and3_1
X_8065_ net298 net278 _2427_ vssd1 vssd1 vccd1 vccd1 _3597_ sky130_fd_sc_hd__or3_4
XANTENNA__6566__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7016_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[6\] _2771_
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[3\] vssd1 vssd1
+ vccd1 vccd1 _2772_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_71_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7973__A1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8967_ net258 net277 _3279_ _4443_ vssd1 vssd1 vccd1 vccd1 _4444_ sky130_fd_sc_hd__or4b_1
XANTENNA__4814__A _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7918_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] team_08_WB.instance_to_wrap.allocation.game.controller.v\[2\]
+ _3458_ vssd1 vssd1 vccd1 vccd1 _3460_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8898_ net190 _2267_ _2271_ net187 _4374_ vssd1 vssd1 vccd1 vccd1 _4375_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7849_ _3413_ vssd1 vssd1 vccd1 vccd1 _3414_ sky130_fd_sc_hd__inv_2
XANTENNA__8005__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4820__Y _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9519_ net394 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_78_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5267__A2 _1215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7008__A3 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput34 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput23 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7770__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6180_ _1591_ _1593_ _1595_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__nand3_1
X_5200_ _0867_ _1097_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5131_ _1073_ _1077_ _1083_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5062_ _1011_ _1014_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6673__X _2547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8821_ _4292_ _4298_ vssd1 vssd1 vccd1 vccd1 _4299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8752_ _4213_ _4222_ vssd1 vssd1 vccd1 vccd1 _4230_ sky130_fd_sc_hd__or2_1
XANTENNA__5449__B _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5964_ _1880_ _1914_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7703_ net174 _3292_ vssd1 vssd1 vccd1 vccd1 _3293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4915_ _0861_ _0867_ _0803_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5895_ _0772_ _0930_ _1846_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8683_ _4119_ _4158_ _4124_ vssd1 vssd1 vccd1 vccd1 _4162_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4846_ _0798_ _0797_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout234_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7634_ _3221_ _3223_ vssd1 vssd1 vccd1 vccd1 _3224_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_99_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7565_ net617 _2554_ _3015_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4777_ _0618_ _0627_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__xnor2_4
X_9304_ clknet_leaf_5_wb_clk_i _0019_ net204 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.slow_clk
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6516_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[8\] _2441_
+ _2429_ vssd1 vssd1 vccd1 vccd1 _2444_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7496_ _3134_ _3023_ _3024_ vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__or3b_1
XFILLER_0_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9235_ clknet_leaf_21_wb_clk_i _0050_ net242 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_6447_ net296 _2392_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9166_ _0141_ _0416_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_6378_ team_08_WB.instance_to_wrap.allocation.game.game.score\[4\] _2328_ vssd1 vssd1
+ vccd1 vccd1 _2329_ sky130_fd_sc_hd__nand2_1
X_9536__492 vssd1 vssd1 vccd1 vccd1 net492 _9536__492/LO sky130_fd_sc_hd__conb_1
XFILLER_0_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5329_ _1279_ _1280_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__nand2b_1
X_8117_ _3628_ _3642_ _3643_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3644_ sky130_fd_sc_hd__o211a_1
XANTENNA__4809__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9097_ clknet_leaf_52_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[27\]
+ net209 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_8048_ _3567_ _3582_ _0570_ vssd1 vssd1 vccd1 vccd1 _3583_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9068__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8371__B2 team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_3__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5822__B _1774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7749__B net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7937__A1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9274__SET_B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _1629_ _1632_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__nor2_1
X_4700_ net576 net295 _0638_ _0655_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4741__X _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4631_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[0\] vssd1
+ vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_44_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7350_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr1\[0\] team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__xnor2_1
X_4562_ _0530_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6301_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[17\]
+ _2199_ _2253_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__o21ba_1
X_4493_ net646 vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__inv_2
X_7281_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[18\]
+ _2958_ net180 vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__o21ai_1
X_6232_ _2144_ _2184_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9020_ clknet_leaf_0_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[2\]
+ net206 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6163_ _2054_ _2064_ _2063_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5114_ _1029_ _1066_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__nand2_1
X_6094_ _2015_ _2017_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5045_ _0794_ _0856_ _0961_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6563__B _2477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6996_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2760_ sky130_fd_sc_hd__nand2_1
XANTENNA__6282__C _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8804_ net175 _3335_ _3888_ _4281_ vssd1 vssd1 vccd1 vccd1 _4282_ sky130_fd_sc_hd__a31o_1
X_9607__471 vssd1 vssd1 vccd1 vccd1 _9607__471/HI net471 sky130_fd_sc_hd__conb_1
X_5947_ _1852_ _1854_ _1853_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_66_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8735_ net186 _3775_ _4212_ vssd1 vssd1 vccd1 vccd1 _4213_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8666_ _4143_ _4144_ vssd1 vssd1 vccd1 vccd1 _4145_ sky130_fd_sc_hd__and2_1
X_5878_ _1829_ _1830_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout237_X net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7617_ _3190_ _3205_ vssd1 vssd1 vccd1 vccd1 _3207_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4829_ _0776_ _0780_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_8597_ _0661_ _3595_ _4075_ vssd1 vssd1 vccd1 vccd1 _4076_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_65_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7548_ net257 _3159_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7479_ net114 _3119_ vssd1 vssd1 vccd1 vccd1 _3120_ sky130_fd_sc_hd__nand2_1
X_9218_ clknet_leaf_19_wb_clk_i _0075_ net229 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9149_ clknet_leaf_36_wb_clk_i net506 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9249__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7919__A1 _0552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4545__Y _0514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8041__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8895__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5833__A _1074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7524__S team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4449__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7083__B2 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8355__S team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 team_08_WB.instance_to_wrap.allocation.game.sync0 vssd1 vssd1 vccd1 vccd1 net499
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6850_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__nand2_1
XANTENNA__8032__B1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7386__A2 _3022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5801_ _1703_ _1704_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__xnor2_2
X_6781_ net634 _2619_ net270 vssd1 vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5732_ _1678_ _1682_ _1683_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8520_ net191 _0556_ net105 net103 vssd1 vssd1 vccd1 vccd1 _3999_ sky130_fd_sc_hd__a31o_1
XANTENNA__8335__A1 _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5663_ _1615_ _1614_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_73_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8451_ _3931_ vssd1 vssd1 vccd1 vccd1 _3932_ sky130_fd_sc_hd__inv_2
X_5594_ _1490_ _1546_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4614_ net313 _0540_ _0572_ net261 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[7\]
+ sky130_fd_sc_hd__o211a_1
X_7402_ _3025_ _3043_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_13_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8382_ _3859_ _3862_ vssd1 vssd1 vccd1 vccd1 _3863_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7333_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[23\]
+ _3000_ vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4545_ _0419_ net290 vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__nor2_2
XFILLER_0_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5743__A _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_29_wb_clk_i_X clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4476_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__inv_2
X_9003_ clknet_leaf_4_wb_clk_i _0167_ net203 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__7310__A2 _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7264_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[12\]
+ _2946_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6215_ _2162_ _2166_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__xnor2_1
X_7195_ net164 _2899_ _2900_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_2__f_wb_clk_i_X clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6146_ _2087_ _2089_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_0_wb_clk_i_X clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6077_ _1989_ _1990_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout187_X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5028_ _0979_ _0980_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8023__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6979_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[21\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[20\]
+ _2744_ _0019_ vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8718_ net260 net208 _4196_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6337__B1 _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8877__A2 _3542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8649_ _2537_ net119 vssd1 vssd1 vccd1 vccd1 _4128_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8317__B2 _3543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5303__A1 _1039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6000_ _1951_ _1952_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__nor2_1
XANTENNA__8253__B1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7951_ _0550_ _3490_ _3482_ vssd1 vssd1 vccd1 vccd1 _3491_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_94_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7882_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[15\]
+ _3435_ vssd1 vssd1 vccd1 vccd1 _3437_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6902_ _2700_ _2701_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__nor2_1
XANTENNA__7777__X _3367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9621_ net264 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
X_6833_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[10\]
+ _2653_ net275 vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__a21oi_1
XANTENNA__7359__A2 _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout147_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9552_ net420 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
X_6764_ _2609_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5715_ _1662_ _1664_ _1667_ _0933_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__o31a_1
X_6695_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[6\]
+ _2562_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__and2_1
X_9483_ net358 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8503_ _3290_ _3302_ _3313_ _3974_ net171 vssd1 vssd1 vccd1 vccd1 _3983_ sky130_fd_sc_hd__o311a_1
X_5646_ _1578_ _1598_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout314_A team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8434_ _3290_ _3302_ _3364_ _3914_ vssd1 vssd1 vccd1 vccd1 _3915_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7672__B _3261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5577_ _1525_ _1529_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__or2_1
X_8365_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] _2874_ _3850_
+ _0561_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__o22a_1
X_4528_ _0487_ _0496_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__nand2_1
X_8296_ net329 _3525_ vssd1 vssd1 vccd1 vccd1 _3789_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout102_X net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7316_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[3\]
+ _2983_ vssd1 vssd1 vccd1 vccd1 _2984_ sky130_fd_sc_hd__or2_1
XANTENNA__5192__B _1144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4459_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _0431_ sky130_fd_sc_hd__inv_2
XANTENNA__8784__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8492__B1 _3971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7247_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[7\]
+ _2936_ vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_57_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7178_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[8\] _2887_ _2889_
+ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6129_ _2080_ _2081_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8795__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4536__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7687__X _3277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8024__A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4552__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6479__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9471__346 vssd1 vssd1 vccd1 vccd1 _9471__346/HI net346 sky130_fd_sc_hd__conb_1
XANTENNA__6485__Y _2423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4727__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9512__387 vssd1 vssd1 vccd1 vccd1 _9512__387/HI net387 sky130_fd_sc_hd__conb_1
XANTENNA__6797__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5558__A _0814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5500_ _0747_ _1452_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8869__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6480_ net295 net137 vssd1 vssd1 vccd1 vccd1 _2420_ sky130_fd_sc_hd__nor2_1
XANTENNA__5293__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5431_ _1355_ _1376_ _1378_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__a21o_2
XFILLER_0_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5362_ _1312_ _1314_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__and2_1
X_8150_ _3669_ _3670_ _3671_ net237 net578 vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_39_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7101_ _2836_ _2839_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8081_ _3610_ vssd1 vssd1 vccd1 vccd1 _3611_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5293_ net129 _1186_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__xnor2_1
X_7032_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[1\] vssd1
+ vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__nand2_2
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8983_ net312 vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7934_ _0491_ _0550_ vssd1 vssd1 vccd1 vccd1 _3475_ sky130_fd_sc_hd__xor2_2
XANTENNA__7300__X _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7865_ _3424_ _3425_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[9\]
+ net166 vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__a2bb2o_1
X_9604_ net468 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_93_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5468__A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6816_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[4\]
+ _2641_ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7796_ _2358_ _2373_ vssd1 vssd1 vccd1 vccd1 _3382_ sky130_fd_sc_hd__nand2_1
X_9535_ net491 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6747_ net690 _2596_ net269 vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6678_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8162__C1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9466_ net341 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
X_5629_ _1572_ _1580_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5915__B _1867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6712__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9397_ clknet_leaf_31_wb_clk_i _0344_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_8417_ _3289_ _3296_ _3884_ _3897_ vssd1 vssd1 vccd1 vccd1 _3898_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8348_ _3511_ _3837_ _3834_ _3479_ vssd1 vssd1 vccd1 vccd1 _3838_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8279_ _3492_ _3520_ _3760_ net196 vssd1 vssd1 vccd1 vccd1 _3773_ sky130_fd_sc_hd__a31o_1
XANTENNA__5650__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4547__A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9445__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9553__421 vssd1 vssd1 vccd1 vccd1 _9553__421/HI net421 sky130_fd_sc_hd__conb_1
XFILLER_0_32_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7532__S team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6656__B _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_16_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7768__A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5980_ net148 _0922_ _1932_ _1930_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4931_ _0850_ _0883_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__nor2_1
XANTENNA__4796__A2 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4862_ _0783_ _0793_ _0814_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__o21ai_4
X_7650_ _3231_ _3239_ vssd1 vssd1 vccd1 vccd1 _3240_ sky130_fd_sc_hd__and2_1
X_6601_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[13\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[14\]
+ _2498_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_25_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4793_ _0719_ _0738_ _0744_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__and3b_4
XFILLER_0_55_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9320_ clknet_leaf_29_wb_clk_i _0290_ net233 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7581_ _0420_ team_08_WB.instance_to_wrap.allocation.game.game.score\[1\] net255
+ _2368_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6532_ _2453_ _2454_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[13\]
+ sky130_fd_sc_hd__nor2_1
X_9251_ clknet_leaf_15_wb_clk_i _0102_ net213 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6463_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[18\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[17\]
+ _2405_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[19\]
+ vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__or4b_1
XFILLER_0_43_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5414_ _0852_ _1215_ _1366_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__a21bo_2
X_9182_ clknet_leaf_11_wb_clk_i _0045_ net226 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_8202_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[4\]
+ _2984_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[5\]
+ vssd1 vssd1 vccd1 vccd1 _3715_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8133_ _0642_ _2386_ net279 vssd1 vssd1 vccd1 vccd1 _3659_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6394_ team_08_WB.instance_to_wrap.allocation.game.game.score\[4\] _2328_ team_08_WB.instance_to_wrap.allocation.game.game.score\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__a21oi_1
X_5345_ net129 _1244_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__or2_1
XANTENNA__5751__A _1012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5276_ _1205_ _1207_ net123 vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_54_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8064_ _0703_ _3595_ vssd1 vssd1 vccd1 vccd1 _3596_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_71_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7015_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[5\] team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[4\] vssd1 vssd1
+ vccd1 vccd1 _2771_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_71_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8966_ net98 _3276_ _4088_ net100 vssd1 vssd1 vccd1 vccd1 _4443_ sky130_fd_sc_hd__a31o_1
X_7917_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] team_08_WB.instance_to_wrap.allocation.game.controller.v\[2\]
+ _3458_ vssd1 vssd1 vccd1 vccd1 _3459_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5198__A _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8897_ net190 _2267_ _4373_ _2264_ _3284_ vssd1 vssd1 vccd1 vccd1 _4374_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7848_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[5\] _3408_
+ vssd1 vssd1 vccd1 vccd1 _3413_ sky130_fd_sc_hd__and3_1
XANTENNA__8005__C net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5736__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7779_ net292 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] net290 vssd1
+ vssd1 vccd1 vccd1 _3368_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8135__C1 _3597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9518_ net393 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_78_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8047__A_N team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9449_ clknet_leaf_45_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[3\]
+ net238 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_61_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7352__S _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8972__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9583__447 vssd1 vssd1 vccd1 vccd1 _9583__447/HI net447 sky130_fd_sc_hd__conb_1
XFILLER_0_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7527__S team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8212__A _3034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4740__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput35 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
Xinput24 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9477__352 vssd1 vssd1 vccd1 vccd1 _9477__352/HI net352 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_70_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6667__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7770__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5130_ _1081_ _1082_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9518__393 vssd1 vssd1 vccd1 vccd1 _9518__393/HI net393 sky130_fd_sc_hd__conb_1
X_5061_ _1012_ _1013_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__and2_2
XFILLER_0_35_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8882__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8820_ _4294_ _4297_ _4295_ vssd1 vssd1 vccd1 vccd1 _4298_ sky130_fd_sc_hd__a21oi_1
X_5963_ _0918_ _1813_ _1812_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__a21o_1
X_8751_ _4226_ _4228_ vssd1 vssd1 vccd1 vccd1 _4229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4914_ _0787_ _0793_ _0788_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__a21bo_4
XTAP_TAPCELL_ROW_36_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7702_ net126 net117 vssd1 vssd1 vccd1 vccd1 _3292_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5894_ _0773_ _0931_ _1846_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8682_ _4119_ _4158_ _4160_ net150 vssd1 vssd1 vccd1 vccd1 _4161_ sky130_fd_sc_hd__a22oi_1
X_4845_ net168 _0756_ _0762_ _0763_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__6915__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7633_ _3210_ _3222_ vssd1 vssd1 vccd1 vccd1 _3223_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9367__RESET_B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7564_ net257 _3168_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__or2_1
X_4776_ _0625_ _0727_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_56_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8117__C1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5465__B _1417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout227_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9303_ clknet_leaf_13_wb_clk_i net336 net214 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_6515_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[8\] _2441_
+ vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7495_ net304 _3071_ _3092_ _3050_ net302 vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__o221a_1
X_9234_ clknet_leaf_21_wb_clk_i _0062_ net241 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6446_ net296 _2392_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__and2_2
XFILLER_0_101_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9165_ _0140_ _0415_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_12_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6377_ team_08_WB.instance_to_wrap.allocation.game.game.score\[3\] _2327_ vssd1 vssd1
+ vccd1 vccd1 _2328_ sky130_fd_sc_hd__and2_1
X_5328_ _1227_ _1278_ _1280_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__or3_1
X_8116_ _0687_ _3614_ vssd1 vssd1 vccd1 vccd1 _3643_ sky130_fd_sc_hd__or2_1
X_9096_ clknet_leaf_52_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[26\]
+ net209 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4809__B _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8047_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] net318 vssd1
+ vssd1 vccd1 vccd1 _3582_ sky130_fd_sc_hd__nand2b_1
X_5259_ _1163_ _1211_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8949_ net177 _3707_ _4425_ vssd1 vssd1 vccd1 vccd1 _4426_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5656__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7871__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8967__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6487__A _2423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7590__B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__7589__Y _3179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[2\]
+ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4630_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[1\] vssd1
+ vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6300_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[17\]
+ _2199_ _2201_ _2252_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4561_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[15\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[14\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[16\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[17\]
+ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_42_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8114__A2 _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4492_ net624 vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__inv_2
X_7280_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[18\]
+ _2958_ vssd1 vssd1 vccd1 vccd1 _2960_ sky130_fd_sc_hd__and2_1
XANTENNA__6668__Y _2544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6231_ _1347_ _1348_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__and2b_1
XANTENNA__4583__A_N team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _2113_ _2114_ _2070_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _1036_ _1065_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6093_ _1882_ _2045_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5044_ _0967_ _0975_ _0976_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8803_ _3313_ _3888_ _3870_ vssd1 vssd1 vccd1 vccd1 _4281_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout177_A _3178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6995_ _2758_ vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5946_ _1895_ _1898_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8734_ net326 _3763_ vssd1 vssd1 vccd1 vccd1 _4212_ sky130_fd_sc_hd__nand2_1
X_5877_ _1826_ _1827_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_66_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8665_ net119 _3608_ vssd1 vssd1 vccd1 vccd1 _4144_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4828_ _0776_ _0780_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__and2b_2
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7616_ _3190_ _3205_ vssd1 vssd1 vccd1 vccd1 _3206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7561__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6364__A1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8596_ _0432_ _0658_ vssd1 vssd1 vccd1 vccd1 _4075_ sky130_fd_sc_hd__or2_1
X_7547_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr1\[1\] team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr1\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.clk1 vssd1
+ vssd1 vccd1 vccd1 _3159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4759_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.state\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.state\[0\] vssd1
+ vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7691__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7478_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\] _3113_
+ _3115_ _3118_ _3022_ vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__a41o_1
X_9217_ clknet_leaf_18_wb_clk_i _0074_ net229 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6429_ _2358_ _2377_ _2351_ _2354_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__a211oi_1
Xclkbuf_leaf_12_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9148_ clknet_leaf_41_wb_clk_i _0249_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__8408__A3 _3888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9079_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[9\]
+ net223 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8041__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9289__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8329__C1 _3635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8344__A2 _2393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8895__A3 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8697__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9589__453 vssd1 vssd1 vccd1 vccd1 _9589__453/HI net453 sky130_fd_sc_hd__conb_1
Xhold2 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.tft_reset vssd1 vssd1
+ vccd1 vccd1 net500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8032__A1 _0505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5800_ _1744_ _1751_ _1752_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__a21oi_2
X_6780_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[6\]
+ _2619_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5731_ _1682_ _1683_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5662_ _1565_ _1566_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__xnor2_1
XANTENNA__6346__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8450_ _3916_ _3930_ _3859_ vssd1 vssd1 vccd1 vccd1 _3931_ sky130_fd_sc_hd__a21oi_2
X_5593_ net131 _1489_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4613_ _0540_ _0571_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__nand2_1
X_8381_ net135 net124 _3861_ vssd1 vssd1 vccd1 vccd1 _3862_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7401_ net307 net309 vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_13_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7332_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[22\]
+ _2999_ vssd1 vssd1 vccd1 vccd1 _3000_ sky130_fd_sc_hd__nor2_1
X_4544_ _0506_ _0507_ _0512_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__nor3_1
XANTENNA__5743__B _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7263_ net566 _2946_ _2948_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4475_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__inv_2
X_6214_ _1011_ _1014_ _1056_ _1058_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__a31oi_1
X_9002_ clknet_leaf_4_wb_clk_i _0166_ net205 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_7194_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[13\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[14\]
+ _2896_ vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6145_ _0724_ _0917_ _2097_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__or3b_1
XFILLER_0_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6076_ _2025_ _2028_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__nand2_1
X_5027_ _0892_ _0894_ _0978_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_68_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8023__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6978_ _2747_ _2417_ _2746_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__and3b_1
X_8717_ _4089_ _4132_ _4174_ _4195_ _4087_ vssd1 vssd1 vccd1 vccd1 _4196_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_24_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5929_ net182 _0905_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9311__RESET_B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8648_ _2536_ _4116_ _4126_ vssd1 vssd1 vccd1 vccd1 _4127_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8579_ _4046_ _4047_ _4049_ _4042_ vssd1 vssd1 vccd1 vccd1 _4058_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6765__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5076__B2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8980__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4587__B1 _0552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8317__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6005__A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6659__B _2532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5303__A2 _1047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4511__A0 team_08_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8253__A1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4907__B _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8253__B2 _0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7950_ _0421_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[1\] vssd1
+ vssd1 vccd1 vccd1 _3490_ sky130_fd_sc_hd__nand2_1
X_7881_ _3435_ _3436_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[14\]
+ net166 vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__a2bb2o_1
X_6901_ net622 _2698_ net267 vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__o21ai_1
X_9620_ net481 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XANTENNA__4923__A _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6832_ _2653_ _2654_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9551_ net419 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6763_ _2606_ _2608_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_100_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5714_ _0936_ _1666_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__xor2_1
X_9482_ net357 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
X_6694_ net272 _2561_ _2562_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__nor3_1
XFILLER_0_57_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8502_ _3308_ _3360_ _3980_ net173 vssd1 vssd1 vccd1 vccd1 _3982_ sky130_fd_sc_hd__o211a_1
X_5645_ _1575_ _1577_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8433_ net149 net124 _3913_ vssd1 vssd1 vccd1 vccd1 _3914_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5576_ _1527_ _1528_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8364_ _3471_ _3849_ _3842_ vssd1 vssd1 vccd1 vccd1 _3850_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6569__B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8295_ _3522_ _3772_ _3786_ _3787_ net193 vssd1 vssd1 vccd1 vccd1 _3788_ sky130_fd_sc_hd__o311a_1
X_4527_ net329 team_08_WB.instance_to_wrap.allocation.game.controller.v\[2\] _0495_
+ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7315_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[2\]
+ _2982_ vssd1 vssd1 vccd1 vccd1 _2983_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4458_ net299 vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__inv_2
X_7246_ net179 _2935_ _2937_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__and3_1
X_7177_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[8\] _2887_ net164
+ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__a21oi_1
X_6128_ _2066_ _2067_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6059_ _1970_ _2010_ _2009_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_29_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5929__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8024__B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4552__B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8975__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5839__A _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8869__B _3542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7773__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5430_ _1335_ _1382_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8171__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5361_ _1263_ _1313_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5292_ net129 _1244_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__nand2_1
X_7100_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[22\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[23\]
+ _2837_ _2838_ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_39_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8080_ _0660_ _0664_ vssd1 vssd1 vccd1 vccd1 _3610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7031_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\] vssd1
+ vssd1 vccd1 vccd1 _2780_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_87_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8982_ net312 vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7933_ team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[1\] _2426_ net277
+ vssd1 vssd1 vccd1 vccd1 _3474_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5460__A1 _1217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7864_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[9\]
+ _3421_ net159 vssd1 vssd1 vccd1 vccd1 _3425_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout257_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6672__B1_N _2544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9603_ net467 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
X_6815_ _2642_ _2643_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7795_ _2398_ _3378_ _3380_ _2375_ vssd1 vssd1 vccd1 vccd1 _3381_ sky130_fd_sc_hd__a211oi_1
X_6746_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[9\]
+ _2596_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9534_ net490 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_18_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6677_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[9\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__or4_1
X_9465_ net340 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
X_5628_ _1580_ _1572_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__and2b_1
X_9396_ clknet_leaf_31_wb_clk_i _0343_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8416_ _3290_ _3879_ _3297_ vssd1 vssd1 vccd1 vccd1 _3897_ sky130_fd_sc_hd__o21ai_1
X_9494__369 vssd1 vssd1 vccd1 vccd1 _9494__369/HI net369 sky130_fd_sc_hd__conb_1
X_5559_ _1509_ _1510_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8347_ _3460_ _3580_ _3835_ _3836_ vssd1 vssd1 vccd1 vccd1 _3837_ sky130_fd_sc_hd__o22a_1
XFILLER_0_41_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4680__C_N team_08_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8278_ _3492_ _3760_ _3520_ vssd1 vssd1 vccd1 vccd1 _3772_ sky130_fd_sc_hd__a21oi_1
X_7229_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[0\]
+ _2922_ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7976__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8940__A2 _3276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output53_A net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7768__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4930_ _0785_ _0846_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4861_ _0810_ _0812_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8931__A2 _3329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6600_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[12\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[13\]
+ _2497_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[14\] vssd1
+ vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__a31o_1
X_4792_ net168 _0743_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__nand2_4
XFILLER_0_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7580_ net290 net692 _3176_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8144__B1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6531_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[13\] _2451_
+ net156 vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9250_ clknet_leaf_15_wb_clk_i _0101_ net214 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6462_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[21\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[20\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[22\]
+ vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__or3b_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8695__A1 _4001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8695__B2 _4036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5413_ _1217_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9181_ clknet_leaf_11_wb_clk_i _0044_ net226 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8201_ _2985_ _3714_ _3713_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6393_ _2341_ _2342_ team_08_WB.instance_to_wrap.allocation.game.game.score\[6\]
+ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__mux2_1
X_5344_ net129 _1296_ _1294_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8132_ _0646_ _2323_ vssd1 vssd1 vccd1 vccd1 _3658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5275_ _0915_ _1227_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8063_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\] _0656_
+ vssd1 vssd1 vccd1 vccd1 _3595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7014_ _0453_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[4\]
+ _2770_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[2\] vssd1
+ vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__a211o_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7958__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8965_ _4406_ _4408_ _4441_ vssd1 vssd1 vccd1 vccd1 _4442_ sky130_fd_sc_hd__a21oi_1
X_7916_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\]
+ net289 team_08_WB.instance_to_wrap.allocation.game.controller.v\[7\] vssd1 vssd1
+ vccd1 vccd1 _3458_ sky130_fd_sc_hd__or4_2
X_8896_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ _0450_ _0451_ net192 vssd1 vssd1 vccd1 vccd1 _4373_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_37_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_7847_ net159 _3411_ _3412_ net165 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7694__A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8922__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7778_ net292 net291 net207 _3367_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4830__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6729_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[3\]
+ _2585_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__and2_1
X_9517_ net392 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_78_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9448_ clknet_leaf_42_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[2\]
+ net238 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__8686__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9379_ clknet_leaf_32_wb_clk_i _0326_ net245 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5006__X _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4845__X _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6773__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6621__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput36 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5060_ net143 _0836_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5962_ _1880_ _1914_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__nor2_1
XANTENNA__5299__A _1039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8750_ net333 net192 vssd1 vssd1 vccd1 vccd1 _4228_ sky130_fd_sc_hd__xor2_1
X_4913_ _0862_ _0865_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_36_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7701_ net124 net116 vssd1 vssd1 vccd1 vccd1 _3291_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5893_ _0761_ _0929_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__nor2_1
X_8681_ _4158_ _4159_ vssd1 vssd1 vccd1 vccd1 _4160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4844_ _0774_ _0795_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7632_ _3206_ _3207_ _3209_ net126 vssd1 vssd1 vccd1 vccd1 _3222_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__8403__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7563_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr2\[1\] team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr2\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.clk1 vssd1
+ vssd1 vccd1 vccd1 _3168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4775_ _0621_ _0626_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9302_ clknet_leaf_13_wb_clk_i _0122_ net214 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_6514_ _2441_ _2442_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9233_ clknet_2_3__leaf_wb_clk_i _0061_ net241 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_7494_ _3025_ _3043_ vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_67_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6445_ net280 _2391_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9164_ _0139_ _0414_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_6376_ team_08_WB.instance_to_wrap.allocation.game.game.score\[2\] team_08_WB.instance_to_wrap.allocation.game.game.score\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.game.score\[1\] vssd1 vssd1 vccd1 vccd1
+ _2327_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5327_ _1256_ _1261_ _1259_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_73_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8115_ _0688_ _3641_ vssd1 vssd1 vccd1 vccd1 _3642_ sky130_fd_sc_hd__nor2_1
X_9095_ clknet_leaf_52_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[25\]
+ net209 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_8046_ _3564_ _3580_ vssd1 vssd1 vccd1 vccd1 _3581_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8840__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5258_ _1148_ _1162_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7689__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5189_ _1140_ _1141_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4825__B net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8948_ _4422_ _4423_ _4424_ vssd1 vssd1 vccd1 vccd1 _4425_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4614__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5937__A _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8879_ _4345_ _4346_ _4354_ _4356_ vssd1 vssd1 vccd1 vccd1 _4357_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9240__SET_B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8967__B net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9077__RESET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8983__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 net181 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_2
XFILLER_0_89_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4735__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6070__A1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6008__A _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5847__A _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8898__B2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8898__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4560_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[7\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[9\]
+ _0527_ _0528_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4491_ net300 vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6230_ _1302_ _2146_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _2068_ _2069_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8893__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _1063_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__nand2_1
XANTENNA__7086__B1 _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6092_ _2033_ _2044_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8822__A1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5043_ _0956_ _0957_ _0989_ _0987_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__a31o_1
XANTENNA__4926__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6833__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8802_ net97 _4266_ _4278_ _4264_ _4277_ vssd1 vssd1 vccd1 vccd1 _4280_ sky130_fd_sc_hd__a221o_1
X_6994_ _0468_ _2756_ vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5945_ _1895_ _1896_ _1897_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__nand3_1
X_8733_ net104 _4208_ _4210_ _4207_ vssd1 vssd1 vccd1 vccd1 _4211_ sky130_fd_sc_hd__a211o_1
X_5876_ _0918_ _1721_ _1719_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5757__A _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8664_ net119 _3608_ vssd1 vssd1 vccd1 vccd1 _4143_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4827_ _0599_ _0601_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7615_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[10\]
+ _3191_ net133 vssd1 vssd1 vccd1 vccd1 _3205_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8595_ net134 _4071_ _4073_ _4065_ vssd1 vssd1 vccd1 vccd1 _4074_ sky130_fd_sc_hd__o211a_1
X_7546_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr1\[0\] net551
+ _3158_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__o21ai_1
X_4758_ team_08_WB.instance_to_wrap.allocation.game.controller.block_done net139 _0712_
+ team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\] vssd1 vssd1 vccd1
+ vccd1 _0005_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout125_X net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5492__A _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4689_ net288 _0643_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__or2_1
X_7477_ net304 _3041_ _3052_ _3117_ vssd1 vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7691__B net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9216_ clknet_leaf_17_wb_clk_i _0073_ net229 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6428_ _2377_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9147_ clknet_leaf_41_wb_clk_i _0248_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6359_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9078_ clknet_leaf_49_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[8\]
+ net224 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_8029_ net194 _3563_ _3564_ vssd1 vssd1 vccd1 vccd1 _3565_ sky130_fd_sc_hd__and3_1
XANTENNA__7092__A3 _2832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__7212__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8329__B1 _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8978__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4746__A team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[0\]
+ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9110__Q team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5730_ _1599_ _1627_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5661_ _1140_ _1600_ _1613_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7400_ net307 net308 vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__or2_1
X_5592_ net132 _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_61_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4612_ _0569_ _0570_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__xnor2_1
X_8380_ net112 _3860_ vssd1 vssd1 vccd1 vccd1 _3861_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9449__SET_B net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7331_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[21\]
+ _2998_ vssd1 vssd1 vccd1 vccd1 _2999_ sky130_fd_sc_hd__or2_1
X_4543_ _0508_ _0509_ _0510_ _0511_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8400__B net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7262_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[12\]
+ _2946_ net179 vssd1 vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4474_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__inv_2
X_6213_ _1038_ _1042_ _2165_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__a21o_1
X_9001_ clknet_leaf_4_wb_clk_i _0165_ net203 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7193_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[13\] _2896_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[14\]
+ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6144_ _2084_ _2096_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__and2_1
X_6075_ _2025_ _2026_ _2027_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__nand3_1
X_5026_ _0892_ _0894_ _0978_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5085__A2 _0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[20\]
+ _2744_ vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5928_ _1866_ _1867_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout242_X net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8716_ net279 _2386_ _4184_ _4194_ vssd1 vssd1 vccd1 vccd1 _4195_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5859_ _1810_ _1811_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8647_ net149 _4119_ _4121_ _4125_ _4118_ vssd1 vssd1 vccd1 vccd1 _4126_ sky130_fd_sc_hd__o311a_1
X_9620__481 vssd1 vssd1 vccd1 vccd1 _9620__481/HI net481 sky130_fd_sc_hd__conb_1
XANTENNA__5545__B1 _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9351__RESET_B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8578_ _3241_ _3596_ _4002_ _4005_ _4053_ vssd1 vssd1 vccd1 vccd1 _4057_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7529_ net532 net502 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5076__A2 _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4587__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9092__RESET_B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8501__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9021__RESET_B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6659__C _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4747__Y _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7880_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[14\]
+ _3433_ _3403_ vssd1 vssd1 vccd1 vccd1 _3436_ sky130_fd_sc_hd__o21ai_1
X_6900_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[4\]
+ _2697_ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6831_ net602 _2652_ net271 vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4923__B _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9550_ net418 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XANTENNA__7764__A1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5100__A _1012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6762_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ _2605_ _2607_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_63_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8501_ net173 _3980_ vssd1 vssd1 vccd1 vccd1 _3981_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9481_ net356 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5713_ _0813_ _0932_ _1665_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__or3_1
XFILLER_0_73_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6693_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[4\]
+ _2558_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5644_ _1553_ _1582_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8432_ net149 net135 _3314_ _3895_ vssd1 vssd1 vccd1 vccd1 _3913_ sky130_fd_sc_hd__or4b_1
X_8363_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] _3470_ vssd1
+ vssd1 vccd1 vccd1 _3849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5575_ _1500_ _1526_ vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7314_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__or2_1
X_8294_ _3522_ _3772_ _3786_ vssd1 vssd1 vccd1 vccd1 _3787_ sky130_fd_sc_hd__o21ai_1
X_4526_ _0489_ _0492_ _0494_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout202_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4457_ net4 vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__inv_2
X_7245_ _2936_ vssd1 vssd1 vccd1 vccd1 _2937_ sky130_fd_sc_hd__inv_2
X_7176_ _2874_ _2887_ _2888_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input7_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6127_ _2079_ _2078_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout192_X net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6058_ _1970_ _2009_ _2010_ vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_29_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ _0819_ _0960_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__and2b_1
XANTENNA__7697__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5929__B _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8180__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5839__B _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4743__B _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5855__A _0814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5360_ _1251_ _1262_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5291_ _1241_ _1242_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__xnor2_1
XANTENNA__6686__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7030_ _0434_ _2778_ _2775_ vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_56_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4477__Y _0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7013__C team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8981_ net312 vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__inv_2
X_7932_ _3468_ net170 net297 vssd1 vssd1 vccd1 vccd1 _3473_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7863_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[9\]
+ _3421_ vssd1 vssd1 vccd1 vccd1 _3424_ sky130_fd_sc_hd__and2_1
XANTENNA__4653__B team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9602_ net466 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_92_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6814_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[3\]
+ _2641_ net271 vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__o21ai_1
X_7794_ _2358_ _3379_ vssd1 vssd1 vccd1 vccd1 _3380_ sky130_fd_sc_hd__xnor2_1
X_6745_ net272 _2595_ _2596_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__nor3_1
X_9533_ net489 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9464_ net339 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_46_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6676_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__or4b_1
XFILLER_0_45_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8162__A1 _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8162__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8415_ _3289_ _3303_ _3895_ _3295_ _3297_ vssd1 vssd1 vccd1 vccd1 _3896_ sky130_fd_sc_hd__o221a_1
X_5627_ _1573_ _1578_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__xnor2_1
X_9395_ clknet_leaf_31_wb_clk_i _0342_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5558_ _0814_ _0906_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__nand2_1
X_8346_ _0570_ _3582_ _3822_ net197 vssd1 vssd1 vccd1 vccd1 _3836_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4509_ net266 vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8277_ net139 _2271_ vssd1 vssd1 vccd1 vccd1 _3771_ sky130_fd_sc_hd__nor2_1
X_5489_ _1440_ _1441_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_76_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7228_ _2924_ _2925_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__nor2_1
XANTENNA__4828__B _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7159_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[0\] net261 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2878_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7976__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8986__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7967__A1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4754__A _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5442__A2 _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4860_ _0809_ _0811_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__nor2_4
XFILLER_0_75_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4791_ _0718_ _0742_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__nand2_2
X_6530_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[13\] _2451_
+ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__and2_1
XANTENNA__8144__A1 _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6461_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[6\]
+ _2403_ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5412_ _0852_ _1215_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9180_ clknet_leaf_17_wb_clk_i _0043_ net227 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_8200_ net557 _2984_ vssd1 vssd1 vccd1 vccd1 _3714_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6392_ team_08_WB.instance_to_wrap.allocation.game.game.score\[3\] _2338_ vssd1 vssd1
+ vccd1 vccd1 _2343_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5343_ _1294_ _1295_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8131_ _0428_ _0646_ net279 vssd1 vssd1 vccd1 vccd1 _3657_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5274_ _0940_ _1226_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_54_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8062_ _3593_ _3594_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[1\]
+ net237 vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__o2bb2a_1
X_7013_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[6\] team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\] team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_71_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8407__Y _3888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9195__RESET_B net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8964_ _4409_ _4417_ _4432_ _4440_ vssd1 vssd1 vccd1 vccd1 _4441_ sky130_fd_sc_hd__o211a_1
X_7915_ net335 _2426_ _3456_ vssd1 vssd1 vccd1 vccd1 _3457_ sky130_fd_sc_hd__a21o_1
X_8895_ _2279_ net96 net102 _4371_ net99 vssd1 vssd1 vccd1 vccd1 _4372_ sky130_fd_sc_hd__o32a_1
X_7846_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[4\]
+ _3408_ vssd1 vssd1 vccd1 vccd1 _3412_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout155_X net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7694__B team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4989_ net128 _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7777_ _3357_ _3362_ _3366_ _3350_ _3274_ vssd1 vssd1 vccd1 vccd1 _3367_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9516_ net391 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_73_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6728_ net272 _2584_ _2585_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9502__377 vssd1 vssd1 vccd1 vccd1 _9502__377/HI net377 sky130_fd_sc_hd__conb_1
X_9447_ clknet_leaf_12_wb_clk_i _0392_ net219 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6659_ net286 _2532_ _2536_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8686__A2 _3622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7894__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9378_ clknet_leaf_33_wb_clk_i _0325_ net247 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.wr
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8329_ _2294_ _2393_ _2426_ _3562_ _3635_ vssd1 vssd1 vccd1 vccd1 _3820_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4839__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5121__A1 _0919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7949__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput37 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
Xinput15 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5692__X _1645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5299__B _1047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5961_ _1881_ _1913_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__nand2_1
X_4912_ _0858_ _0864_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4771__X _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7700_ net149 net133 vssd1 vssd1 vccd1 vccd1 _3290_ sky130_fd_sc_hd__nand2_2
X_8680_ net286 net283 _0643_ net281 vssd1 vssd1 vccd1 vccd1 _4159_ sky130_fd_sc_hd__a31o_1
X_5892_ _1843_ _1844_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__nor2_1
XANTENNA__8365__A1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7631_ _3218_ _3220_ vssd1 vssd1 vccd1 vccd1 _3221_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4843_ _0795_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7562_ _3166_ _3167_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__nor2_1
X_4774_ _0624_ _0725_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__nor2_2
XFILLER_0_55_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9301_ clknet_leaf_13_wb_clk_i _0121_ net217 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6513_ net677 _2439_ _2429_ vssd1 vssd1 vccd1 vccd1 _2442_ sky130_fd_sc_hd__o21ai_1
X_7493_ _3109_ _3121_ _3132_ net114 net502 vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__o32a_1
XFILLER_0_71_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9232_ clknet_leaf_21_wb_clk_i _0060_ net241 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6444_ _2387_ _2388_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5351__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9163_ _0138_ _0413_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_6375_ team_08_WB.instance_to_wrap.allocation.game.game.score\[0\] team_08_WB.instance_to_wrap.allocation.game.game.score\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__and2_2
XFILLER_0_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5326_ _1227_ _1278_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8114_ _0675_ _0686_ net162 vssd1 vssd1 vccd1 vccd1 _3641_ sky130_fd_sc_hd__o21ba_1
X_9094_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[24\]
+ net209 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5257_ _1193_ _1209_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__nand2_1
X_8045_ net314 _3559_ vssd1 vssd1 vccd1 vccd1 _3580_ sky130_fd_sc_hd__xnor2_2
XANTENNA__9376__RESET_B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7689__B net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5188_ _0824_ _0839_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__xor2_2
XANTENNA__4862__B1 _0814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7041__Y _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9305__RESET_B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8947_ net177 _3707_ vssd1 vssd1 vccd1 vccd1 _4424_ sky130_fd_sc_hd__nor2_1
X_9543__411 vssd1 vssd1 vccd1 vccd1 _9543__411/HI net411 sky130_fd_sc_hd__conb_1
XFILLER_0_65_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7159__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8878_ _4281_ _4355_ vssd1 vssd1 vccd1 vccd1 _4356_ sky130_fd_sc_hd__nor2_1
X_7829_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\]
+ _3401_ _3400_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8967__C _3279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9630__483 vssd1 vssd1 vccd1 vccd1 _9630__483/HI net483 sky130_fd_sc_hd__conb_1
Xfanout170 _3472_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_4
Xfanout181 _2923_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__9046__RESET_B net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout192 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[1\]
+ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8595__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6070__A2 _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8347__A1 _3460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8504__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4490_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _2080_ _2081_ _2112_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__a21oi_1
X_5111_ _1061_ _1062_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__or2_1
XANTENNA__4766__X _0719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8893__B net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6694__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6091_ _2041_ _2042_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__xor2_1
XANTENNA__8822__A2 _0425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5042_ _0992_ _0994_ _0991_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5103__A _1047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8801_ net314 _3266_ vssd1 vssd1 vccd1 vccd1 _4279_ sky130_fd_sc_hd__or2_1
X_6993_ _0467_ _0468_ _2757_ _2754_ _2753_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__o32a_2
XTAP_TAPCELL_ROW_49_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5944_ _1849_ _1894_ _1893_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__a21o_1
X_8732_ _4209_ vssd1 vssd1 vccd1 vccd1 _4210_ sky130_fd_sc_hd__inv_2
XANTENNA__8414__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5875_ _1826_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__and2b_1
XANTENNA__5757__B _0926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4661__B team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8663_ net127 _3681_ vssd1 vssd1 vccd1 vccd1 _4142_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout232_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4826_ _0772_ _0774_ _0778_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7614_ _3202_ _3203_ vssd1 vssd1 vccd1 vccd1 _3204_ sky130_fd_sc_hd__and2b_1
X_8594_ net155 _4067_ _4068_ vssd1 vssd1 vccd1 vccd1 _4073_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7545_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr1\[0\] _3157_
+ net257 vssd1 vssd1 vccd1 vccd1 _3158_ sky130_fd_sc_hd__a21oi_1
XANTENNA__7972__B _3472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5572__A1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4757_ team_08_WB.instance_to_wrap.allocation.game.controller.block_done _0711_ vssd1
+ vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__nand2b_1
XANTENNA__8420__Y _3901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7313__A2 _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4688_ net286 _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__nor2_2
X_7476_ net307 _3041_ _3071_ _0440_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__o211a_1
XANTENNA__5492__B _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9215_ clknet_leaf_17_wb_clk_i _0072_ net229 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_6427_ _2368_ _2371_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6358_ _2308_ _2309_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_8_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9146_ clknet_leaf_37_wb_clk_i _0247_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_9614__478 vssd1 vssd1 vccd1 vccd1 _9614__478/HI net478 sky130_fd_sc_hd__conb_1
X_5309_ _1256_ _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7077__A1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6289_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[7\]
+ _2217_ _2220_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__a22o_1
XANTENNA__4676__X _0634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9077_ clknet_leaf_49_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[7\]
+ net224 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_8028_ net321 _3534_ _3561_ vssd1 vssd1 vccd1 vccd1 _3564_ sky130_fd_sc_hd__or3_1
X_9467__342 vssd1 vssd1 vccd1 vccd1 _9467__342/HI net342 sky130_fd_sc_hd__conb_1
XFILLER_0_98_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6588__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8324__A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5667__B net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9508__383 vssd1 vssd1 vccd1 vccd1 _9508__383/HI net383 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_27_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_49_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6779__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9227__RESET_B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7607__A3 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4826__A0 _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[5\] vssd1
+ vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5660_ _1611_ _1612_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ net313 team_08_WB.instance_to_wrap.allocation.game.controller.v\[7\] vssd1
+ vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__xnor2_4
XANTENNA__8740__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5593__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5591_ _1540_ _1542_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7330_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[20\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[19\]
+ _2996_ vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__or3_1
X_4542_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[14\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[17\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[16\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[15\]
+ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__or4b_1
X_4473_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7261_ _2946_ _2947_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6212_ _1039_ _1041_ _0861_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9000_ clknet_leaf_4_wb_clk_i _0164_ net203 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8256__A0 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7192_ net582 _2896_ _2898_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4937__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6143_ _2034_ _2083_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__or2_1
X_6074_ _1986_ _1997_ _2024_ vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__a21o_1
X_5025_ _0967_ _0977_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8008__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8559__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6976_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[20\]
+ _2744_ vssd1 vssd1 vccd1 vccd1 _2746_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5927_ _1865_ _1869_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8715_ _4190_ _4192_ _4193_ vssd1 vssd1 vccd1 vccd1 _4194_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5858_ _0923_ _1762_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8731__B2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8646_ _4120_ _4122_ _4123_ net153 _4124_ vssd1 vssd1 vccd1 vccd1 _4125_ sky130_fd_sc_hd__o221a_1
X_5789_ _1739_ _1740_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__xor2_1
X_4809_ net144 _0761_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__or2_4
XFILLER_0_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8577_ _0695_ _4043_ _0694_ vssd1 vssd1 vccd1 vccd1 _4056_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7528_ net537 net521 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__mux2_1
X_7459_ net309 _3091_ _3100_ vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9129_ clknet_leaf_37_wb_clk_i _0230_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__8798__A1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7997__C1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6830_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[9\]
+ _2652_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6761_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_63_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5712_ _0809_ _0930_ _0928_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5100__B _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8500_ net153 net133 _3291_ _3895_ _3364_ vssd1 vssd1 vccd1 vccd1 _3980_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_100_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6692_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[4\]
+ _2558_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9480_ net355 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_100_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5643_ _1591_ _1593_ _1595_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8431_ _3312_ _3909_ _3910_ _3911_ vssd1 vssd1 vccd1 vccd1 _3912_ sky130_fd_sc_hd__a22o_1
X_5574_ _1500_ _1526_ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8362_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[2\] _2875_ _3848_
+ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__a21o_1
XANTENNA__7308__A _2972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4525_ net329 team_08_WB.instance_to_wrap.allocation.game.controller.v\[2\] vssd1
+ vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__xnor2_2
X_7313_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[5\] _2975_ _2977_
+ _2980_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8293_ _0485_ _3530_ _3785_ vssd1 vssd1 vccd1 vccd1 _3786_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4456_ net293 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7244_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[5\]
+ _2932_ vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7175_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[6\] _2885_ net687
+ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__a21oi_1
X_6126_ _1882_ _2045_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6057_ _1967_ _1969_ _1968_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5008_ _0960_ _0819_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_29_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7697__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6959_ _0462_ _2734_ vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4569__A2 _0505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9579__443 vssd1 vssd1 vccd1 vccd1 _9579__443/HI net443 sky130_fd_sc_hd__conb_1
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8629_ _4090_ _4091_ _4104_ _4107_ vssd1 vssd1 vccd1 vccd1 _4108_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout98_X net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_X clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5855__B _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6706__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5290_ _1236_ _1240_ _1242_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__a21o_1
XANTENNA__5196__A_N _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8980_ net311 vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__inv_2
X_7931_ _0522_ _3458_ _3471_ vssd1 vssd1 vccd1 vccd1 _3472_ sky130_fd_sc_hd__nor3_4
X_9601_ net465 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7862_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[8\]
+ net165 net159 _3423_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__a22o_1
XANTENNA__8934__B2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6813_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[3\]
+ _2641_ vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7793_ _2364_ _2372_ vssd1 vssd1 vccd1 vccd1 _3379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6744_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[8\]
+ _2592_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__and3_1
X_9532_ net407 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XFILLER_0_19_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6675_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9463_ net338 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
X_5626_ _1573_ _1578_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8414_ net110 _3865_ vssd1 vssd1 vccd1 vccd1 _3895_ sky130_fd_sc_hd__nor2_2
X_9394_ clknet_leaf_30_wb_clk_i _0341_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_5557_ net142 _0909_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__nand2_1
X_8345_ _3582_ _3822_ _0570_ vssd1 vssd1 vccd1 vccd1 _3835_ sky130_fd_sc_hd__a21oi_1
X_4508_ _0473_ _0474_ _0475_ _0478_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__or4_1
X_5488_ _1435_ _1438_ _1439_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__and3_1
X_8276_ _3479_ _3757_ _3770_ net235 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout100_X net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7227_ net614 _2922_ net180 vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__o21ai_1
X_7158_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[1\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[0\]
+ net261 vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6109_ _2021_ _2061_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__xor2_1
X_7089_ _2829_ _2830_ _2779_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__o21a_1
XANTENNA__8083__D1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7976__A2 _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4860__A _0809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8332__A _0505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7593__D net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6787__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8456__A3 _3888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9560__428 vssd1 vssd1 vccd1 vccd1 _9560__428/HI net428 sky130_fd_sc_hd__conb_1
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4790_ _0718_ _0742_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__and2_4
XFILLER_0_68_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8242__A _3034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8144__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6460_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[5\]
+ _2401_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__and3_1
XANTENNA__7352__A0 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5411_ _0959_ _1222_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6391_ _2334_ _2340_ vssd1 vssd1 vccd1 vccd1 _2342_ sky130_fd_sc_hd__or2_1
X_5342_ _1290_ _1292_ _1293_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_58_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8130_ _0696_ _3645_ _3655_ vssd1 vssd1 vccd1 vccd1 _3656_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8061_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\] net137
+ _0654_ net237 vssd1 vssd1 vccd1 vccd1 _3594_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5273_ _0914_ _1223_ _1225_ _0915_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_54_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7012_ _0460_ _2769_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[1\]
+ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_71_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7958__A2 _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9569__497 vssd1 vssd1 vccd1 vccd1 net497 _9569__497/LO sky130_fd_sc_hd__conb_1
XANTENNA__4664__B team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8963_ _2293_ net99 _4124_ _4439_ vssd1 vssd1 vccd1 vccd1 _4440_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7914_ net299 team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\] _3455_
+ vssd1 vssd1 vccd1 vccd1 _3456_ sky130_fd_sc_hd__or3_2
XFILLER_0_37_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8894_ _2280_ net102 vssd1 vssd1 vccd1 vccd1 _4371_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout262_A _0514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7845_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[4\]
+ _3408_ vssd1 vssd1 vccd1 vccd1 _3411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4988_ _0818_ _0912_ _0915_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__a21oi_1
X_9515_ net390 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XANTENNA_fanout148_X net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7776_ _3335_ _3363_ _3365_ net175 vssd1 vssd1 vccd1 vccd1 _3366_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6727_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__and3_1
XANTENNA__7991__A team_08_WB.instance_to_wrap.allocation.game.controller.v\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9446_ clknet_leaf_12_wb_clk_i _0391_ net219 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6658_ net286 _2536_ vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__or2_1
XANTENNA__7894__A1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5609_ _0792_ _0906_ _1560_ _1558_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__a31o_1
X_9377_ clknet_leaf_32_wb_clk_i _0402_ net247 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.init_done
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_46_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8328_ net198 _3814_ _3818_ _3540_ vssd1 vssd1 vccd1 vccd1 _3819_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6589_ _2493_ _2494_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8259_ net300 _3752_ _3754_ _3474_ vssd1 vssd1 vccd1 vccd1 _3755_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_79_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_2
XANTENNA__8327__A _3460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4861__Y _0814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6909__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5686__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7582__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput16 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xinput38 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6310__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8062__B2 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9484__359 vssd1 vssd1 vccd1 vccd1 _9484__359/HI net359 sky130_fd_sc_hd__conb_1
X_5960_ _1910_ _1912_ _1908_ _1909_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__a2bb2o_1
X_4911_ _0851_ _0855_ _0857_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__and3_1
X_5891_ _1790_ _1796_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__xnor2_2
XANTENNA_clkbuf_2_0__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8365__A2 _2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7630_ _3191_ _3219_ vssd1 vssd1 vccd1 vccd1 _3220_ sky130_fd_sc_hd__xor2_1
X_4842_ net167 _0756_ _0762_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__mux2_2
XANTENNA__7573__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7561_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.clk1
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr2\[0\] team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr2\[1\]
+ net258 vssd1 vssd1 vccd1 vccd1 _3167_ sky130_fd_sc_hd__a31o_1
X_4773_ _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9300_ clknet_leaf_13_wb_clk_i _0120_ net217 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6512_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[7\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[6\]
+ _2437_ vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__and3_1
X_7492_ _3023_ _3131_ vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9231_ clknet_leaf_21_wb_clk_i _0059_ net241 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6443_ _0649_ _2385_ vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkload47_A clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout108_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9162_ _0137_ _0133_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_6374_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.state\[0\] _0420_
+ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__nor2_4
X_5325_ _0940_ _1226_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_73_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8113_ _3629_ _3637_ _3640_ net244 net592 vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__o32a_1
X_9093_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[23\]
+ net209 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_5256_ _1207_ _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8044_ _3481_ _3570_ _3579_ net241 net567 vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_3_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5187_ _0749_ _1139_ _0745_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4614__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7986__A _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8946_ net127 _3678_ vssd1 vssd1 vccd1 vccd1 _4423_ sky130_fd_sc_hd__nor2_1
XANTENNA__7800__B2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7800__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9345__RESET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8877_ net318 _3542_ _4279_ _4283_ _3931_ vssd1 vssd1 vccd1 vccd1 _4355_ sky130_fd_sc_hd__a311o_1
XFILLER_0_4_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7828_ _2781_ _3397_ vssd1 vssd1 vccd1 vccd1 _3401_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7759_ _3342_ _3346_ _3348_ _3326_ vssd1 vssd1 vccd1 vccd1 _3349_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_85_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8610__A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9429_ clknet_leaf_39_wb_clk_i _0374_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input38_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4856__Y _0809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 _0716_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_4
Xfanout160 _3403_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_4
Xfanout171 net172 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout193 net195 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4872__X _0825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4605__A1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5110_ _1061_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__nand2_1
X_6090_ _2041_ _2042_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__nor2_1
XANTENNA__7086__A2 _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8893__C _4370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5041_ _0991_ _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4495__A team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9566__434 vssd1 vssd1 vccd1 vccd1 _9566__434/HI net434 sky130_fd_sc_hd__conb_1
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
X_8800_ net314 net99 vssd1 vssd1 vccd1 vccd1 _4278_ sky130_fd_sc_hd__nor2_2
X_6992_ _2755_ _2756_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8731_ net103 _4205_ _4208_ net104 vssd1 vssd1 vccd1 vccd1 _4209_ sky130_fd_sc_hd__o2bb2a_1
X_5943_ net142 _0922_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5874_ _1772_ _1777_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8662_ _4137_ _4140_ vssd1 vssd1 vccd1 vccd1 _4141_ sky130_fd_sc_hd__nand2_1
X_4825_ _0738_ net148 vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__nand2_4
X_7613_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[10\]
+ net133 vssd1 vssd1 vccd1 vccd1 _3203_ sky130_fd_sc_hd__or2_1
X_8593_ net125 _4070_ _4071_ net134 vssd1 vssd1 vccd1 vccd1 _4072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7544_ net550 team_08_WB.instance_to_wrap.allocation.game.cactus1size.lfsr1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout225_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4756_ _0706_ _0710_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4687_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\] _0642_ vssd1
+ vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__or2_2
X_7475_ _0439_ net304 vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9573__438 vssd1 vssd1 vccd1 vccd1 _9573__438/HI net438 sky130_fd_sc_hd__conb_1
X_9214_ clknet_leaf_17_wb_clk_i _0071_ net231 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6426_ _2358_ _2372_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6357_ net331 _2306_ _2307_ net327 vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_8_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9145_ clknet_leaf_37_wb_clk_i net512 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5308_ _1259_ _1260_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__nor2_1
XANTENNA__7077__A2 _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6288_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[6\]
+ _2220_ _2222_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__o22ai_1
XANTENNA__7052__Y _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9076_ clknet_leaf_49_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[6\]
+ net224 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_5239_ net143 _1144_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__or2_1
X_8027_ net321 _3534_ _3561_ vssd1 vssd1 vccd1 vccd1 _3563_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8329__A2 _2393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8929_ _2278_ _3265_ vssd1 vssd1 vccd1 vccd1 _4406_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9209__Q team_08_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8576__A_N _3261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6795__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4586__Y _0552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8804__A3 _3888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5204__A _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[23\]
+ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8515__A team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4610_ net316 team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] _0536_
+ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8740__A2 _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5590_ _1540_ _1542_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8250__A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4541_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[19\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[20\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[18\] vssd1 vssd1
+ vccd1 vccd1 _0510_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_13_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4472_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__inv_2
X_7260_ net651 _2944_ net179 vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6211_ net129 _2163_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7191_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[13\] _2896_ _0523_
+ vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__o21ai_1
X_6142_ _2092_ _2093_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6073_ _1935_ _1937_ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__nand2_1
X_5024_ _0975_ _0976_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4953__A _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout175_A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6975_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[19\]
+ _2743_ _2745_ _2417_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__o211a_1
X_5926_ _1876_ _1877_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_85_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8714_ _4116_ _4183_ _4191_ vssd1 vssd1 vccd1 vccd1 _4193_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8645_ net279 net173 vssd1 vssd1 vccd1 vccd1 _4124_ sky130_fd_sc_hd__nand2_2
XFILLER_0_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5857_ _1808_ _1809_ _1806_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_63_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5788_ _1736_ _1738_ _1740_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__a21o_1
XANTENNA__5545__A2 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4808_ _0753_ _0759_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8576_ _3261_ _4053_ _4054_ _4004_ vssd1 vssd1 vccd1 vccd1 _4055_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_72_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7527_ net531 net517 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__mux2_1
X_4739_ net280 _0693_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__nand2_2
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7458_ net307 _0440_ _3043_ vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__or3_1
XANTENNA__8495__A1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6409_ _2344_ _2359_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__nor2_1
X_7389_ net650 _3036_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_101_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4847__B _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9128_ clknet_leaf_38_wb_clk_i _0229_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_9059_ clknet_leaf_34_wb_clk_i _0194_ net246 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8486__A1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9448__RESET_B net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6990__A_N team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6972__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6760_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[9\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__or4_1
X_5711_ _0936_ _1663_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6691_ net681 _2558_ _2560_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__o21a_1
XANTENNA__8174__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5642_ _1545_ _1594_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_80_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7921__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8430_ _3292_ _3307_ _3885_ vssd1 vssd1 vccd1 vccd1 _3911_ sky130_fd_sc_hd__or3_1
X_5573_ _0940_ _1473_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8361_ _3470_ _3847_ _3843_ vssd1 vssd1 vccd1 vccd1 _3848_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5109__A _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4524_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[2\] net329 vssd1
+ vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__nand2b_1
X_7312_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[4\] _2974_ _2979_
+ _2981_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__o211a_1
X_8292_ _0485_ _0500_ vssd1 vssd1 vccd1 vccd1 _3785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4455_ net282 vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__inv_2
X_7243_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[4\]
+ _2930_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__a31o_1
X_7174_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[6\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[7\]
+ _2885_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__and3_1
X_6125_ _2076_ _2077_ _2075_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__a21o_1
X_6056_ _2006_ _2007_ _2005_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_29_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _0794_ _0856_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout178_X net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6958_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[13\]
+ _2733_ _2734_ net158 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__o211a_1
X_5909_ _1860_ _1861_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__nand2_1
X_6889_ _2692_ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8628_ _4052_ _4106_ vssd1 vssd1 vccd1 vccd1 _4107_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8559_ net113 _3603_ _4037_ vssd1 vssd1 vccd1 vccd1 _4038_ sky130_fd_sc_hd__o21ba_1
XANTENNA__5019__A _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_86_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4858__A _0573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input20_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4864__Y _0817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_95_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8065__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5871__B _1774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4768__A _0719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9282__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9211__RESET_B net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5599__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7930_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] _3470_ vssd1
+ vssd1 vccd1 vccd1 _3471_ sky130_fd_sc_hd__or2_2
X_7861_ _3421_ _3422_ vssd1 vssd1 vccd1 vccd1 _3423_ sky130_fd_sc_hd__nor2_1
X_9600_ net464 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4790__X _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6812_ net275 _2640_ _2641_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__nor3_1
XANTENNA__8395__B1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7792_ _2368_ _2376_ _2382_ vssd1 vssd1 vccd1 vccd1 _3378_ sky130_fd_sc_hd__o21ai_1
X_6743_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[7\]
+ _2592_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__a21oi_1
X_9531_ net406 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_42_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9462_ net337 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_73_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6674_ team_08_WB.instance_to_wrap.allocation.game.det team_08_WB.instance_to_wrap.allocation.game.dinoJump.button
+ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_6_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5625_ _1575_ _1577_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout138_A _0817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8413_ net105 _3352_ _3355_ net103 vssd1 vssd1 vccd1 vccd1 _3894_ sky130_fd_sc_hd__a31o_1
XANTENNA__8762__A2_N net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9393_ clknet_leaf_28_wb_clk_i _0340_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5556_ net140 net145 vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__nand2b_1
X_8344_ _2293_ _2393_ _2426_ _3580_ _3635_ vssd1 vssd1 vccd1 vccd1 _3834_ sky130_fd_sc_hd__a221o_1
X_4507_ net29 net28 _0476_ _0477_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__or4_2
X_5487_ _1435_ _1438_ _1439_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__a21oi_1
X_8275_ _3498_ _3766_ _3768_ _3769_ vssd1 vssd1 vccd1 vccd1 _3770_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6476__A3 _2261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7226_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[0\]
+ _2922_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6893__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7157_ net645 net256 _2876_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__a21bo_1
X_6108_ _2019_ _2048_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__nand2_1
X_7088_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[6\]
+ _2799_ _2825_ _2828_ vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__a211o_1
XANTENNA__8622__A1 _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6039_ _1987_ _1988_ _1991_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8172__X _3691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8613__A _0685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5972__A _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4859__Y _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8310__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6872__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9385__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8523__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8129__B1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5410_ _1361_ _1362_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__nor2_2
XFILLER_0_3_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6390_ _2335_ _2340_ _0452_ _2330_ vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__o2bb2a_1
X_5341_ _1290_ _1292_ _1293_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_58_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8301__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8060_ _0432_ net139 vssd1 vssd1 vccd1 vccd1 _3593_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5666__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5272_ _1220_ _1223_ _1224_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__nand3_1
X_7011_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[2\] _2767_
+ _2768_ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8604__A1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8962_ net281 net153 _4438_ vssd1 vssd1 vccd1 vccd1 _4439_ sky130_fd_sc_hd__o21ai_1
XANTENNA__6615__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7913_ _3017_ _3454_ vssd1 vssd1 vccd1 vccd1 _3455_ sky130_fd_sc_hd__nor2_1
XANTENNA__8907__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8893_ net262 net236 _4370_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7844_ net159 _3409_ _3410_ net165 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout255_A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5506__A_N _1215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7775_ _3313_ _3363_ _3364_ vssd1 vssd1 vccd1 vccd1 _3365_ sky130_fd_sc_hd__a21oi_1
X_4987_ _0939_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__inv_6
X_6726_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__a21oi_1
X_9514_ net389 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XANTENNA__7991__B _3527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5792__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9445_ clknet_leaf_12_wb_clk_i _0390_ net217 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_6657_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[4\] _2537_ _2532_
+ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[4\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9376_ clknet_leaf_23_wb_clk_i _0324_ net253 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_5608_ _1558_ _1560_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__and2b_1
X_6588_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[9\] _2492_ net262
+ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__o21ai_1
X_5539_ _1074_ _1437_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__xnor2_2
X_8327_ _3460_ _3815_ _3817_ vssd1 vssd1 vccd1 vccd1 _3818_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8258_ net197 _3475_ _3753_ _3466_ net297 vssd1 vssd1 vccd1 vccd1 _3754_ sky130_fd_sc_hd__o221a_1
XANTENNA__8843__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_7209_ _0523_ _2908_ _2909_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__and3_1
X_8189_ net280 _0651_ vssd1 vssd1 vccd1 vccd1 _3706_ sky130_fd_sc_hd__xor2_1
Xfanout331 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[2\] vssd1
+ vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_2
Xfanout320 net323 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4855__B net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7512__A _0134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4590__B _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput39 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6310__B team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output51_A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4910_ _0810_ _0860_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__or2_2
X_5890_ _1795_ _1837_ _1842_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__nand3_2
XFILLER_0_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4841_ _0789_ _0793_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7560_ net625 team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr2\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr2\[0\] vssd1 vssd1 vccd1
+ vccd1 _3166_ sky130_fd_sc_hd__a21oi_1
X_4772_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[0\] vssd1
+ vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7491_ _3024_ _3074_ _3128_ _3130_ vssd1 vssd1 vccd1 vccd1 _3131_ sky130_fd_sc_hd__o211a_1
X_6511_ _2439_ _2440_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[6\]
+ sky130_fd_sc_hd__nor2_1
X_9230_ clknet_leaf_21_wb_clk_i _0058_ net240 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6442_ _0427_ _0641_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9161_ _0136_ _0132_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8112_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\] _3632_ _3639_
+ team_08_WB.instance_to_wrap.allocation.game.controller.state\[2\] vssd1 vssd1 vccd1
+ vccd1 _3640_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6373_ net261 _2324_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.collides
+ sky130_fd_sc_hd__and2_1
X_5324_ net128 _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_73_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9092_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[22\]
+ net209 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5255_ _1200_ _1206_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__or2_1
X_8043_ net318 _2426_ _3578_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[4\]
+ _3016_ vssd1 vssd1 vccd1 vccd1 _3579_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5186_ _0772_ _0859_ _0797_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__a21oi_2
XANTENNA__8147__B net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6890__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7986__B _0423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8945_ net126 _3678_ _4419_ _4421_ vssd1 vssd1 vccd1 vccd1 _4422_ sky130_fd_sc_hd__a211o_1
XANTENNA__5787__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout160_X net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8876_ _4234_ _4278_ _4348_ net98 _4353_ vssd1 vssd1 vccd1 vccd1 _4354_ sky130_fd_sc_hd__a221o_1
XANTENNA__8163__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4691__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7827_ _3395_ _3399_ vssd1 vssd1 vccd1 vccd1 _3400_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7758_ _3288_ _3306_ _3321_ _3324_ _3347_ vssd1 vssd1 vccd1 vccd1 _3348_ sky130_fd_sc_hd__o311a_1
XFILLER_0_85_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6709_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[10\]
+ _2568_ vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7689_ net99 net96 vssd1 vssd1 vccd1 vccd1 _3279_ sky130_fd_sc_hd__nor2_2
XFILLER_0_19_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8610__B _3280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9428_ clknet_leaf_39_wb_clk_i _0373_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9359_ clknet_leaf_26_wb_clk_i _0307_ net249 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6130__B _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4866__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout161 _2394_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_4
Xfanout183 _0668_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_2
Xfanout150 net151 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout172 net173 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7004__B1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8801__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5040_ _0901_ _0951_ _0990_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__nor3_1
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6991_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5942_ _1849_ _1893_ _1894_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_49_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8730_ _0421_ _3789_ _4197_ vssd1 vssd1 vccd1 vccd1 _4208_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5873_ _1818_ _1823_ _1824_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8661_ net135 _4136_ _4139_ vssd1 vssd1 vccd1 vccd1 _4140_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4824_ _0771_ _0775_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7612_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[10\]
+ net133 vssd1 vssd1 vccd1 vccd1 _3202_ sky130_fd_sc_hd__and2_1
X_8592_ _0686_ _4062_ vssd1 vssd1 vccd1 vccd1 _4071_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7543_ net550 _2581_ _3015_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__mux2_1
X_4755_ net163 _0696_ _0709_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9213_ clknet_leaf_18_wb_clk_i _0070_ net230 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4686_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__or2_2
X_7474_ _3044_ _3057_ _3074_ _3114_ vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__or4b_1
XFILLER_0_12_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6425_ net259 _2360_ _2375_ _2325_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__a32o_1
XANTENNA__9315__Q team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4957__Y _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6356_ net331 _2306_ _2307_ net327 vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9144_ clknet_leaf_36_wb_clk_i net510 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_5307_ _1052_ _1258_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__nor2_1
X_9075_ clknet_leaf_49_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[5\]
+ net236 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5134__X _1087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6287_ _2223_ _2226_ _2229_ _2239_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__or4_1
X_8026_ _3561_ vssd1 vssd1 vccd1 vccd1 _3562_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5238_ _1189_ _1190_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__and2b_1
X_5169_ _0903_ _0950_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__and2_1
XANTENNA__4973__X _0926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8928_ _3916_ _4401_ _4402_ net177 _0697_ vssd1 vssd1 vccd1 vccd1 _4405_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8859_ net186 _0519_ _4335_ vssd1 vssd1 vccd1 vccd1 _4337_ sky130_fd_sc_hd__nor3_1
XFILLER_0_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_30_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6 _0212_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7700__A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5220__A _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9236__RESET_B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6316__A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8250__B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[7\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[9\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_13_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9135__Q team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4471_ net627 vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__inv_2
X_6210_ _0943_ net123 vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__xor2_1
X_7190_ _2874_ _2896_ _2897_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6141_ _2092_ _2093_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__or2_1
XANTENNA__5867__A_N _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9319__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6072_ _1986_ _1997_ _2024_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__nand3_1
X_9533__489 vssd1 vssd1 vccd1 vccd1 net489 _9533__489/LO sky130_fd_sc_hd__conb_1
XANTENNA__7464__B1 _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5023_ _0746_ _0769_ _0974_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__nand3_1
XANTENNA__4793__X _0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout168_A _0723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6974_ _2744_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5925_ _1876_ _1877_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_85_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7519__A1 _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8713_ net136 _4181_ vssd1 vssd1 vccd1 vccd1 _4192_ sky130_fd_sc_hd__xnor2_1
X_5856_ _1804_ _1805_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8441__A _3355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8644_ _4121_ _4122_ vssd1 vssd1 vccd1 vccd1 _4123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4807_ _0753_ _0759_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__and2_4
XANTENNA__8192__A1 _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5787_ net131 _1688_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8575_ net109 _3596_ vssd1 vssd1 vccd1 vccd1 _4054_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout123_X net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4738_ _0680_ _0682_ _0681_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__o21bai_2
X_7526_ net511 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet vssd1 vssd1
+ vccd1 vccd1 _0246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6896__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4669_ _0620_ _0626_ _0619_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7457_ _0440_ _3054_ _3079_ vssd1 vssd1 vccd1 vccd1 _3099_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6408_ _2354_ _2358_ _2351_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7388_ _3023_ _3028_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__or2_1
X_9127_ clknet_leaf_38_wb_clk_i _0228_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_6339_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[2\] vssd1 vssd1 vccd1
+ vccd1 _2291_ sky130_fd_sc_hd__a21o_1
X_9058_ clknet_leaf_34_wb_clk_i _0193_ net246 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8009_ net196 _3545_ _3540_ vssd1 vssd1 vccd1 vccd1 _3546_ sky130_fd_sc_hd__o21ai_1
XANTENNA__8616__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6966__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8486__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7414__B net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4845__A1_N net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5869__B _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6046__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9070__RESET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5710_ _1660_ _1661_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5885__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9604__468 vssd1 vssd1 vccd1 vccd1 _9604__468/HI net468 sky130_fd_sc_hd__conb_1
X_6690_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[4\]
+ _2558_ net276 vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5641_ net132 _1544_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7921__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5572_ net128 _1524_ _1522_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8360_ team_08_WB.instance_to_wrap.allocation.game.controller.v\[2\] _3469_ vssd1
+ vssd1 vccd1 vccd1 _3847_ sky130_fd_sc_hd__nand2_1
X_4523_ net334 team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] _0491_
+ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__nand3_1
X_7311_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[3\] _2975_ _2978_
+ _2980_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__a211o_1
X_8291_ net139 _2275_ vssd1 vssd1 vccd1 vccd1 _3784_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7242_ net552 _2932_ _2934_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__a21oi_1
X_4454_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[4\] vssd1 vssd1
+ vccd1 vccd1 _0427_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7173_ net583 _2885_ _2886_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6124_ _2073_ _2074_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__xor2_1
X_6055_ _2005_ _2007_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__and2b_1
XANTENNA__5463__A2 _1410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5006_ _0785_ _0847_ _0884_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__a21o_2
XFILLER_0_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6957_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[12\]
+ _2730_ vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__nand3_2
XFILLER_0_64_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5908_ _1836_ _1845_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__xnor2_1
X_6888_ _2689_ _2691_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__or2_1
X_5839_ _0724_ _0910_ _1791_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8627_ net120 _4105_ vssd1 vssd1 vccd1 vccd1 _4106_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8558_ net118 _3606_ vssd1 vssd1 vccd1 vccd1 _4037_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7509_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\] _3143_
+ _3145_ _3022_ vssd1 vssd1 vccd1 vccd1 _3146_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8489_ net120 _3288_ vssd1 vssd1 vccd1 vccd1 _3969_ sky130_fd_sc_hd__nand2_1
XANTENNA__4858__B _0602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5151__A1 _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8065__B net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4593__B team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8928__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8156__A1 _3597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5914__B1 _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9251__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7860_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[7\]
+ _3416_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _3422_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8919__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6811_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8395__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7791_ net292 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1 vssd1
+ vccd1 vccd1 _3377_ sky130_fd_sc_hd__or2_1
X_6742_ net674 _2592_ _2594_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9530_ net405 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_9_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6673_ team_08_WB.instance_to_wrap.allocation.game.det team_08_WB.instance_to_wrap.allocation.game.dinoJump.button
+ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__and2b_1
X_9461_ clknet_leaf_37_wb_clk_i _0399_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.internalSck
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__8698__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5624_ _1499_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__nor2_1
X_9392_ clknet_leaf_20_wb_clk_i _0339_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_8412_ net99 _3892_ _3891_ _3330_ vssd1 vssd1 vccd1 vccd1 _3893_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8343_ net195 _3830_ _3832_ net170 vssd1 vssd1 vccd1 vccd1 _3833_ sky130_fd_sc_hd__a211o_1
XANTENNA__7370__A2 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5555_ _0907_ _1464_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4506_ net26 net25 vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__nand2_1
X_9539__495 vssd1 vssd1 vccd1 vccd1 net495 _9539__495/LO sky130_fd_sc_hd__conb_1
X_5486_ net129 _1390_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8274_ _2306_ net161 vssd1 vssd1 vccd1 vccd1 _3769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout200_A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9323__Q team_08_WB.instance_to_wrap.allocation.game.controller.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7225_ _2837_ _2922_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__nand2_1
X_7156_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[0\] net256 net164
+ _0539_ vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input5_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6107_ _1998_ _2012_ _2011_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_10_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7087_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[6\]
+ _2792_ _0429_ vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout190_X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6038_ _1990_ _1989_ vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__and2b_1
XANTENNA__5302__B _1254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8386__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7989_ _3524_ _3525_ vssd1 vssd1 vccd1 vccd1 _3527_ sky130_fd_sc_hd__or2_2
XANTENNA__8613__B net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8138__A1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5972__B _0926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8310__A1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7899__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8523__B net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4938__A1 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9640__487 vssd1 vssd1 vccd1 vccd1 _9640__487/HI net487 sky130_fd_sc_hd__conb_1
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5882__B _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5340_ _1237_ _1239_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_58_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7155__A _2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5271_ _0852_ _1222_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5666__A2 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7010_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[6\] team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5403__A _1353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8961_ _4435_ _4436_ _4437_ _4120_ vssd1 vssd1 vccd1 vccd1 _4438_ sky130_fd_sc_hd__o211a_1
X_7912_ net298 team_08_WB.instance_to_wrap.allocation.game.controller.state\[0\] _2427_
+ vssd1 vssd1 vccd1 vccd1 _3454_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8892_ _4231_ _4286_ _4288_ _4311_ _4369_ vssd1 vssd1 vccd1 vccd1 _4370_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7843_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[1\] team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[3\] vssd1
+ vssd1 vccd1 vccd1 _3410_ sky130_fd_sc_hd__a31o_1
X_4986_ _0919_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout150_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7774_ net153 net126 net116 _3359_ vssd1 vssd1 vccd1 vccd1 _3364_ sky130_fd_sc_hd__a31o_1
X_9513_ net388 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XANTENNA__5051__B1 _0999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6725_ net270 _2580_ _2582_ _2583_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout248_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9444_ clknet_leaf_6_wb_clk_i _0389_ net217 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6656_ _0649_ _2536_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9375_ clknet_leaf_23_wb_clk_i _0323_ net252 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_5607_ net141 net145 _0909_ net147 vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__a22o_1
XANTENNA__5792__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4689__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6587_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[9\] _2492_ vssd1
+ vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5538_ _1488_ _1490_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__nand2_1
X_8326_ net318 _3801_ vssd1 vssd1 vccd1 vccd1 _3817_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8257_ _2268_ net197 vssd1 vssd1 vccd1 vccd1 _3753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5469_ _1402_ _1421_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__xnor2_1
X_7208_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[19\] _2906_ vssd1
+ vssd1 vccd1 vccd1 _2909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout332 net333 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_2
Xfanout321 net323 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_4
X_8188_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\] _0692_ _0699_
+ vssd1 vssd1 vccd1 vccd1 _3705_ sky130_fd_sc_hd__and3_1
Xfanout310 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_2
XANTENNA__8056__B1 _3511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7139_ _2850_ _2868_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4599__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4856__B1 _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8093__X _3622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8534__A _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4840_ net144 net140 vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__nor2_4
XFILLER_0_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6989__A team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5893__A _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6781__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4771_ _0721_ _0722_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__or2_4
XFILLER_0_56_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6510_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[6\] _2437_
+ _2429_ vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7490_ _0440_ _3054_ _3057_ _3129_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6441_ _0427_ _0641_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_77_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5887__A2 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6372_ _0645_ _2320_ _2322_ _2323_ _2290_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__a41o_2
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9160_ _0135_ _0131_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_5323_ _1272_ _1274_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__xnor2_1
X_8111_ _0646_ _3638_ vssd1 vssd1 vccd1 vccd1 _3639_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9091_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[21\]
+ net222 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8709__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5254_ _1200_ _1206_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__nand2_1
X_8042_ net199 _3575_ _3576_ _3577_ vssd1 vssd1 vccd1 vccd1 _3578_ sky130_fd_sc_hd__a31o_1
X_5185_ _1136_ _1137_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout198_A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8589__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_8944_ net134 _4418_ _4420_ vssd1 vssd1 vccd1 vccd1 _4421_ sky130_fd_sc_hd__o21ai_1
X_8875_ _4349_ _4352_ net98 _4348_ vssd1 vssd1 vccd1 vccd1 _4353_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_66_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7826_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[0\] team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\] vssd1
+ vssd1 vccd1 vccd1 _3399_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_35_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8761__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4969_ _0727_ _0920_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__or2_4
XFILLER_0_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7757_ _3286_ _3287_ net153 vssd1 vssd1 vccd1 vccd1 _3347_ sky130_fd_sc_hd__a21o_1
X_6708_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[10\]
+ _2568_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7688_ net104 net101 vssd1 vssd1 vccd1 vccd1 _3278_ sky130_fd_sc_hd__nand2_2
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6639_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[28\] _2524_
+ net255 vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__a21oi_1
X_9427_ clknet_leaf_43_wb_clk_i _0372_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9358_ clknet_leaf_27_wb_clk_i _0306_ net251 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_9289_ clknet_leaf_14_wb_clk_i _0108_ net213 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_8309_ net325 net322 _3776_ vssd1 vssd1 vccd1 vccd1 _3801_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4866__B _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9550__418 vssd1 vssd1 vccd1 vccd1 _9550__418/HI net418 sky130_fd_sc_hd__conb_1
XFILLER_0_100_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout140 _0791_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_4
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_2
Xfanout151 net152 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_2
Xfanout173 _3179_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_2
XANTENNA__5978__A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout195 _3460_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_4
Xfanout184 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[12\]
+ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7004__A1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8801__B _3266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7307__A2 _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5218__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9095__RESET_B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9024__RESET_B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8529__A _3261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9490__365 vssd1 vssd1 vccd1 vccd1 _9490__365/HI net365 sky130_fd_sc_hd__conb_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8070__A2_N net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6991__B team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6990_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__and2b_1
XANTENNA__4792__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6336__X _2288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5941_ net147 _0927_ _1847_ _1848_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5872_ _1823_ _1824_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_8660_ _4120_ _4133_ _4138_ vssd1 vssd1 vccd1 vccd1 _4139_ sky130_fd_sc_hd__a21bo_1
X_4823_ _0771_ _0775_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7611_ _3195_ _3198_ _3199_ vssd1 vssd1 vccd1 vccd1 _3201_ sky130_fd_sc_hd__or3_1
X_8591_ _4062_ _4069_ vssd1 vssd1 vccd1 vccd1 _4070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4754_ _0686_ _0707_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7542_ _0443_ net543 _2545_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7473_ net306 _3051_ _3060_ net307 vssd1 vssd1 vccd1 vccd1 _3114_ sky130_fd_sc_hd__o22a_1
X_9212_ clknet_leaf_18_wb_clk_i _0069_ net230 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4685_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6424_ _2364_ _2374_ vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout113_A _3234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6355_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[3\] _2291_ vssd1
+ vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_8_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9143_ clknet_leaf_36_wb_clk_i net527 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__8439__A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5306_ _1052_ _1199_ _1257_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__and3_1
X_6286_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[3\]
+ _2228_ _2231_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[2\]
+ _2238_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9074_ clknet_leaf_44_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[4\]
+ net236 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5237_ _1187_ _1188_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8025_ _3559_ _3560_ vssd1 vssd1 vccd1 vccd1 _3561_ sky130_fd_sc_hd__nand2_2
XANTENNA__5493__A0 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5168_ _1115_ _1120_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5099_ _1051_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout270_X net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8927_ _0696_ _3179_ _4097_ vssd1 vssd1 vccd1 vccd1 _4404_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8858_ _0519_ _4335_ net186 vssd1 vssd1 vccd1 vccd1 _4336_ sky130_fd_sc_hd__o21a_1
X_7809_ _2972_ _3386_ vssd1 vssd1 vccd1 vccd1 _3390_ sky130_fd_sc_hd__nor2_1
X_8789_ net323 _4262_ vssd1 vssd1 vccd1 vccd1 _4267_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6422__A _2368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9474__349 vssd1 vssd1 vccd1 vccd1 _9474__349/HI net349 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_18_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataShift\[1\]
+ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7700__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6316__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5507__B1_N _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8812__A _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8731__A1_N net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8725__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6736__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8725__B2 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8531__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7715__X _3305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4470_ net308 vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4787__A _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6140_ _2078_ _2079_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__xor2_1
XANTENNA__8815__A_N net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7464__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6071_ _1982_ _2022_ _2023_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__and3_1
X_5022_ _0746_ _0769_ _0974_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8413__B1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8706__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5411__A _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6973_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[19\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[18\]
+ _2741_ vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__and3_1
X_5924_ _1829_ _1830_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_85_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8712_ _0427_ net119 vssd1 vssd1 vccd1 vccd1 _4191_ sky130_fd_sc_hd__or2_1
X_5855_ _0814_ _0922_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_24_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8643_ net283 net281 _2538_ vssd1 vssd1 vccd1 vccd1 _4122_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout230_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4806_ _0583_ _0596_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5786_ _1736_ _1738_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8574_ _4037_ _4051_ _4052_ vssd1 vssd1 vccd1 vccd1 _4053_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9326__Q team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4737_ _0687_ _0690_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7525_ net509 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet vssd1 vssd1
+ vccd1 vccd1 _0245_ sky130_fd_sc_hd__mux2_1
XANTENNA__4968__Y _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4668_ _0623_ _0624_ _0622_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7456_ net516 net115 _3070_ _3098_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout116_X net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4697__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6407_ _2328_ _2348_ _2357_ _2356_ _2334_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__o32a_4
XFILLER_0_101_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4599_ net256 _0535_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7387_ net630 _3028_ _3035_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9126_ clknet_leaf_41_wb_clk_i _0227_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_6338_ net315 _2278_ _2288_ _2289_ _0684_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__a2111oi_1
X_6269_ _2111_ _2221_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__nand2_1
X_9057_ clknet_leaf_35_wb_clk_i _0192_ net245 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_8008_ net321 _3544_ _3534_ vssd1 vssd1 vccd1 vccd1 _3545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7520__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5941__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9556__424 vssd1 vssd1 vccd1 vccd1 _9556__424/HI net424 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_10_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8526__B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8542__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5758__A1_N net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5885__B _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5640_ net131 _1592_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5571_ _1522_ _1523_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9496__371 vssd1 vssd1 vccd1 vccd1 _9496__371/HI net371 sky130_fd_sc_hd__conb_1
XFILLER_0_54_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8290_ _3479_ _3771_ _3783_ net235 net675 vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__o32a_1
X_4522_ _0489_ _0490_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__and2_2
X_7310_ net636 _2974_ _2981_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4453_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\] vssd1 vssd1
+ vccd1 vccd1 _0426_ sky130_fd_sc_hd__inv_2
X_7241_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[5\]
+ _2932_ net181 vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7172_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[6\] _2885_ _0523_
+ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6123_ _0761_ _0917_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__nor2_1
X_6054_ _1964_ _2004_ _2003_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5005_ _0956_ _0957_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6660__A2 _2532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A _0637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8937__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6956_ _2733_ net157 _2732_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__and3b_1
XFILLER_0_48_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5907_ _0919_ _1859_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6887_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ _2688_ _2690_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__or4b_1
XFILLER_0_37_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5838_ _0718_ net146 vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8626_ _0668_ _3602_ _4090_ vssd1 vssd1 vccd1 vccd1 _4105_ sky130_fd_sc_hd__a21o_1
X_5769_ _0919_ _1721_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8557_ _3355_ _3901_ net102 _3280_ vssd1 vssd1 vccd1 vccd1 _4036_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_86_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7508_ net302 _0442_ _3144_ _0438_ vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__a211o_1
XANTENNA__4698__Y _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7515__B _3040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8488_ _3282_ _3338_ _3967_ vssd1 vssd1 vccd1 vccd1 _3968_ sky130_fd_sc_hd__nor3_1
XANTENNA__8873__B1 _3272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7439_ _3082_ vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9109_ clknet_leaf_40_wb_clk_i net504 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__8627__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4874__B _0825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8928__A1 _3916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8928__B2 _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7706__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9530__405 vssd1 vssd1 vccd1 vccd1 _9530__405/HI net405 sky130_fd_sc_hd__conb_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8919__B2 _0674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5896__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6810_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9291__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7790_ team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] _2325_ _3376_ net261
+ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__a22o_1
X_6741_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[7\]
+ _2592_ net272 vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9460_ clknet_leaf_45_wb_clk_i _0398_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_floor
+ sky130_fd_sc_hd__dfxtp_1
X_6672_ net563 _2546_ _2544_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__a21bo_1
X_5623_ _0749_ _1498_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__and2_1
X_9391_ clknet_leaf_28_wb_clk_i _0338_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8411_ _0425_ _0558_ net104 vssd1 vssd1 vccd1 vccd1 _3892_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8342_ net314 _3817_ _3831_ net198 vssd1 vssd1 vccd1 vccd1 _3832_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5554_ _0786_ _1506_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_42_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5485_ net131 _1437_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__nand2_1
X_4505_ net22 net21 net24 net23 vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__or4_1
XANTENNA__5136__A _1087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8273_ net330 net194 _3511_ _3767_ vssd1 vssd1 vccd1 vccd1 _3768_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7054__C team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7224_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.state\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.state\[0\] vssd1
+ vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__and2b_1
XANTENNA__6330__B2 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6330__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7155_ _2874_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__inv_2
X_6106_ _2057_ _2058_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7086_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[6\]
+ _2789_ _2800_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[6\]
+ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__a22o_1
X_6037_ _1987_ _1988_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7988_ _3524_ _3525_ vssd1 vssd1 vccd1 vccd1 _3526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6939_ _2404_ _2722_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7897__A1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8609_ net190 _3284_ _3271_ net187 vssd1 vssd1 vccd1 vccd1 _4088_ sky130_fd_sc_hd__a211o_1
XANTENNA__4502__X _0473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9589_ net453 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_84_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8310__A2 _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9633__484 vssd1 vssd1 vccd1 vccd1 _9633__484/HI net484 sky130_fd_sc_hd__conb_1
XANTENNA__4885__A _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout96_X net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8074__A1 _3597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8092__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7585__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8129__A2 _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5270_ _0852_ _1222_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8960_ net281 net155 net136 net285 vssd1 vssd1 vccd1 vccd1 _4437_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_7911_ net559 _0713_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8891_ _4225_ _4327_ _4328_ _4357_ _4368_ vssd1 vssd1 vccd1 vccd1 _4369_ sky130_fd_sc_hd__a311o_1
XFILLER_0_77_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7842_ _3408_ vssd1 vssd1 vccd1 vccd1 _3409_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4985_ _0934_ _0937_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__nor2_2
XANTENNA__4929__A2 _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7773_ net153 net133 _3291_ vssd1 vssd1 vccd1 vccd1 _3363_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout143_A _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6724_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__nand2_1
X_9512_ net387 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_74_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9443_ clknet_leaf_6_wb_clk_i _0388_ net211 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6655_ _0426_ _2535_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__nor2_2
X_9374_ clknet_leaf_24_wb_clk_i _0322_ net252 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_5606_ net140 _0905_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6586_ _2492_ _2478_ _2491_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[8\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_15_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5537_ net131 _1489_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__nand2_1
X_8325_ net320 net316 vssd1 vssd1 vccd1 vccd1 _3816_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8256_ net333 _3476_ net195 vssd1 vssd1 vccd1 vccd1 _3752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5468_ _0940_ _1374_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__xnor2_4
X_7207_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[19\] _2906_ vssd1
+ vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5399_ _1349_ _1350_ _1351_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__or3_1
Xfanout300 team_08_WB.instance_to_wrap.allocation.game.controller.state\[4\] vssd1
+ vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_4
X_8187_ _0710_ _3703_ _2418_ vssd1 vssd1 vccd1 vccd1 _3704_ sky130_fd_sc_hd__a21o_1
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout311 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.frameBufferLowNibble
+ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_8
XANTENNA__8056__A1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout333 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[1\] vssd1
+ vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7138_ _2868_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__inv_2
XANTENNA__4992__X _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7069_ net293 _2814_ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8359__A2 _2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__8640__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput19 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5504__A _1217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6989__B team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4770_ _0721_ _0722_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6440_ _0648_ _2386_ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_77_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6371_ _0428_ net279 vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__and2_1
X_5322_ _1274_ _1272_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_51_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8110_ net283 _0645_ vssd1 vssd1 vccd1 vccd1 _3638_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9090_ clknet_leaf_50_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[20\]
+ net222 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8709__B _3241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5253_ _1202_ _1204_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__xnor2_1
X_8041_ net318 net194 net170 vssd1 vssd1 vccd1 vccd1 _3577_ sky130_fd_sc_hd__a21o_1
XANTENNA__7613__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5184_ _1133_ _1135_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8943_ net152 _3696_ vssd1 vssd1 vccd1 vccd1 _4420_ sky130_fd_sc_hd__or2_1
X_8874_ net101 _3543_ _4350_ _3526_ _4351_ vssd1 vssd1 vccd1 vccd1 _4352_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout260_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7825_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[1\]
+ _3395_ _3396_ _3398_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9329__Q team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4968_ _0727_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__nor2_4
X_7756_ net174 net117 _3325_ _3345_ vssd1 vssd1 vccd1 vccd1 _3346_ sky130_fd_sc_hd__o31a_1
XFILLER_0_80_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4899_ _0808_ _0815_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__nand2_4
XFILLER_0_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6707_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[10\]
+ _2568_ _2570_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7687_ _3263_ _3275_ vssd1 vssd1 vccd1 vccd1 _3277_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9426_ clknet_leaf_43_wb_clk_i _0371_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_6638_ _2524_ _2525_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[27\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_22_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9357_ clknet_leaf_26_wb_clk_i _0305_ net249 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8308_ _3798_ _3799_ vssd1 vssd1 vccd1 vccd1 _3800_ sky130_fd_sc_hd__and2_1
X_6569_ _2481_ net263 _2480_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[2\]
+ sky130_fd_sc_hd__and3b_1
X_9288_ clknet_leaf_14_wb_clk_i _0107_ net213 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8239_ _3034_ _3739_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__nand2_1
Xfanout130 net132 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_1
XANTENNA__5324__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9323__RESET_B net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout141 _0782_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
Xfanout163 _0684_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_2
Xfanout174 net175 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_2
Xfanout152 _3187_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_4
Xfanout196 net199 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__buf_2
XANTENNA__5978__B _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7004__A2 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6212__B1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8370__A team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6602__B net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6279__B1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9064__RESET_B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7779__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4792__B _0743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5940_ _1890_ _1891_ _1846_ _1889_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5871_ _1773_ _1774_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_66_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7610_ _3195_ _3198_ _3199_ vssd1 vssd1 vccd1 vccd1 _3200_ sky130_fd_sc_hd__nor3_2
X_4822_ _0577_ _0598_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8590_ net178 _4061_ vssd1 vssd1 vccd1 vccd1 _4069_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4753_ _0707_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7541_ net593 _3156_ _2545_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7472_ _3048_ _3112_ _3059_ _3056_ vssd1 vssd1 vccd1 vccd1 _3113_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9211_ clknet_leaf_18_wb_clk_i net587 net231 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4684_ net287 net284 vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__or2_1
X_6423_ _2358_ _2373_ _2363_ vssd1 vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8259__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6354_ _2291_ _2305_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_8_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9142_ clknet_leaf_38_wb_clk_i _0243_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout106_A _3252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5305_ _1199_ _1257_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6285_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[2\]
+ _2231_ _2233_ _2237_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__o211ai_1
X_9073_ clknet_leaf_49_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[3\]
+ net224 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5236_ _1187_ _1188_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8024_ net321 net317 _3524_ vssd1 vssd1 vccd1 vccd1 _3560_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6690__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5167_ _1118_ _1119_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__nand2_1
XANTENNA__4983__A _0809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5098_ _1012_ _1050_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8926_ net169 _3200_ _4100_ _4396_ vssd1 vssd1 vccd1 vccd1 _4403_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8857_ net331 _0422_ vssd1 vssd1 vccd1 vccd1 _4335_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7808_ net628 _2975_ _3388_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__a21o_1
XANTENNA__8190__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8788_ _4264_ _4265_ vssd1 vssd1 vccd1 vccd1 _4266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7739_ _3265_ _3276_ vssd1 vssd1 vccd1 vccd1 _3329_ sky130_fd_sc_hd__nand2_2
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9409_ clknet_leaf_31_wb_clk_i _0356_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input36_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold8 _0250_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8812__B _0425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8186__B1 _0696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7933__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4787__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6070_ net182 _0860_ _1980_ _1981_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__o22ai_1
XANTENNA__8661__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5021_ _0972_ _0973_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8413__A1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6972_ _2743_ net158 _2742_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__and3b_1
XFILLER_0_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8711_ _0427_ net119 _4186_ _4189_ vssd1 vssd1 vccd1 vccd1 _4190_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_85_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5923_ _1872_ _1875_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5854_ _0813_ _0921_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8642_ net283 _2538_ net281 vssd1 vssd1 vccd1 vccd1 _4121_ sky130_fd_sc_hd__a21oi_1
X_4805_ _0757_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__inv_2
X_8573_ net111 _3603_ vssd1 vssd1 vccd1 vccd1 _4052_ sky130_fd_sc_hd__xnor2_1
X_5785_ net132 _1737_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7524_ net526 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.data\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet vssd1 vssd1
+ vccd1 vccd1 _0244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout223_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4736_ net169 _0690_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4667_ _0623_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__and2_1
X_7455_ _3023_ _3096_ _3097_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7386_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\] _3022_
+ _3028_ _3034_ vssd1 vssd1 vccd1 vccd1 _3035_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout109_X net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6406_ team_08_WB.instance_to_wrap.allocation.game.game.score\[3\] _2327_ vssd1 vssd1
+ vccd1 vccd1 _2357_ sky130_fd_sc_hd__nor2_1
X_4598_ _0492_ _0559_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__and2_1
X_6337_ _2282_ _2283_ _2284_ _0697_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__a31o_1
X_9125_ clknet_leaf_40_wb_clk_i _0226_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.tft_reset
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6268_ _2095_ _2102_ _2110_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__nand3_1
X_9056_ clknet_leaf_34_wb_clk_i _0191_ net248 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_6199_ _1137_ _2150_ _1136_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__a21o_1
X_5219_ _0943_ _1171_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__nand2_1
X_8007_ _3541_ _3542_ vssd1 vssd1 vccd1 vccd1 _3544_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5602__A _1087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8909_ _0689_ net118 _4010_ vssd1 vssd1 vccd1 vccd1 _4386_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5049__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5016__A_N _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9388__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8823__A _0423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5570_ _1507_ _1519_ _1521_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4521_ net332 team_08_WB.instance_to_wrap.allocation.game.controller.v\[1\] vssd1
+ vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4452_ net185 vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__inv_2
X_7240_ _2932_ _2933_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7171_ net164 _2884_ _2885_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6122_ _2073_ _2074_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_0_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6053_ _0761_ _0921_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_37_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6645__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5004_ _0943_ _0955_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__or2_1
XANTENNA__5422__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout173_A _3179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6955_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[12\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[11\]
+ _2729_ vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__and3_1
X_5906_ _1856_ _1857_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6886_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2690_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8625_ _4090_ _4091_ _4099_ _4103_ vssd1 vssd1 vccd1 vccd1 _4104_ sky130_fd_sc_hd__a211oi_1
X_5837_ _1746_ _1748_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5768_ _1719_ _1720_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8556_ _4027_ _4034_ _4001_ vssd1 vssd1 vccd1 vccd1 _4035_ sky130_fd_sc_hd__o21a_1
X_4719_ _0672_ _0673_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__xor2_2
X_7507_ _3091_ _3122_ _3093_ net303 vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__a211oi_1
X_8487_ net185 _0555_ net188 vssd1 vssd1 vccd1 vccd1 _3967_ sky130_fd_sc_hd__or3b_1
XFILLER_0_86_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5699_ _0772_ net145 _1648_ _1651_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7438_ net305 _3042_ _3044_ _3059_ _3081_ vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__o311a_1
XFILLER_0_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_7369_ net277 _2421_ _2423_ vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_55_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9108_ clknet_leaf_40_wb_clk_i _0211_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_9039_ clknet_leaf_7_wb_clk_i _0174_ net211 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoMovement
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7061__B1 _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5072__C1 _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8930__X _4407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5914__A2 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7706__B net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5242__A _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_9610__474 vssd1 vssd1 vccd1 vccd1 _9610__474/HI net474 sky130_fd_sc_hd__conb_1
XANTENNA__8919__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6740_ _2592_ _2593_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6671_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[1\] _2545_
+ vssd1 vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__and3_1
X_5622_ _0747_ _1574_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__nor2_1
X_9390_ clknet_leaf_28_wb_clk_i _0337_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8410_ _3887_ _3889_ vssd1 vssd1 vccd1 vccd1 _3891_ sky130_fd_sc_hd__nor2_1
X_5553_ _1465_ _1466_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__xnor2_1
X_8341_ net314 _3817_ vssd1 vssd1 vccd1 vccd1 _3831_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4504_ net13 net12 net14 net15 vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__or4b_1
XFILLER_0_53_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5484_ _1435_ _1436_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_91_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8272_ net193 _3495_ vssd1 vssd1 vccd1 vccd1 _3767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5136__B _1088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6866__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7223_ _2911_ _2919_ _2920_ _2921_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7154_ net256 _0546_ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__nor2_4
XFILLER_0_1_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6105_ _2028_ _2056_ _2055_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5152__A _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7085_ _2819_ _2825_ _2827_ _2818_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__o31a_1
XANTENNA__8083__A2 _3608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6036_ _1901_ _1904_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4991__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5841__A1 _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout176_X net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7987_ net328 net325 vssd1 vssd1 vccd1 vccd1 _3525_ sky130_fd_sc_hd__nor2_1
X_6938_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[6\]
+ _2403_ net157 vssd1 vssd1 vccd1 vccd1 _2722_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6869_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[8\]
+ _2675_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9588_ net452 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8608_ _4035_ _4060_ _4085_ _4086_ _0694_ vssd1 vssd1 vccd1 vccd1 _4087_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_49_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8539_ _4016_ _4017_ vssd1 vssd1 vccd1 vccd1 _4018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8357__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5062__A _1011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7585__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7717__A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8298__C1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9440__Q team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7812__A2 _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8283__A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7910_ net547 _0713_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__and2_1
X_8890_ _4323_ _4367_ vssd1 vssd1 vccd1 vccd1 _4368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7841_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[1\] team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[3\] vssd1
+ vssd1 vccd1 vccd1 _3408_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_19_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4984_ _0921_ _0926_ _0929_ _0931_ _0810_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__a41o_1
XFILLER_0_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7772_ net176 _3361_ vssd1 vssd1 vccd1 vccd1 _3362_ sky130_fd_sc_hd__nor2_1
X_6723_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2582_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9511_ net386 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9442_ clknet_leaf_5_wb_clk_i _0387_ net214 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_6654_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5605_ net141 _0909_ _1557_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout136_A _3200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9373_ clknet_leaf_24_wb_clk_i _0321_ net252 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6585_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[7\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[8\]
+ _2488_ vssd1 vssd1 vccd1 vccd1 _2492_ sky130_fd_sc_hd__and3_1
X_5536_ _1486_ _1487_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__xnor2_1
X_8324_ net318 _3801_ vssd1 vssd1 vccd1 vccd1 _3815_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5467_ _0939_ _1419_ _1418_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__a21o_1
XANTENNA__4986__A _0919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8255_ net615 net242 _3020_ _3751_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7206_ net570 _2904_ _2907_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__o21a_1
X_5398_ _0766_ _0971_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__nor2_1
X_8186_ net163 _0709_ _0696_ vssd1 vssd1 vccd1 vccd1 _3703_ sky130_fd_sc_hd__o21ai_1
Xfanout323 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[5\] vssd1
+ vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_2
Xfanout301 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_4
Xfanout312 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.frameBufferLowNibble
+ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_4
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7137_ _2865_ _2867_ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__nor2_2
X_7068_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\]
+ _2781_ _2790_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__or3_1
X_6019_ _1931_ _1932_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5610__A _0825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8640__B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8819__B2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6351__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9435__Q team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6370_ net287 _0648_ net285 vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__a21oi_1
X_5321_ _1225_ _1273_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8040_ _3548_ _3552_ _3571_ _3574_ vssd1 vssd1 vccd1 vccd1 _3576_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9616__480 vssd1 vssd1 vccd1 vccd1 _9616__480/HI net480 sky130_fd_sc_hd__conb_1
X_5252_ _1202_ _1204_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5183_ _1133_ _1135_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8942_ net152 _3696_ _4418_ net134 vssd1 vssd1 vccd1 vccd1 _4419_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8873_ _3526_ _4350_ _3272_ vssd1 vssd1 vccd1 vccd1 _4351_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout253_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7824_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\]
+ _2781_ _2793_ _2795_ vssd1 vssd1 vccd1 vccd1 _3398_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_35_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4967_ _0624_ _0725_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7755_ _3344_ vssd1 vssd1 vccd1 vccd1 _3345_ sky130_fd_sc_hd__inv_2
X_4898_ _0846_ _0850_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__or2_1
X_6706_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[10\]
+ _2568_ net273 vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout139_X net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7686_ _3263_ _3275_ vssd1 vssd1 vccd1 vccd1 _3276_ sky130_fd_sc_hd__nor2_4
XFILLER_0_62_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9425_ clknet_leaf_43_wb_clk_i _0370_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_6637_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[27\] _2523_
+ net260 vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9356_ clknet_leaf_26_wb_clk_i _0304_ net249 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4535__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6568_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _2481_ sky130_fd_sc_hd__and3_1
XANTENNA__7644__X _3234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4987__Y _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5519_ _1470_ _1471_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8307_ _3555_ _3785_ _3787_ vssd1 vssd1 vccd1 vccd1 _3799_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5605__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9287_ clknet_leaf_14_wb_clk_i _0130_ net214 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8188__A team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6499_ _2431_ _2432_ net156 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_30_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8238_ _2996_ _3738_ net122 vssd1 vssd1 vccd1 vccd1 _3739_ sky130_fd_sc_hd__a21o_1
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_4
X_8169_ net284 _3677_ _0650_ vssd1 vssd1 vccd1 vccd1 _3688_ sky130_fd_sc_hd__a21boi_1
Xfanout120 _3224_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_4
Xfanout142 _0782_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
Xfanout164 _0524_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_4
Xfanout153 net154 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_4
Xfanout197 net199 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_4
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_2
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_2
XFILLER_0_96_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8651__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6212__A1 _1039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7960__A1 _2393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5058__Y _1011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5515__A _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6279__B2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8826__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7779__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5250__A _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5870_ _1822_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4821_ _0738_ _0772_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_66_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6668__A_N team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6081__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4752_ _0669_ net178 vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7540_ _3154_ _3155_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4683_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.cactusMovement net294
+ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__nand2_1
X_7471_ _3084_ _3092_ vssd1 vssd1 vccd1 vccd1 _3112_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9210_ clknet_leaf_18_wb_clk_i _0063_ net230 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6422_ _2368_ _2371_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__nand2_1
X_9141_ clknet_leaf_38_wb_clk_i _0242_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6353_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[2\] team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusHeight1\[0\] vssd1 vssd1 vccd1
+ vccd1 _2305_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5304_ _1197_ _1198_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nand2_1
X_6284_ _2234_ _2235_ _2236_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__and3_1
X_9072_ clknet_leaf_49_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[2\]
+ net224 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5235_ _1074_ _1132_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5144__B _0825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8023_ net321 _3524_ net317 vssd1 vssd1 vccd1 vccd1 _3559_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_41_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5166_ _0943_ _1117_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__or2_1
X_5097_ _1048_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8925_ _0705_ net118 _4397_ vssd1 vssd1 vccd1 vccd1 _4402_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8856_ _3789_ _4329_ vssd1 vssd1 vccd1 vccd1 _4334_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5999_ _1948_ _1949_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__xor2_1
X_7807_ _0450_ _2974_ _3389_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__o21ai_1
X_8787_ net324 net323 _4261_ net316 vssd1 vssd1 vccd1 vccd1 _4265_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7738_ _3311_ _3327_ _3285_ vssd1 vssd1 vccd1 vccd1 _3328_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7815__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9408_ clknet_leaf_31_wb_clk_i _0355_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_7669_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[4\]
+ _3247_ _3254_ _3258_ vssd1 vssd1 vccd1 vccd1 _3259_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9339_ clknet_leaf_26_wb_clk_i _0004_ net249 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5054__B _0998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold9 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.dataDc vssd1
+ vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8422__A2 _3355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8186__A1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8381__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7933__A1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7709__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5172__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5245__A _1194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9285__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5020_ _0748_ _0971_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9214__RESET_B net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6971_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[18\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[17\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[16\]
+ _2737_ vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8710_ _4187_ _4188_ _4185_ vssd1 vssd1 vccd1 vccd1 _4189_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_85_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5922_ _1874_ _1873_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8291__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9540__408 vssd1 vssd1 vccd1 vccd1 _9540__408/HI net408 sky130_fd_sc_hd__conb_1
X_5853_ _1805_ _1804_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8641_ net279 net173 vssd1 vssd1 vccd1 vccd1 _4120_ sky130_fd_sc_hd__or2_2
X_5784_ _1734_ _1735_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4804_ net144 _0750_ net167 _0741_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__o31a_2
X_8572_ net118 _3606_ _4042_ _4050_ vssd1 vssd1 vccd1 vccd1 _4051_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_90_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4735_ _0663_ net178 _0689_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__and3_1
X_7523_ net303 _3152_ net301 vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout216_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4666_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[1\] vssd1
+ vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7454_ _3059_ _3094_ _3090_ _3057_ vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_101_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5163__A1 _1087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4597_ net334 team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] _0491_
+ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7385_ _3028_ _3033_ vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__or2_2
X_6405_ _2343_ _2355_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6336_ net315 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[6\] _2285_
+ _2287_ _0685_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__a221o_1
X_9124_ clknet_leaf_41_wb_clk_i _0225_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_9055_ clknet_leaf_34_wb_clk_i _0190_ net246 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4994__A _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6267_ _2112_ _2219_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__or2_1
X_6198_ _1138_ _2150_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__nand2_1
X_5218_ net123 _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__xor2_1
X_8006_ _3541_ _3542_ vssd1 vssd1 vccd1 vccd1 _3543_ sky130_fd_sc_hd__nor2_2
X_5149_ _1096_ _1098_ _1100_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__or3b_1
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8908_ _4379_ _4384_ vssd1 vssd1 vccd1 vccd1 _4385_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7915__A1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8839_ _0521_ _3816_ net95 vssd1 vssd1 vccd1 vccd1 _4317_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9480__355 vssd1 vssd1 vccd1 vccd1 _9480__355/HI net355 sky130_fd_sc_hd__conb_1
XFILLER_0_19_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9521__396 vssd1 vssd1 vccd1 vccd1 _9521__396/HI net396 sky130_fd_sc_hd__conb_1
XFILLER_0_34_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7832__X _3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8823__B net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7158__C net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5264__A2_N _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6590__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4798__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4520_ net332 team_08_WB.instance_to_wrap.allocation.game.controller.v\[1\] vssd1
+ vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9443__Q team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4451_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__inv_2
X_7170_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[5\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[4\]
+ _2881_ vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6121_ _2039_ _2040_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8557__Y _4036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5262__X _1215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5703__A _1048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7190__A _2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8095__B1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6052_ _1964_ _2003_ _2004_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5003_ _0943_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9464__339 vssd1 vssd1 vccd1 vccd1 _9464__339/HI net339 sky130_fd_sc_hd__conb_1
XFILLER_0_89_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6954_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[12\]
+ _2730_ vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout166_A _3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5905_ _1856_ _1857_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6885_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[9\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_17_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8624_ _4092_ _4095_ _4102_ vssd1 vssd1 vccd1 vccd1 _4103_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_101_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5836_ _1753_ _1788_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout333_A team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8570__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4989__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5767_ _1715_ _1717_ _1718_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7365__A team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8555_ _4008_ _4011_ _4026_ _4033_ vssd1 vssd1 vccd1 vccd1 _4034_ sky130_fd_sc_hd__a31o_1
X_5698_ net147 _0906_ _1650_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4718_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[4\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[4\]
+ _0666_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__a21oi_2
X_7506_ _0437_ _3142_ _3134_ net301 vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__a211o_1
X_8486_ net99 net104 _3965_ _3330_ vssd1 vssd1 vccd1 vccd1 _3966_ sky130_fd_sc_hd__o31a_1
XFILLER_0_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4649_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[6\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[6\] vssd1
+ vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__and2b_1
X_7437_ net309 _3080_ _3079_ vssd1 vssd1 vccd1 vccd1 _3081_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7368_ net565 net244 _2423_ _3019_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__o22a_1
X_7299_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.drawDoneCactus _2323_
+ vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__and2_1
X_6319_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[3\] _2265_ vssd1
+ vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__xnor2_2
X_9107_ clknet_leaf_39_wb_clk_i _0210_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5613__A _1087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9038_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[20\]
+ net208 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4647__B1 _0573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7061__B2 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9562__430 vssd1 vssd1 vccd1 vccd1 _9562__430/HI net430 sky130_fd_sc_hd__conb_1
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7364__A2 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_86_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7355__A2 _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6670_ _2545_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__inv_2
X_5621_ net141 _0859_ _1088_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__a21oi_1
XANTENNA__6801__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5552_ _1502_ _1504_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__or2_1
X_8340_ _3828_ _3829_ vssd1 vssd1 vccd1 vccd1 _3830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4503_ net18 net17 net20 net19 vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__or4_1
XANTENNA__8304__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8304__B2 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8271_ net196 _3761_ _3765_ _3540_ vssd1 vssd1 vccd1 vccd1 _3766_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5483_ _1429_ _1433_ _1434_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7222_ net316 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[6\]
+ vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7153_ net294 team_08_WB.instance_to_wrap.allocation.game.controller.state\[0\] vssd1
+ vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6104_ _2028_ _2055_ _2056_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__and3_1
X_7084_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[5\]
+ _2789_ _2799_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[5\]
+ _2826_ vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6035_ _1922_ _1947_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout283_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5841__A2 _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9546__414 vssd1 vssd1 vccd1 vccd1 _9546__414/HI net414 sky130_fd_sc_hd__conb_1
XANTENNA__7579__C1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7986_ _0422_ _0423_ vssd1 vssd1 vccd1 vccd1 _3524_ sky130_fd_sc_hd__nor2_2
XFILLER_0_95_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6937_ _2403_ _2721_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6868_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[7\]
+ _2675_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8543__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9587_ net451 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_92_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5776__A_N _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5819_ _1771_ _1770_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__and2b_1
X_8607_ _0695_ _4063_ vssd1 vssd1 vccd1 vccd1 _4086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6799_ net519 _2630_ net270 vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8538_ net163 _4012_ vssd1 vssd1 vccd1 vccd1 _4017_ sky130_fd_sc_hd__or2_1
X_9592__456 vssd1 vssd1 vccd1 vccd1 _9592__456/HI net456 sky130_fd_sc_hd__conb_1
XFILLER_0_5_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8469_ _3279_ _3894_ _3947_ _3949_ vssd1 vssd1 vccd1 vccd1 _3950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8638__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5062__B _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9486__361 vssd1 vssd1 vccd1 vccd1 _9486__361/HI net361 sky130_fd_sc_hd__conb_1
XFILLER_0_28_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7717__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8564__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7840_ net159 _3406_ _3407_ net165 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_19_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4983_ _0809_ _0927_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7771_ net149 net125 _3358_ _3360_ vssd1 vssd1 vccd1 vccd1 _3361_ sky130_fd_sc_hd__o211a_1
X_9510_ net385 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
X_6722_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ net268 _2580_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__and3b_1
XANTENNA__6812__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9441_ clknet_leaf_6_wb_clk_i _0386_ net211 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7627__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6653_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[3\] _2533_ _2532_
+ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[3\]
+ sky130_fd_sc_hd__mux2_1
X_5604_ net147 net145 vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout129_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9372_ clknet_leaf_24_wb_clk_i _0320_ net252 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6584_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[7\] _2488_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5535_ _1486_ _1487_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_83_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8323_ _3812_ _3813_ vssd1 vssd1 vccd1 vccd1 _3814_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5466_ _1416_ _1417_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8254_ net298 _3748_ _3750_ _3457_ vssd1 vssd1 vccd1 vccd1 _3751_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7205_ _2874_ _2906_ vssd1 vssd1 vccd1 vccd1 _2907_ sky130_fd_sc_hd__nor2_1
X_5397_ _0960_ _1197_ _0961_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__a21o_1
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_8
X_8185_ _3698_ _3700_ _3702_ net243 net568 vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__o32a_1
Xfanout302 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_2
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_4
Xfanout335 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[0\] vssd1
+ vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7136_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[16\]
+ _2856_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__xor2_1
XANTENNA_input3_A gpio_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7067_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[2\]
+ _2789_ _2792_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[2\]
+ _2812_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__a221o_1
X_6018_ _1967_ _1970_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6775__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7969_ _0487_ _3493_ vssd1 vssd1 vccd1 vccd1 _3508_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9639_ net264 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5057__B _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5750__A1 _0835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7553__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8384__A _3241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7728__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5248__A _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9575__440 vssd1 vssd1 vccd1 vccd1 _9575__440/HI net440 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5320_ _1223_ _1224_ _1220_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__a21o_1
X_5251_ _1157_ _1203_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5182_ _1077_ _1134_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8941_ _2322_ _2390_ vssd1 vssd1 vccd1 vccd1 _4418_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8872_ _4290_ _4298_ _4291_ vssd1 vssd1 vccd1 vccd1 _4350_ sky130_fd_sc_hd__o21ai_1
XANTENNA__6757__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7823_ _3395_ _3396_ _0457_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7754_ net174 _3343_ vssd1 vssd1 vccd1 vccd1 _3344_ sky130_fd_sc_hd__nor2_1
X_4966_ _0809_ _0916_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__nand2_8
X_6705_ _2568_ _2569_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout246_A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7357__B _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4897_ net138 _0849_ _0848_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__o21ai_4
XANTENNA__5980__A1 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7685_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[4\]
+ _3260_ _3254_ vssd1 vssd1 vccd1 vccd1 _3275_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9424_ clknet_leaf_43_wb_clk_i _0369_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_6636_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[27\] _2523_
+ vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__and2_1
X_9355_ clknet_leaf_27_wb_clk_i _0303_ net253 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4535__A2 team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6567_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _2480_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5518_ _1413_ _1414_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8306_ _3785_ _3787_ _3555_ vssd1 vssd1 vccd1 vccd1 _3798_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7373__A team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout201_X net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5605__B _0909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9286_ clknet_leaf_13_wb_clk_i _0129_ net214 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6498_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[1\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[2\] vssd1 vssd1
+ vccd1 vccd1 _2432_ sky130_fd_sc_hd__a21o_1
X_5449_ _1399_ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__and2_1
X_8237_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[18\]
+ _2995_ vssd1 vssd1 vccd1 vccd1 _3738_ sky130_fd_sc_hd__nand2_1
X_8168_ _0690_ _3627_ _0691_ vssd1 vssd1 vccd1 vccd1 _3687_ sky130_fd_sc_hd__o21a_1
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_2
XFILLER_0_11_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout110 _3235_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout132 _1075_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_4
Xfanout143 _0742_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_4
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_2
X_7119_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[10\]
+ _2848_ vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__xor2_2
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout198 net199 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlymetal6s2s_1
X_8099_ _0675_ _0686_ vssd1 vssd1 vccd1 vccd1 _3627_ sky130_fd_sc_hd__xnor2_2
Xfanout176 _3178_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_2
Xfanout187 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_4
XANTENNA__8491__X _3971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7548__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9332__RESET_B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9598__462 vssd1 vssd1 vccd1 vccd1 _9598__462/HI net462 sky130_fd_sc_hd__conb_1
XFILLER_0_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7715__A_N _3261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6279__A2 _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5487__B1 _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8826__B net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7779__A2 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8728__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6739__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8728__B2 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ _0760_ _0770_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__xnor2_4
XANTENNA__9073__RESET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6081__B _0926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9446__Q team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4751_ _0661_ net183 _0703_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4682_ net294 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoMovement team_08_WB.instance_to_wrap.allocation.game.controller.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_43_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7470_ net517 net115 _3111_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8900__A1 _3271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6421_ _2371_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__inv_2
X_9140_ clknet_leaf_38_wb_clk_i _0241_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6352_ _2303_ _2302_ _2299_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__or3b_1
X_5303_ _1039_ _1047_ _1255_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__a21o_1
X_6283_ _2103_ _2232_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9439__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9071_ clknet_leaf_49_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[1\]
+ net224 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5234_ net130 _1186_ _1184_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__a21o_1
X_8022_ _3481_ _3547_ _3558_ net241 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__o32a_1
X_5165_ _0943_ _1117_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout196_A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5096_ _0746_ _0765_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__or2_1
X_8924_ _0661_ net111 net183 vssd1 vssd1 vccd1 vccd1 _4401_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8855_ net321 _4329_ vssd1 vssd1 vccd1 vccd1 _4333_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7806_ _3386_ _3388_ vssd1 vssd1 vccd1 vccd1 _3389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5998_ _0918_ _1859_ _1858_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8786_ _4263_ vssd1 vssd1 vccd1 vccd1 _4264_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout151_X net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4949_ _0844_ _0874_ _0900_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__nor3_1
XFILLER_0_90_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7737_ _3320_ _3326_ _3317_ vssd1 vssd1 vccd1 vccd1 _3327_ sky130_fd_sc_hd__o21a_1
X_7668_ _3257_ vssd1 vssd1 vccd1 vccd1 _3258_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9407_ clknet_leaf_31_wb_clk_i _0354_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6619_ _2513_ net260 _2512_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[20\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_90_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7599_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[11\]
+ _3185_ _3180_ vssd1 vssd1 vccd1 vccd1 _3189_ sky130_fd_sc_hd__a21oi_1
X_9338_ clknet_leaf_33_wb_clk_i _0003_ net249 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_9269_ clknet_leaf_12_wb_clk_i _0078_ net220 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6433__A2 _2325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9526__401 vssd1 vssd1 vccd1 vccd1 _9526__401/HI net401 sky130_fd_sc_hd__conb_1
XFILLER_0_84_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8381__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7933__A2 _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8343__C1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5085__X _1038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8837__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8949__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8413__A3 _3355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6970_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[18\]
+ _2741_ vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__or2_1
X_5921_ _1870_ _1871_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_85_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5852_ _1757_ _1758_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8640_ net279 net173 vssd1 vssd1 vccd1 vccd1 _4119_ sky130_fd_sc_hd__nor2_1
X_5783_ _1735_ _1734_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4803_ net144 net167 vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8571_ net127 _3619_ _4049_ vssd1 vssd1 vccd1 vccd1 _4050_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7916__A team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4734_ _0658_ _0665_ _0669_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__o21a_2
X_7522_ _0437_ _3152_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8334__C1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4665_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[0\] vssd1
+ vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__nand2b_2
XANTENNA__4611__Y _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7453_ net303 _3043_ _3095_ _0438_ vssd1 vssd1 vccd1 vccd1 _3096_ sky130_fd_sc_hd__a211o_1
XANTENNA__5163__A2 _1088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6360__B2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6360__A1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7384_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[2\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _3033_ sky130_fd_sc_hd__or3b_1
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout111_A _3235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4596_ _0557_ _0558_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__nor2_1
X_6404_ team_08_WB.instance_to_wrap.allocation.game.game.score\[3\] _2338_ vssd1 vssd1
+ vccd1 vccd1 _2355_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6335_ _0663_ _0689_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9123_ clknet_leaf_40_wb_clk_i _0224_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9054_ clknet_leaf_35_wb_clk_i _0189_ net245 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6266_ _2082_ _2094_ _2111_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__and3_1
X_8005_ net326 net324 net319 vssd1 vssd1 vccd1 vccd1 _3542_ sky130_fd_sc_hd__and3_2
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6197_ _1191_ _1248_ _2148_ _1189_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__a31o_1
X_5217_ _1142_ _1158_ _1160_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout199_X net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5148_ _1096_ _1098_ _1099_ _0855_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5079_ _1030_ _1031_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__nor2_1
X_8907_ _2285_ net125 _4383_ vssd1 vssd1 vccd1 vccd1 _4384_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4515__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8838_ _4289_ _4304_ _4302_ _4301_ vssd1 vssd1 vccd1 vccd1 _4316_ sky130_fd_sc_hd__a211o_1
XANTENNA__7376__B1 _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7915__A2 _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8769_ net105 _4246_ vssd1 vssd1 vccd1 vccd1 _4247_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7385__X _3034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4450_ net653 vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6120_ net168 _0922_ _2072_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8095__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6051_ _1961_ _1963_ _1962_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__a21o_1
X_5002_ _0953_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6953_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[11\]
+ _2729_ _2731_ net157 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__o211a_1
X_5904_ _1807_ _1809_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6884_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__or4_1
X_5835_ _1744_ _1751_ _1752_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout159_A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8623_ net162 _4093_ _4101_ _0694_ vssd1 vssd1 vccd1 vccd1 _4102_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_17_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5766_ _1715_ _1717_ _1718_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout326_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8554_ _4020_ _4021_ _4023_ _4015_ _4032_ vssd1 vssd1 vccd1 vccd1 _4033_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5697_ _1603_ _1648_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8858__B1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4717_ _0670_ _0671_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__nand2_1
X_7505_ net306 _3044_ _3074_ _3089_ vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__o31ai_1
X_8485_ net191 net188 net185 vssd1 vssd1 vccd1 vccd1 _3965_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5166__A _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4648_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[7\] vssd1
+ vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7436_ _3045_ _3051_ _0440_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7367_ net296 net277 _3018_ vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__or3_1
X_4579_ net164 _0534_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__nor2_2
X_9106_ clknet_leaf_39_wb_clk_i _0209_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__7381__A team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8477__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6318_ net330 _2267_ _2269_ _2264_ _2268_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__o221a_1
X_7298_ _0644_ _2971_ vssd1 vssd1 vccd1 vccd1 _2972_ sky130_fd_sc_hd__nand2_2
X_6249_ _2125_ _2126_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__xor2_1
XANTENNA__4647__A1 _0602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9037_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[19\]
+ net210 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6725__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5072__A1 _0959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5804__A _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8387__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6619__B net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8834__B net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold90 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[2\]
+ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8552__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7466__A team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_dino vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5620_ net128 _1524_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5551_ _1453_ _1503_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4574__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4502_ _0469_ _0470_ _0471_ _0472_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__or4_1
X_8270_ net194 _3762_ _3764_ vssd1 vssd1 vccd1 vccd1 _3765_ sky130_fd_sc_hd__or3b_1
X_5482_ _1429_ _1433_ _1434_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__o21ai_2
X_7221_ net319 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__xor2_1
XANTENNA__8297__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7152_ net670 net37 net39 vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__and3b_1
XFILLER_0_67_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6103_ _2025_ _2027_ _2026_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__a21o_1
X_7083_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[5\]
+ _2792_ _2800_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6034_ _1984_ _1986_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout276_A _2547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7985_ _0485_ _3521_ _3522_ vssd1 vssd1 vccd1 vccd1 _3523_ sky130_fd_sc_hd__nor3_1
XFILLER_0_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6936_ net609 _2402_ net157 vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8760__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5448__X _1401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6867_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[7\]
+ _2675_ _2677_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9586_ net450 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5818_ _1722_ _1723_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6798_ _2630_ _2631_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8606_ _4065_ _4068_ _4072_ _4074_ _4084_ vssd1 vssd1 vccd1 vccd1 _4085_ sky130_fd_sc_hd__a221o_1
X_5749_ _1701_ _1700_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__nand2b_1
XANTENNA__4512__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8537_ net162 _4012_ vssd1 vssd1 vccd1 vccd1 _4016_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7649__A4 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8468_ _3354_ _3900_ _3948_ vssd1 vssd1 vccd1 vccd1 _3949_ sky130_fd_sc_hd__a21oi_1
X_7419_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_over team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_idle
+ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_win team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_cloud
+ vssd1 vssd1 vccd1 vccd1 _3064_ sky130_fd_sc_hd__or4_4
X_8399_ net116 net94 vssd1 vssd1 vccd1 vccd1 _3880_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8654__B net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7886__B1_N net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8670__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__5821__X _1774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4982_ _0924_ _0933_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7770_ net154 net135 vssd1 vssd1 vccd1 vccd1 _3360_ sky130_fd_sc_hd__nand2_2
XFILLER_0_92_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4795__A0 _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6721_ _2580_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_3_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9440_ clknet_leaf_5_wb_clk_i _0385_ net205 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_6652_ _0641_ _0647_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9371_ clknet_leaf_24_wb_clk_i _0319_ net252 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_5603_ _1511_ _1512_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_30_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8322_ _3553_ _3798_ _3811_ vssd1 vssd1 vccd1 vccd1 _3813_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_30_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6583_ net571 _2488_ _2490_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[7\]
+ sky130_fd_sc_hd__a21oi_1
X_5534_ _1430_ _1432_ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5465_ _1416_ _1417_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__and2b_1
XFILLER_0_83_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8253_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\] _0450_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[9\]
+ _0449_ _3749_ vssd1 vssd1 vccd1 vccd1 _3750_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9450__RESET_B net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7204_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[17\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[18\]
+ _2903_ vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8184_ _0702_ _3695_ _3701_ _2419_ vssd1 vssd1 vccd1 vccd1 _3702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5396_ _0766_ _0971_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__and2_1
Xfanout314 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[7\] vssd1
+ vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_4
Xfanout303 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_2
X_7135_ _2865_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__inv_2
Xfanout325 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[4\] vssd1
+ vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_4
XANTENNA__8755__A _3542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7066_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[2\]
+ _2800_ vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__and2_1
X_6017_ _1967_ _1968_ _1969_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7968_ _3503_ _3504_ _3506_ net170 vssd1 vssd1 vccd1 vccd1 _3507_ sky130_fd_sc_hd__a211o_1
XANTENNA__6562__X _2477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7899_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[19\]
+ net160 _3444_ vssd1 vssd1 vccd1 vccd1 _3449_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6722__B net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4786__B1 _0634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6919_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[10\]
+ _2709_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9638_ net486 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4523__A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9600__464 vssd1 vssd1 vccd1 vccd1 _9600__464/HI net464 sky130_fd_sc_hd__conb_1
X_9569_ net497 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
XFILLER_0_45_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8384__B _3864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6913__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7728__B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5250_ _0862_ _1156_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__or2_1
XANTENNA__8140__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5181_ net130 _1076_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8575__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_79_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8940_ _2296_ _3276_ _4416_ vssd1 vssd1 vccd1 vccd1 _4417_ sky130_fd_sc_hd__a21oi_1
XANTENNA__6454__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8871_ net103 _3544_ vssd1 vssd1 vccd1 vccd1 _4349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7822_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ _3395_ vssd1 vssd1 vccd1 vccd1 _3397_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4965_ _0810_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7753_ net126 _3290_ vssd1 vssd1 vccd1 vccd1 _3343_ sky130_fd_sc_hd__nor2_1
XANTENNA__5439__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6704_ net643 _2567_ net268 vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4896_ _0793_ _0813_ _0819_ net140 vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout239_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5980__A2 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9423_ clknet_leaf_42_wb_clk_i _0368_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7684_ net185 net97 _3273_ net100 vssd1 vssd1 vccd1 vccd1 _3274_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6635_ _2523_ net260 _2522_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[26\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_13_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9354_ clknet_leaf_26_wb_clk_i _0302_ net249 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6566_ net262 _2473_ _2479_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[1\]
+ sky130_fd_sc_hd__and3_1
X_5517_ _0807_ _1457_ _1469_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__a21oi_1
X_9285_ clknet_leaf_14_wb_clk_i _0128_ net213 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_8305_ _3784_ _3796_ _3797_ net230 net612 vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__o32a_1
XFILLER_0_6_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8131__B1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8236_ _3727_ _3737_ _3711_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__o21a_1
X_6497_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[1\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[2\] vssd1 vssd1
+ vccd1 vccd1 _2431_ sky130_fd_sc_hd__and3_1
X_5448_ _1352_ _1400_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5379_ _1330_ _1331_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__or2_1
X_8167_ net613 net243 _3686_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__o21ba_1
Xfanout122 _3001_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_2
Xfanout100 _3265_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_4
Xfanout111 _3235_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_2
Xfanout144 _0739_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_4
X_8098_ net620 net243 _3620_ _3626_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__o22a_1
X_7118_ _2848_ _2849_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__nor2_1
Xfanout155 _3186_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_4
Xfanout133 net134 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
Xfanout166 _3402_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
Xfanout199 _3459_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
X_7049_ _2787_ _2791_ net293 vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__o21a_1
Xfanout188 net190 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
Xfanout177 _3178_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9372__RESET_B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4513__A_N team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7564__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9301__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8379__B net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9535__491 vssd1 vssd1 vccd1 vccd1 net491 _9535__491/LO sky130_fd_sc_hd__conb_1
XANTENNA__8425__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6627__B net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6436__B1 _2325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7739__A _3265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4750_ _0661_ net183 vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4681_ _0637_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.reset
+ sky130_fd_sc_hd__inv_2
XFILLER_0_71_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6420_ _2333_ _2369_ _2370_ _2335_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__a2bb2o_2
X_6351_ net325 _2301_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5302_ _1252_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6282_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[0\]
+ _0716_ _0917_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__or3_1
X_9070_ clknet_leaf_49_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[0\]
+ net224 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5233_ _1184_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8021_ net322 _2426_ _3557_ net300 _3016_ vssd1 vssd1 vccd1 vccd1 _3558_ sky130_fd_sc_hd__a221o_1
X_5164_ net123 _1116_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__xor2_1
X_5095_ _0746_ _0765_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout189_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8923_ _0661_ net111 _4395_ _4399_ vssd1 vssd1 vccd1 vccd1 _4400_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8854_ _4330_ _4331_ vssd1 vssd1 vccd1 vccd1 _4332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7805_ _2972_ _3387_ vssd1 vssd1 vccd1 vccd1 _3388_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5997_ _1949_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8785_ _0521_ _4262_ vssd1 vssd1 vccd1 vccd1 _4263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4948_ _0844_ _0874_ _0900_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout144_X net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7736_ _3294_ _3307_ _3325_ _3323_ vssd1 vssd1 vccd1 vccd1 _3326_ sky130_fd_sc_hd__o31a_1
XFILLER_0_90_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4879_ _0831_ _0807_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__and2b_1
X_7667_ _3238_ _3256_ vssd1 vssd1 vccd1 vccd1 _3257_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9406_ clknet_leaf_31_wb_clk_i _0353_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_6618_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[19\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[20\]
+ _2509_ vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7598_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[11\]
+ _3180_ net150 vssd1 vssd1 vccd1 vccd1 _3188_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9337_ clknet_leaf_26_wb_clk_i _0002_ net249 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6549_ _2464_ _2465_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[19\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__7671__X _3261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9268_ clknet_leaf_12_wb_clk_i _0090_ net220 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9199_ clknet_leaf_16_wb_clk_i _0033_ net221 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6728__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8219_ _2990_ _3725_ net121 vssd1 vssd1 vccd1 vccd1 _3726_ sky130_fd_sc_hd__a21o_1
XANTENNA__8943__A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7091__B1 _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7559__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9606__470 vssd1 vssd1 vccd1 vccd1 _9606__470/HI net470 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_26_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4904__B1 _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5261__B _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5920_ _0918_ _1766_ _1765_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__a21bo_1
XANTENNA__6373__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5851_ _1801_ _1803_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9294__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5782_ _1678_ _1684_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__xnor2_1
X_4802_ net167 vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8570_ net136 _4041_ _4046_ _4048_ vssd1 vssd1 vccd1 vccd1 _4049_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7916__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4733_ _0675_ _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__nor2_1
X_7521_ _3151_ _3152_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7452_ net305 _3042_ _3044_ _3080_ _0437_ vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__o311a_1
XFILLER_0_12_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5699__A1 _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4664_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[1\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[1\] vssd1
+ vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__and2b_1
XANTENNA__8885__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6403_ _2329_ _2353_ _2352_ _2334_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__8885__B2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7383_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[2\] team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__or2_1
X_4595_ net191 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ net188 vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6334_ _2285_ vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__inv_2
X_9122_ clknet_leaf_42_wb_clk_i _0223_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA_fanout104_A _3272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6265_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[7\]
+ _2217_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__nor2_1
X_9053_ clknet_leaf_35_wb_clk_i _0188_ net245 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_5216_ _1167_ _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__or2_1
XANTENNA__5452__A _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8004_ net320 _3524_ vssd1 vssd1 vccd1 vccd1 _3541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6196_ _1191_ _1248_ _2148_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__and3_1
X_5147_ _0855_ _1099_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__nand2_1
XANTENNA__8763__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5078_ _1027_ _1028_ _1029_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8906_ net134 _3627_ _4380_ _4382_ vssd1 vssd1 vccd1 vccd1 _4383_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4515__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8837_ net100 _4314_ vssd1 vssd1 vccd1 vccd1 _4315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8768_ _4232_ _4245_ vssd1 vssd1 vccd1 vccd1 _4246_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7719_ net175 _3300_ vssd1 vssd1 vccd1 vccd1 _3309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8699_ _2386_ _4177_ vssd1 vssd1 vccd1 vccd1 _4178_ sky130_fd_sc_hd__or2_1
XANTENNA__6336__C1 _0685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8876__B2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5914__X _1867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9636__485 vssd1 vssd1 vccd1 vccd1 _9636__485/HI net485 sky130_fd_sc_hd__conb_1
XFILLER_0_31_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6639__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input34_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4851__A_N _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6921__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5537__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8867__B2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6050_ _2000_ _2001_ _1999_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__a21bo_1
X_5001_ net123 _0952_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__nand2_1
XANTENNA__8583__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6374__Y _2325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6952_ _2730_ vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5903_ _1852_ _1855_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6883_ net520 _2685_ _2687_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7358__A1 _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5834_ _1785_ _1786_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8622_ _0686_ _4095_ _4100_ vssd1 vssd1 vccd1 vccd1 _4101_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7646__B net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5765_ _0923_ _1668_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8553_ _4031_ _4024_ _4015_ vssd1 vssd1 vccd1 vccd1 _4032_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout221_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5696_ net147 _0906_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4716_ net288 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout319_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7504_ net525 net114 _3121_ _3141_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__o22a_1
X_8484_ _3890_ _3956_ _3963_ _3960_ _3958_ vssd1 vssd1 vccd1 vccd1 _3964_ sky130_fd_sc_hd__a32o_1
X_4647_ _0602_ _0603_ _0573_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__a21o_2
X_7435_ _0440_ _3078_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_15_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7366_ _2427_ _3017_ vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4578_ _0489_ _0492_ _0494_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__and3_1
X_6317_ net335 _0450_ _0451_ net333 vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9105_ clknet_leaf_43_wb_clk_i _0208_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout107_X net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8477__B _3284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7297_ net283 team_08_WB.instance_to_wrap.allocation.game.cactusMove.drawDoneCactus
+ net262 _2323_ vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__and4_1
XANTENNA__8653__A_N _3261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6248_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[16\]
+ _2200_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__nor2_1
X_9036_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[18\]
+ net207 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8589__A1_N net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6179_ _1642_ _2131_ _1640_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4813__X _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_33_Left_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5804__B _0926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold91 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[7\]
+ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[3\]
+ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6635__B net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7466__B _3064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5550_ _0747_ _1452_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4501_ net9 net8 net11 net10 vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__or4_1
X_5481_ _1384_ _1385_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7220_ _2912_ _2913_ _2917_ _2918_ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__or4_1
XANTENNA__8297__B _3776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8068__A2 _0702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7151_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.internalSck
+ net3 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.cs vssd1 vssd1
+ vccd1 vccd1 net66 sky130_fd_sc_hd__and3_1
X_9470__345 vssd1 vssd1 vccd1 vccd1 _9470__345/HI net345 sky130_fd_sc_hd__conb_1
X_6102_ _2051_ _2054_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7082_ team_08_WB.instance_to_wrap.allocation.game.controller.color\[11\] _2796_
+ _2809_ team_08_WB.instance_to_wrap.allocation.game.controller.color\[10\] vssd1
+ vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6033_ _1984_ _1985_ _1980_ vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__or3b_1
X_9511__386 vssd1 vssd1 vccd1 vccd1 _9511__386/HI net386 sky130_fd_sc_hd__conb_1
X_7984_ _0488_ _0493_ vssd1 vssd1 vccd1 vccd1 _3522_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6935_ _2402_ _2720_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout269_A _2548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7594__A4 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8956__A2_N _3214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6866_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[7\]
+ _2675_ net273 vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__a21oi_1
X_9585_ net449 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5817_ _1753_ _1754_ _1769_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__a21o_1
X_6797_ net632 _2629_ net270 vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8605_ _4078_ _4081_ _4083_ vssd1 vssd1 vccd1 vccd1 _4084_ sky130_fd_sc_hd__a21oi_1
XANTENNA__7751__A1 _3284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5748_ _0835_ _1695_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout224_X net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8536_ net127 _3685_ _4014_ net136 vssd1 vssd1 vccd1 vccd1 _4015_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5679_ _1630_ _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8467_ _3279_ _3901_ _3916_ _3880_ _3882_ vssd1 vssd1 vccd1 vccd1 _3948_ sky130_fd_sc_hd__o2111a_1
X_7418_ _3053_ _3062_ _3022_ vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8398_ net110 _3865_ vssd1 vssd1 vccd1 vccd1 _3879_ sky130_fd_sc_hd__nand2_1
X_7349_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr1\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusDist.lfsr2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8059__A2 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9019_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[1\]
+ net208 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5640__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9326__RESET_B net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5045__A2 _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7423__A_N team_08_WB.instance_to_wrap.allocation.game.lcdOutput.r_dino vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8519__B1 _2325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7742__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8398__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_75_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5550__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8758__B1 _0425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4981_ _0924_ _0933_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6720_ _2577_ _2578_ _2579_ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6651_ _0641_ _0647_ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__nor2_1
X_5602_ _1087_ _1554_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__nand2_1
X_9370_ clknet_leaf_24_wb_clk_i _0318_ net252 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_6582_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[7\] _2488_ _2478_
+ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5533_ _1483_ _1485_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__nor2_1
X_8321_ _3553_ _3798_ _3811_ vssd1 vssd1 vccd1 vccd1 _3812_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5464_ _1367_ _1368_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_78_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8252_ _0551_ net195 _3747_ _0463_ vssd1 vssd1 vccd1 vccd1 _3749_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5395_ _1343_ _1345_ _1346_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9552__420 vssd1 vssd1 vccd1 vccd1 _9552__420/HI net420 sky130_fd_sc_hd__conb_1
X_7203_ _2904_ _2905_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__nor2_1
X_8183_ net163 _0709_ vssd1 vssd1 vccd1 vccd1 _3701_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7940__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout304 net306 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_2
XFILLER_0_2_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7134_ _2857_ _2859_ _2864_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__and3_1
Xfanout326 net328 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
Xfanout315 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[7\] vssd1
+ vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
X_7065_ _2808_ _2810_ _2811_ _2806_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__o31a_1
X_6016_ _1927_ _1966_ _1965_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__a21o_1
XANTENNA__8771__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7967_ net327 _3487_ _3505_ net196 vssd1 vssd1 vccd1 vccd1 _3506_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_49_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7898_ _3447_ _3448_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__and2_1
X_6918_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[10\]
+ _2709_ _2711_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__o21a_1
X_9637_ net266 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6849_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ net269 _2665_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__and3b_1
XANTENNA__4523__B team_08_WB.instance_to_wrap.allocation.game.controller.v\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9568_ net496 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_0_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8519_ _3972_ _3993_ _3998_ _2325_ net210 vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__o311a_1
X_9499_ net374 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__8011__A team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8946__A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8665__B _3608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6999__C1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7728__C _3305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8140__A1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8856__A _3789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5180_ net131 _1132_ _1130_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__a21o_1
XANTENNA__6454__A1 _0419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8870_ _4234_ _4347_ vssd1 vssd1 vccd1 vccd1 _4348_ sky130_fd_sc_hd__nand2_1
X_9582__446 vssd1 vssd1 vccd1 vccd1 _9582__446/HI net446 sky130_fd_sc_hd__conb_1
XFILLER_0_94_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7821_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\]
+ _3395_ vssd1 vssd1 vccd1 vccd1 _3396_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4964_ _0623_ _0726_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_35_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7752_ _3288_ _3290_ _3294_ _3306_ _3298_ vssd1 vssd1 vccd1 vccd1 _3342_ sky130_fd_sc_hd__o41a_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6703_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[9\]
+ _2567_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4895_ net140 net138 vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8903__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9422_ clknet_leaf_42_wb_clk_i _0367_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7683_ _3254_ _3262_ _3270_ vssd1 vssd1 vccd1 vccd1 _3273_ sky130_fd_sc_hd__and3_1
XANTENNA__5717__B1 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6634_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[25\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[26\]
+ _2519_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9353_ clknet_leaf_26_wb_clk_i _0301_ net249 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6565_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[1\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5516_ _1460_ _1467_ _1468_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__a21oi_1
X_9284_ clknet_leaf_13_wb_clk_i _0127_ net213 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_8304_ net297 _3791_ _3795_ net300 vssd1 vssd1 vccd1 vccd1 _3797_ sky130_fd_sc_hd__a22o_1
X_9476__351 vssd1 vssd1 vccd1 vccd1 _9476__351/HI net351 sky130_fd_sc_hd__conb_1
X_6496_ _0506_ _2428_ _2430_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[1\]
+ sky130_fd_sc_hd__and3_1
X_5447_ _1349_ _1351_ _1350_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__o21ai_1
X_8235_ _2994_ _3736_ net122 vssd1 vssd1 vccd1 vccd1 _3737_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8766__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5378_ _1322_ _1324_ _1329_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__nor3_1
X_8166_ _2286_ net137 _3685_ _0701_ _3682_ vssd1 vssd1 vccd1 vccd1 _3686_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9517__392 vssd1 vssd1 vccd1 vccd1 _9517__392/HI net392 sky130_fd_sc_hd__conb_1
Xfanout101 _3277_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_4
Xfanout112 _3234_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_4
Xfanout123 _0945_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_4
Xfanout145 _0908_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_4
X_8097_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\] _3614_ _3615_
+ _3625_ vssd1 vssd1 vccd1 vccd1 _3626_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7117_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[9\]
+ _2846_ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__nor2_1
Xfanout156 _2428_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_2
Xfanout134 _3201_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_4
Xfanout167 _0754_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_4
X_7048_ _2794_ _2795_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__nor2_1
Xfanout178 _0674_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
Xfanout189 net190 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_97_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5189__X _1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8999_ clknet_leaf_3_wb_clk_i _0163_ net203 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6436__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7298__Y _2972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7739__B _3276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6643__B net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4680_ net4 net1 team_08_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__or3b_4
XANTENNA__8897__C1 _3284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4922__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6350_ net321 _2296_ _2301_ net325 vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5301_ _0850_ _1253_ _1040_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6281_ net182 _0917_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8586__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5232_ _1178_ _1182_ _1183_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__and3_1
X_8020_ net322 net195 _3472_ _3556_ vssd1 vssd1 vccd1 vccd1 _3557_ sky130_fd_sc_hd__a211o_1
XANTENNA__9011__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5163_ _1087_ _1088_ _1106_ _1108_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__a31oi_2
X_5094_ _1045_ _1046_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__nor2_2
XANTENNA__4906__X _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8922_ _0660_ net113 _4397_ _4398_ vssd1 vssd1 vccd1 vccd1 _4399_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8853_ net321 _4329_ net317 vssd1 vssd1 vccd1 vccd1 _4331_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5938__B1 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7804_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr1\[0\] team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3387_ sky130_fd_sc_hd__xor2_2
XANTENNA_fanout251_A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5996_ _1881_ _1913_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8784_ net325 _4261_ vssd1 vssd1 vccd1 vccd1 _4262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4947_ _0881_ _0898_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7735_ net108 net106 _3261_ net110 vssd1 vssd1 vccd1 vccd1 _3325_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4878_ _0745_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7666_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[6\]
+ net108 _3255_ vssd1 vssd1 vccd1 vccd1 _3256_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9405_ clknet_leaf_30_wb_clk_i _0352_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6617_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[19\] _2509_
+ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[20\] vssd1 vssd1 vccd1
+ vccd1 _2512_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9336_ clknet_leaf_32_wb_clk_i _0001_ net249 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_41_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7597_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\]
+ _3182_ _3185_ vssd1 vssd1 vccd1 vccd1 _3187_ sky130_fd_sc_hd__a21o_1
X_6548_ net644 _2462_ net156 vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__o21ai_1
X_9267_ clknet_leaf_12_wb_clk_i _0089_ net219 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_6479_ net137 vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9198_ clknet_leaf_16_wb_clk_i _0032_ net221 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_8218_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[10\]
+ _2989_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[11\]
+ vssd1 vssd1 vccd1 vccd1 _3725_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5191__Y _1144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4529__A _0423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8149_ _0663_ _0702_ _2393_ _2534_ vssd1 vssd1 vccd1 vccd1 _3671_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7918__A1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8343__A1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4551__X _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5095__A _0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7469__B _3110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4445__Y _0419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6373__B _2324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5850_ net142 _0927_ _1801_ _1802_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__nand4_1
XFILLER_0_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5781_ _1726_ _1731_ _1732_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4801_ _0721_ _0752_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_57_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4902__A _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7916__C net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4732_ net162 net169 vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__nand2_1
X_7520_ net305 _3040_ _3054_ vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4663_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7451_ net308 _3093_ _3091_ net305 vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5699__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6402_ team_08_WB.instance_to_wrap.allocation.game.game.score\[4\] _2328_ _2347_
+ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7382_ _3030_ _3031_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__or2_1
X_4594_ _0425_ _0557_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__xnor2_1
XANTENNA__6829__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9121_ clknet_leaf_30_wb_clk_i _0222_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.color\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_6333_ _0675_ _0708_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6264_ _2113_ _2114_ vssd1 vssd1 vccd1 vccd1 _2217_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9052_ clknet_leaf_34_wb_clk_i _0187_ net246 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_5215_ _1164_ _1166_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8003_ net170 net297 vssd1 vssd1 vccd1 vccd1 _3540_ sky130_fd_sc_hd__and2b_1
X_6195_ _1302_ _2146_ _1249_ _1300_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout299_A team_08_WB.instance_to_wrap.allocation.game.controller.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9588__452 vssd1 vssd1 vccd1 vccd1 _9588__452/HI net452 sky130_fd_sc_hd__conb_1
X_5146_ _0852_ _0854_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__or2_1
X_5077_ _1027_ _1028_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__nor3_1
X_8905_ net155 _3642_ _4381_ vssd1 vssd1 vccd1 vccd1 _4382_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8482__C _3284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout254_X net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8836_ _4198_ _4313_ vssd1 vssd1 vccd1 vccd1 _4314_ sky130_fd_sc_hd__or2_1
XANTENNA__7376__A2 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5979_ _1928_ _1929_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4653__A_N team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8767_ _0423_ _4212_ vssd1 vssd1 vccd1 vccd1 _4245_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_23_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7718_ _3300_ _3302_ vssd1 vssd1 vccd1 vccd1 _3308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8698_ net286 net285 net281 vssd1 vssd1 vccd1 vccd1 _4177_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8003__B net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7649_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[7\]
+ _3217_ _3227_ net110 _3229_ vssd1 vssd1 vccd1 vccd1 _3239_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_91_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9319_ clknet_leaf_29_wb_clk_i _0289_ net233 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8261__B1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7603__A3 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8316__A1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6649__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5000_ net123 _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__or2_1
XANTENNA__6655__Y _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6951_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[9\]
+ _2725_ vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5902_ _1852_ _1854_ _1853_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__or3b_1
XFILLER_0_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6882_ net520 _2685_ net269 vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__o21ai_1
X_5833_ _1074_ _1737_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4903__Y _0856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9444__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8621_ _4093_ _4096_ _4097_ vssd1 vssd1 vccd1 vccd1 _4100_ sky130_fd_sc_hd__nand3_1
XFILLER_0_91_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8552_ _0663_ net113 _4009_ _4025_ _4030_ vssd1 vssd1 vccd1 vccd1 _4031_ sky130_fd_sc_hd__o311a_1
XFILLER_0_5_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5764_ _0923_ _1716_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__nand2_1
X_7503_ _3135_ _3139_ _3140_ net114 vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_16_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5695_ _0761_ _0910_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4715_ net288 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__nand2_1
X_8483_ _3280_ _3961_ _3962_ vssd1 vssd1 vccd1 vccd1 _3963_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4646_ _0573_ _0603_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7434_ _3045_ _3051_ net310 vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7365_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[1\] net296 vssd1
+ vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__or2_1
X_4577_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.state\[0\] _0544_
+ net290 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[5\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6316_ net335 net333 vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__or2_2
X_9104_ clknet_leaf_43_wb_clk_i _0207_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_7296_ net538 _2968_ _2970_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__a21oi_1
X_6247_ _2127_ _2128_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9035_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[17\]
+ net209 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8774__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6178_ _1693_ _2130_ _1691_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5129_ net130 _1080_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8819_ _0421_ net192 _4296_ net334 vssd1 vssd1 vccd1 vccd1 _4297_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_36_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7506__C1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold92 team_08_WB.instance_to_wrap.allocation.game.controller.state\[3\] vssd1 vssd1
+ vccd1 vccd1 net590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[7\]
+ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[21\]
+ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8859__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4500_ net36 net35 net7 net6 vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__or4_1
X_5480_ _1432_ _1430_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7763__A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_1 _3613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7150_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.cs net3 vssd1
+ vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__and2b_1
X_6101_ _2051_ _2052_ _2053_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__nand3_1
XFILLER_0_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7081_ _2778_ _2806_ _2823_ _2824_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__o22a_1
X_6032_ _1946_ _1957_ _1983_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__a21oi_1
X_7983_ _3493_ _3520_ vssd1 vssd1 vccd1 vccd1 _3521_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4914__X _0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6934_ net667 _2401_ net157 vssd1 vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_1_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5458__A _0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6865_ _2675_ _2676_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__nor2_1
X_8604_ net116 _4077_ _4082_ _4072_ vssd1 vssd1 vccd1 vccd1 _4083_ sky130_fd_sc_hd__a211o_1
X_9584_ net448 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_91_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5816_ _1767_ _1768_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__and2b_1
X_6796_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[12\]
+ _2629_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5747_ net167 _0910_ _1647_ _1699_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__o31ai_2
X_8535_ _4012_ _4013_ vssd1 vssd1 vccd1 vccd1 _4014_ sky130_fd_sc_hd__nor2_1
XANTENNA__8769__A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8466_ _3924_ _3943_ _3946_ _3907_ vssd1 vssd1 vccd1 vccd1 _3947_ sky130_fd_sc_hd__a31o_1
X_5678_ _1597_ _1628_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5464__Y _1417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7417_ net309 _3024_ _3058_ _3061_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__o2111a_1
XANTENNA__8700__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5193__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4629_ _0585_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8397_ _3876_ _3877_ _3874_ vssd1 vssd1 vccd1 vccd1 _3878_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7348_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[22\]
+ _2999_ net503 vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__o21a_1
X_7279_ net180 _2957_ _2959_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5817__A2 _1754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9018_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[0\]
+ net207 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4808__Y _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7019__A1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4789__C1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7742__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5753__A1 _1012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5815__B _1754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9493__368 vssd1 vssd1 vccd1 vccd1 _9493__368/HI net368 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_58_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_37_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4980_ _0927_ _0932_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6650_ _0426_ _2532_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_pixel\[2\]
+ sky130_fd_sc_hd__xnor2_1
X_5601_ _1514_ _1515_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6581_ _2488_ _2489_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5532_ _1476_ _1479_ _1483_ _1484_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_82_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4910__A _0810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8320_ _3548_ _3574_ vssd1 vssd1 vccd1 vccd1 _3811_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7497__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5463_ _0882_ _1410_ _1415_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__a21oi_1
X_8251_ _0552_ net195 _3472_ _3747_ vssd1 vssd1 vccd1 vccd1 _3748_ sky130_fd_sc_hd__a211o_1
X_5394_ _1343_ _1345_ _1346_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7202_ net693 _2903_ _2875_ vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__o21ai_1
X_8182_ _0651_ _3699_ _0654_ vssd1 vssd1 vccd1 vccd1 _3700_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7940__B net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_2
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7133_ _2862_ _2863_ _2861_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__a21o_1
XANTENNA__6837__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_4
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_4
X_7064_ _2780_ _2788_ _2797_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6015_ _0773_ _0921_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout281_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7939__Y _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4644__X _0602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7957__C1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout167_X net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7966_ net327 _3487_ vssd1 vssd1 vccd1 vccd1 _3505_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7897_ net160 _3444_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[19\]
+ vssd1 vssd1 vccd1 vccd1 _3448_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6917_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[10\]
+ _2709_ net272 vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__a21oi_1
X_9636_ net485 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6848_ _2665_ vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9567_ net435 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
X_6779_ net274 _2618_ _2619_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__nor3_1
XFILLER_0_18_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8518_ _3955_ _3964_ _3986_ _3274_ _3997_ vssd1 vssd1 vccd1 vccd1 _3998_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9498_ net373 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_33_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8011__B _3543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__7488__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8449_ net175 net124 _3359_ vssd1 vssd1 vccd1 vccd1 _3930_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4819__X _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5651__A _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9391__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6999__B1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8452__A3 _3888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5098__A _1012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6151__A1 _0723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9288__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4448__Y _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6454__A2 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7820_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\] _3393_
+ _3394_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.init_done
+ vssd1 vssd1 vccd1 vccd1 _3395_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4963_ _0623_ _0726_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_35_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7751_ _3284_ _3339_ _3340_ vssd1 vssd1 vccd1 vccd1 _3341_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_80_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6702_ net276 _2566_ _2567_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__nor3_1
XFILLER_0_50_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7682_ _3262_ _3270_ vssd1 vssd1 vccd1 vccd1 _3272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4894_ _0846_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6633_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[25\] team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[24\]
+ _2518_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[26\] vssd1
+ vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__a31o_1
X_9421_ clknet_leaf_41_wb_clk_i _0366_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9352_ clknet_leaf_27_wb_clk_i _0300_ net251 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__6331__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6564_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[0\] _2478_ vssd1
+ vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[0\]
+ sky130_fd_sc_hd__and2b_1
XANTENNA__7654__C net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout127_A _3214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5455__B _1407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5515_ _0807_ _1457_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9283_ clknet_leaf_14_wb_clk_i _0126_ net213 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_8303_ _2301_ net161 _2425_ _3527_ _3636_ vssd1 vssd1 vccd1 vccd1 _3796_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_14_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6495_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[1\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2430_ sky130_fd_sc_hd__nand2_1
X_5446_ _0885_ _1396_ _1398_ _0837_ _0769_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8234_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[16\]
+ _2993_ vssd1 vssd1 vccd1 vccd1 _3736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7890__B2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5377_ _1322_ _1324_ _1329_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__o21a_1
Xfanout102 _3277_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_2
X_8165_ _3683_ _3684_ vssd1 vssd1 vccd1 vccd1 _3685_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout113 _3234_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_2
Xfanout146 _0908_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_1
X_8096_ net299 _3622_ _3623_ _3624_ _3597_ vssd1 vssd1 vccd1 vccd1 _3625_ sky130_fd_sc_hd__a221o_1
X_7116_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[9\]
+ _2846_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__and2_1
Xfanout124 net125 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input1_A gpio_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout168 _0723_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_4
X_7047_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[2\] vssd1
+ vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__nand2_1
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
XANTENNA__8782__A _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout179 net181 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8998_ clknet_leaf_3_wb_clk_i _0162_ net202 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9386__Q team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7949_ net199 _3485_ _3487_ _3488_ vssd1 vssd1 vccd1 vccd1 _3489_ sky130_fd_sc_hd__a22o_1
XANTENNA__8006__B _3542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9559__427 vssd1 vssd1 vccd1 vccd1 _9559__427/HI net427 sky130_fd_sc_hd__conb_1
X_9619_ net264 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_98_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4550__A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7881__B2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4731__Y _0686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4460__A team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9499__374 vssd1 vssd1 vccd1 vccd1 _9499__374/HI net374 sky130_fd_sc_hd__conb_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4922__A2 _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5300_ _0852_ _0862_ _0815_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8113__A2 _3637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6280_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[1\]
+ _2103_ _2232_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5231_ _1178_ _1182_ _1183_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5162_ _1113_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__nand2b_1
X_5093_ _1044_ _0846_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__and2b_1
X_8921_ net183 net118 vssd1 vssd1 vccd1 vccd1 _4398_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8852_ _0520_ _4329_ vssd1 vssd1 vccd1 vccd1 _4330_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5938__A1 _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7803_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr1\[1\] team_08_WB.instance_to_wrap.allocation.game.cactus2size.lfsr2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3386_ sky130_fd_sc_hd__xnor2_1
X_8783_ _0422_ _3486_ vssd1 vssd1 vccd1 vccd1 _4261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5995_ _1922_ _1947_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__and2b_1
XANTENNA__5938__B2 _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7734_ _3323_ vssd1 vssd1 vccd1 vccd1 _3324_ sky130_fd_sc_hd__inv_2
X_4946_ _0881_ _0898_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_75_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4610__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout244_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4877_ _0828_ _0829_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7665_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[6\]
+ net108 net106 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[5\]
+ vssd1 vssd1 vccd1 vccd1 _3255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9404_ clknet_leaf_31_wb_clk_i _0351_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6363__A1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6616_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[19\] _2509_
+ _2511_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[19\]
+ sky130_fd_sc_hd__o21a_1
X_7596_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\]
+ _3182_ _3185_ vssd1 vssd1 vccd1 vccd1 _3186_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6547_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[19\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[18\]
+ _2461_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__and3_1
X_9335_ clknet_leaf_0_wb_clk_i _0018_ net201 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9266_ clknet_leaf_12_wb_clk_i _0088_ net219 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6478_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\] _0711_ vssd1
+ vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5429_ _1332_ _1334_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__and2_1
X_9197_ clknet_leaf_16_wb_clk_i _0031_ net221 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_8217_ net121 _3724_ _3036_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8148_ net299 _0653_ _2533_ _3597_ vssd1 vssd1 vccd1 vccd1 _3670_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4529__B net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8079_ _0642_ _2535_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[9\]
+ vssd1 vssd1 vccd1 vccd1 _3609_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7091__A2 _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4545__A _0419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7530__S team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4455__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4800_ _0721_ _0752_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__and2_2
XFILLER_0_57_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5780_ _1731_ _1732_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4731_ _0678_ _0679_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4662_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[2\] vssd1
+ vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__nand2b_1
X_7450_ _3050_ _3092_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7772__Y _3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6401_ team_08_WB.instance_to_wrap.allocation.game.game.score\[4\] _2343_ vssd1 vssd1
+ vccd1 vccd1 _2352_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9120_ clknet_leaf_31_wb_clk_i _0221_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.color\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7381_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\] _3028_
+ vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4593_ net191 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ net188 vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6332_ net318 _2279_ _2281_ net321 vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__o2bb2a_1
X_6263_ _2117_ _2215_ vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__or2_1
X_9051_ clknet_leaf_35_wb_clk_i _0186_ net245 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5214_ _1164_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8002_ _0483_ _0498_ _3516_ net196 vssd1 vssd1 vccd1 vccd1 _3539_ sky130_fd_sc_hd__o31a_1
X_6194_ _1302_ _2146_ _1300_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5145_ _0867_ _1097_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout194_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5076_ _0914_ _0940_ _0944_ net138 vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__o22a_1
XANTENNA__5084__A1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8904_ _0698_ _3178_ vssd1 vssd1 vccd1 vccd1 _4381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8022__B2 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8835_ net314 _0520_ vssd1 vssd1 vccd1 vccd1 _4313_ sky130_fd_sc_hd__nor2_1
X_5978_ net148 _0922_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8766_ net103 _4243_ vssd1 vssd1 vccd1 vccd1 _4244_ sky130_fd_sc_hd__xnor2_1
X_4929_ _0824_ _0826_ _0828_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_43_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7717_ net149 net135 vssd1 vssd1 vccd1 vccd1 _3307_ sky130_fd_sc_hd__nand2_2
X_8697_ net176 _4175_ vssd1 vssd1 vccd1 vccd1 _4176_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6336__A1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7648_ _0454_ _3233_ _3236_ vssd1 vssd1 vccd1 vccd1 _3238_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_62_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7682__Y _3272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7579_ team_08_WB.instance_to_wrap.allocation.game.game.score\[0\] _2347_ _3175_
+ _2335_ net255 vssd1 vssd1 vccd1 vccd1 _3176_ sky130_fd_sc_hd__a221o_1
X_9318_ clknet_leaf_23_wb_clk_i _0020_ _0152_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9249_ clknet_leaf_15_wb_clk_i _0100_ net214 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4546__Y _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8970__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9325__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6489__X _2426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7525__S team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6649__B _2477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7055__A2 _2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8252__A1 _0551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6950_ _2729_ net157 _2728_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__and3b_1
XFILLER_0_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5901_ _1803_ _1851_ _1850_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6881_ _2685_ _2686_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__nor2_1
X_5832_ _1781_ _1784_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__nor2_1
XANTENNA__4913__A _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8620_ _4094_ _4095_ _4098_ _4092_ vssd1 vssd1 vccd1 vccd1 _4099_ sky130_fd_sc_hd__o31a_1
X_5763_ _1713_ _1714_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4577__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8960__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8551_ _4011_ _4029_ vssd1 vssd1 vccd1 vccd1 _4030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4714_ _0658_ net183 vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__nand2_1
X_7502_ net304 net308 _3048_ _3125_ net301 vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__o311a_1
X_5694_ _0761_ net146 vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_44_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8482_ net189 _3278_ _3284_ vssd1 vssd1 vccd1 vccd1 _3962_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4645_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[8\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[8\] vssd1
+ vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__nand2b_1
X_7433_ net305 _3073_ _3076_ vssd1 vssd1 vccd1 vccd1 _3077_ sky130_fd_sc_hd__a21o_1
XANTENNA__5744__A _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7364_ net556 net242 _3016_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__o21a_1
X_4576_ net319 _0541_ _0543_ _0503_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__o2bb2a_1
X_6315_ _2265_ _2266_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__and2_1
X_9103_ clknet_leaf_43_wb_clk_i _0206_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7295_ net538 _2968_ net180 vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_9034_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[16\]
+ net209 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6246_ _1742_ _2129_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__xnor2_1
X_6177_ _1742_ _2129_ _1741_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4647__X _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5128_ net130 _1080_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4807__B _0759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5059_ _0742_ _0836_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__nand2_4
XANTENNA__4804__A1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8790__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8818_ _0421_ net192 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 _4296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8749_ _4226_ vssd1 vssd1 vccd1 vccd1 _4227_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5654__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold71 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[5\] vssd1 vssd1
+ vccd1 vccd1 net569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 team_08_WB.instance_to_wrap.allocation.game.dinoJump.button vssd1 vssd1 vccd1
+ vccd1 net558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.idle vssd1 vssd1
+ vccd1 vccd1 net580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[4\]
+ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6100_ _2024_ _2050_ _2049_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7080_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[4\]
+ _2792_ _2799_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[4\]
+ _0429_ vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8473__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4908__A _0809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6031_ _1946_ _1957_ _1983_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5039__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4793__A_N _0719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7982_ _3500_ _3502_ vssd1 vssd1 vccd1 vccd1 _3520_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_1_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6933_ _2401_ net157 _2719_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__and3b_1
X_6864_ net640 _2674_ net269 vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5458__B _1215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5815_ _1753_ _1754_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout157_A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8603_ net125 _4070_ _4074_ vssd1 vssd1 vccd1 vccd1 _4082_ sky130_fd_sc_hd__o21ai_1
X_9583_ net447 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XFILLER_0_92_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6795_ net274 _2628_ _2629_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__nor3_1
XFILLER_0_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5746_ _1697_ _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout324_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8534_ _0686_ _3683_ vssd1 vssd1 vccd1 vccd1 _4013_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5677_ _1620_ _1622_ _1624_ _1626_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_60_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8465_ _3887_ _3936_ _3944_ _3945_ _3874_ vssd1 vssd1 vccd1 vccd1 _3946_ sky130_fd_sc_hd__o2111a_1
X_4628_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[2\] vssd1
+ vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7416_ _3046_ _3060_ _3059_ vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout112_X net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8396_ _3282_ _3338_ _3355_ vssd1 vssd1 vccd1 vccd1 _3877_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_38_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4559_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[6\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__nor2_1
X_7347_ _3000_ _3008_ _3002_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7278_ _2958_ vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__inv_2
X_6229_ _2147_ _2181_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__nor2_1
X_9017_ clknet_leaf_6_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[7\]
+ net211 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_86_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4789__B1 _0634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4553__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9335__RESET_B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4961__B1 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9076__RESET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5600_ _1502_ _1552_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6580_ net621 _2486_ net263 vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5531_ _1427_ _1482_ _1481_ _1454_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4910__B _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8250_ net335 net195 vssd1 vssd1 vccd1 vccd1 _3747_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5462_ _1414_ _1413_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__and2b_1
X_7201_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[17\] _2903_ vssd1
+ vssd1 vccd1 vccd1 _2904_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8694__A1 _3305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5393_ net129 _1296_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8181_ net282 _0650_ vssd1 vssd1 vccd1 vccd1 _3699_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7132_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[11\]
+ _2850_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__nand2_1
XANTENNA__4909__Y _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7063_ team_08_WB.instance_to_wrap.allocation.game.controller.color\[10\] _2796_
+ _2809_ team_08_WB.instance_to_wrap.allocation.game.controller.color\[11\] vssd1
+ vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__a22o_1
Xfanout328 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[3\] vssd1
+ vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_2
Xfanout317 net318 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_8
XANTENNA__8892__X _4370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6014_ _1927_ _1965_ _1966_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout274_A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7965_ _3500_ _0487_ _3484_ vssd1 vssd1 vccd1 vccd1 _3504_ sky130_fd_sc_hd__mux2_1
X_7896_ net160 _3446_ net166 vssd1 vssd1 vccd1 vccd1 _3447_ sky130_fd_sc_hd__a21o_1
X_6916_ _2709_ _2710_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__nor2_1
X_9635_ net265 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6847_ _2661_ _2662_ _2663_ _2664_ vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__or4_4
XFILLER_0_43_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9566_ net434 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XFILLER_0_76_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6778_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[5\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[4\]
+ _2615_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5729_ _1679_ _1681_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5475__Y _1428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8517_ _3994_ _3996_ _3989_ vssd1 vssd1 vccd1 vccd1 _3997_ sky130_fd_sc_hd__o21ba_1
XANTENNA__4820__B _0770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9497_ net372 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__8685__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8448_ _3920_ _3928_ _3902_ vssd1 vssd1 vccd1 vccd1 _3929_ sky130_fd_sc_hd__a21oi_1
X_8379_ net174 net117 vssd1 vssd1 vccd1 vccd1 _3860_ sky130_fd_sc_hd__nand2_1
XANTENNA__7690__Y _3280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5651__B _0910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6448__A0 _2393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6999__A1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7297__C net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5098__B _1050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8373__B1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9501__376 vssd1 vssd1 vccd1 vccd1 _9501__376/HI net376 sky130_fd_sc_hd__conb_1
XFILLER_0_24_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__8676__A1 _3864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4729__Y _0684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7769__A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8061__C1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5414__A1 _0852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9257__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4962_ _0818_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7750_ net101 _3339_ _3280_ vssd1 vssd1 vccd1 vccd1 _3340_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4893_ _0821_ _0823_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__nor2_2
X_6701_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[7\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[8\]
+ _2563_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7681_ _3262_ _3270_ vssd1 vssd1 vccd1 vccd1 _3271_ sky130_fd_sc_hd__and2_2
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8903__A2 _3179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6632_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[25\] _2519_
+ _2521_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[25\]
+ sky130_fd_sc_hd__o21a_1
X_9420_ clknet_leaf_42_wb_clk_i _0365_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9351_ clknet_leaf_27_wb_clk_i _0299_ net253 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6563_ net258 _2477_ vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__nor2_2
X_5514_ _1465_ _1466_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__nand2b_1
X_8302_ net193 _3792_ _3793_ _3794_ vssd1 vssd1 vccd1 vccd1 _3795_ sky130_fd_sc_hd__a31o_1
X_9282_ clknet_leaf_5_wb_clk_i _0125_ net213 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6494_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[0\] _2429_
+ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[0\]
+ sky130_fd_sc_hd__and2b_1
X_5445_ _0769_ _0837_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__xor2_2
XANTENNA__6848__A _2665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8233_ _3733_ _3735_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8164_ net178 _3672_ vssd1 vssd1 vccd1 vccd1 _3684_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5376_ _1327_ _1328_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7115_ _2846_ _2847_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__nor2_1
Xfanout103 _3276_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_4
Xfanout147 net148 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
X_8095_ net288 _0642_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[9\]
+ vssd1 vssd1 vccd1 vccd1 _3624_ sky130_fd_sc_hd__o21a_1
Xfanout125 _3215_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_4
Xfanout114 _0236_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_4
Xfanout136 _3200_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
X_7046_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[4\]
+ _2793_ vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__or2_1
Xfanout158 _2417_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
Xfanout169 _0685_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_2
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8997_ clknet_leaf_3_wb_clk_i _0161_ net202 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_7948_ net330 _3466_ net193 vssd1 vssd1 vccd1 vccd1 _3488_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9618_ net264 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7879_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[14\]
+ _3433_ vssd1 vssd1 vccd1 vccd1 _3435_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_46_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4550__B _0422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9549_ net417 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_21_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8658__B2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold190 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8973__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8830__A1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9542__410 vssd1 vssd1 vccd1 vccd1 _9542__410/HI net410 sky130_fd_sc_hd__conb_1
XFILLER_0_95_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7528__S team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8897__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5556__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5230_ _1125_ _1127_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__xor2_2
XFILLER_0_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5161_ _1093_ _1110_ _1112_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__or3b_1
XFILLER_0_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5092_ _0821_ _0823_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6674__Y _2548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8920_ _4091_ _4092_ _4100_ vssd1 vssd1 vccd1 vccd1 _4397_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8107__B net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8851_ net330 net327 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[4\]
+ vssd1 vssd1 vccd1 vccd1 _4329_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5994_ _1942_ _1946_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7802_ net300 net298 net294 vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__mux2_1
X_8782_ _0422_ _3486_ vssd1 vssd1 vccd1 vccd1 _4260_ sky130_fd_sc_hd__and2_1
XANTENNA__9020__RESET_B net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4945_ _0841_ _0896_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7946__B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7733_ net171 _3322_ vssd1 vssd1 vccd1 vccd1 _3323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4610__A2 team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _0820_ _0827_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout237_A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8123__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7664_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[5\]
+ _3251_ _3253_ vssd1 vssd1 vccd1 vccd1 _3254_ sky130_fd_sc_hd__o21a_1
XANTENNA__8888__A1 _3888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5466__B _1417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9403_ clknet_leaf_31_wb_clk_i _0350_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6615_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[19\] _2509_
+ net255 vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7595_ _2855_ _3177_ _3184_ vssd1 vssd1 vccd1 vccd1 _3185_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_41_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9334_ clknet_leaf_53_wb_clk_i _0017_ net200 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_6546_ _2462_ _2463_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[18\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9265_ clknet_leaf_12_wb_clk_i _0087_ net226 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6477_ _0429_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[3\] _0635_
+ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5428_ _1363_ _1380_ _1361_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__a21o_1
X_9196_ clknet_leaf_16_wb_clk_i _0030_ net228 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_8216_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[10\]
+ _2989_ vssd1 vssd1 vccd1 vccd1 _3724_ sky130_fd_sc_hd__xor2_1
X_5359_ _1055_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__nor2_1
X_8147_ _0663_ net137 vssd1 vssd1 vccd1 vccd1 _3669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7076__B1 _2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8078_ _0643_ _2389_ vssd1 vssd1 vccd1 vccd1 _3608_ sky130_fd_sc_hd__and2_2
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7029_ _0435_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[2\]
+ _2777_ vssd1 vssd1 vccd1 vccd1 _2778_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4545__B net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5392__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9613__477 vssd1 vssd1 vccd1 vccd1 _9613__477/HI net477 sky130_fd_sc_hd__conb_1
XFILLER_0_40_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9466__341 vssd1 vssd1 vccd1 vccd1 _9466__341/HI net341 sky130_fd_sc_hd__conb_1
XFILLER_0_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8319__B1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4742__Y _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7790__A1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7790__B2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9507__382 vssd1 vssd1 vccd1 vccd1 _9507__382/HI net382 sky130_fd_sc_hd__conb_1
X_4730_ _0678_ _0679_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__xor2_2
XFILLER_0_71_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4661_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[2\] vssd1
+ vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7380_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\] _3028_
+ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7782__A _2368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6400_ _2335_ _2340_ _2349_ _2347_ _2346_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6331_ team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[6\] _2279_ net314
+ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4592_ net188 net185 vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6262_ _2065_ _2116_ _2115_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9050_ clknet_leaf_35_wb_clk_i _0185_ net245 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_6193_ _1348_ _2145_ _1347_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__a21o_1
X_5213_ _1110_ _1165_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8001_ _0498_ _3516_ _0483_ vssd1 vssd1 vccd1 vccd1 _3538_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_2_2__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5144_ _0820_ _0825_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9272__RESET_B net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5075_ _0979_ _0984_ _1026_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__and3_1
XANTENNA__9201__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6281__A1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8903_ _0699_ _3179_ net155 _3642_ vssd1 vssd1 vccd1 vccd1 _4380_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8022__A2 _3547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8834_ _0521_ net95 _3816_ vssd1 vssd1 vccd1 vccd1 _4312_ sky130_fd_sc_hd__and3_1
X_5977_ _1929_ _1928_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8765_ _4233_ _4242_ vssd1 vssd1 vccd1 vccd1 _4243_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_23_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4928_ _0879_ _0880_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout142_X net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8696_ net279 _2386_ vssd1 vssd1 vccd1 vccd1 _4175_ sky130_fd_sc_hd__xnor2_1
X_7716_ _3305_ vssd1 vssd1 vccd1 vccd1 _3306_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7647_ _3227_ _3236_ vssd1 vssd1 vccd1 vccd1 _3237_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _0573_ _0602_ _0781_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__nand3_4
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6336__A2 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7692__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7578_ team_08_WB.instance_to_wrap.allocation.game.game.score\[0\] _2336_ vssd1 vssd1
+ vccd1 vccd1 _3175_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_91_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9317_ clknet_leaf_3_wb_clk_i _0288_ net202 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_6529_ _2451_ _2452_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[12\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9248_ clknet_leaf_15_wb_clk_i _0099_ net218 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9179_ clknet_leaf_17_wb_clk_i _0042_ net227 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__7049__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4827__Y _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8797__B1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8028__A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8721__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5850__A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8252__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4466__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5900_ _0791_ _0921_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6880_ net635 _2684_ net269 vssd1 vssd1 vccd1 vccd1 _2686_ sky130_fd_sc_hd__o21ai_1
X_5831_ _1782_ _1783_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__and2b_1
XANTENNA__7496__B _3023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5762_ _1714_ _1713_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__nand2b_1
XANTENNA__5297__A _1048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8960__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8550_ _4005_ _4028_ vssd1 vssd1 vccd1 vccd1 _4029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_4713_ _0666_ _0667_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__or2_1
X_7501_ _3060_ _3138_ _3059_ vssd1 vssd1 vccd1 vccd1 _3139_ sky130_fd_sc_hd__o21a_1
X_5693_ _1605_ _1606_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8481_ net186 _3278_ vssd1 vssd1 vccd1 vccd1 _3961_ sky130_fd_sc_hd__nor2_1
X_4644_ _0599_ _0600_ _0574_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__a21o_4
X_7432_ _3044_ _3057_ _3074_ _3075_ vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5744__B _0905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4575_ _0483_ _0502_ _0540_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__o21ai_1
X_7363_ net233 net161 vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__nand2_2
X_6314_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[2\] _2264_ vssd1
+ vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__nand2_1
X_7294_ net180 _2967_ _2969_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout102_A _3277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9102_ clknet_leaf_43_wb_clk_i _0205_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_6245_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[18\]
+ _2196_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__and2_1
XANTENNA__5829__A1 _0919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9033_ clknet_leaf_52_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[15\]
+ net207 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6856__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6176_ _2127_ _2128_ _1787_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__a21oi_1
X_5127_ _1078_ _1079_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5058_ _0825_ _1010_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__xnor2_4
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4823__B _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8817_ net189 net331 vssd1 vssd1 vccd1 vccd1 _4295_ sky130_fd_sc_hd__and2b_1
XANTENNA__7974__X _3513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8748_ net335 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 _4226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5000__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5935__A _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8679_ _0643_ _2386_ vssd1 vssd1 vccd1 vccd1 _4158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input32_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst0.clk1
+ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8981__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1__f_wb_clk_i_X clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold72 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[18\] vssd1 vssd1
+ vccd1 vccd1 net570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.idx\[5\]
+ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[6\]
+ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_11_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6030_ _1982_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__inv_2
XANTENNA__4908__B _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7981_ net297 _3517_ _3518_ vssd1 vssd1 vccd1 vccd1 _3519_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6932_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[3\]
+ _2400_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6863_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[6\]
+ _2674_ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5814_ _0918_ _1766_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8602_ net111 _4076_ _4079_ _4080_ vssd1 vssd1 vccd1 vccd1 _4081_ sky130_fd_sc_hd__a2bb2o_1
X_9582_ net446 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XFILLER_0_88_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6794_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[10\]
+ _2625_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5745_ _1647_ _1696_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8533_ _0686_ _3683_ vssd1 vssd1 vccd1 vccd1 _4012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5676_ _1597_ _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout317_A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7673__C _3261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8464_ _3860_ _3895_ _3870_ _3345_ vssd1 vssd1 vccd1 vccd1 _3945_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_60_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4627_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[2\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[2\] vssd1
+ vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7415_ net304 net309 vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8395_ net101 _3875_ net99 vssd1 vssd1 vccd1 vccd1 _3876_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4558_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[10\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[12\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_38_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7346_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[22\]
+ _2999_ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout105_X net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5490__A _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4489_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[24\]
+ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__inv_2
X_7277_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[17\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[16\]
+ _2954_ vssd1 vssd1 vccd1 vccd1 _2958_ sky130_fd_sc_hd__and3_1
XANTENNA__8464__A2 _3895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6228_ _1247_ _1249_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__nor2_1
X_9016_ clknet_leaf_7_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[6\]
+ net211 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[6\]
+ sky130_fd_sc_hd__dfstp_4
XANTENNA__4818__B _0770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6159_ _2094_ _2111_ _2082_ vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_86_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7975__A1 _3513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7356__S _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4961__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9375__RESET_B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8976__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_75_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6662__C _2532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ _1454_ _1481_ _1482_ _1427_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_30_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5461_ _0882_ _1410_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8143__A1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7200_ net164 _2902_ _2903_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__nor3_1
XFILLER_0_42_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9045__RESET_B net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5392_ net129 _1344_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__nand2_1
X_8180_ net278 _2391_ _3697_ _3016_ vssd1 vssd1 vccd1 vccd1 _3698_ sky130_fd_sc_hd__o31a_1
XANTENNA__4704__A1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.pixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7131_ net184 _2851_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7062_ _2788_ _2795_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__nor2_1
Xfanout318 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[6\] vssd1
+ vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_4
Xfanout329 net331 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_4
Xfanout307 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
XFILLER_0_94_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6013_ _1924_ _1926_ _1925_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7964_ net193 _3501_ vssd1 vssd1 vccd1 vccd1 _3503_ sky130_fd_sc_hd__nor2_1
XANTENNA__7301__Y _2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5469__B _1421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6915_ net649 _2708_ net268 vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout267_A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7895_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[19\]
+ _3444_ vssd1 vssd1 vccd1 vccd1 _3446_ sky130_fd_sc_hd__nand2_1
XANTENNA__5266__A_N _1217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9634_ net265 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6846_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[11\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[10\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[13\]
+ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9565_ net433 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_92_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6777_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[4\]
+ _2615_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5485__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5728_ _1623_ _1680_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8516_ _3330_ _3995_ _3890_ _3274_ vssd1 vssd1 vccd1 vccd1 _3996_ sky130_fd_sc_hd__o211a_1
X_9496_ net371 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5659_ _1140_ _1600_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8447_ _3874_ _3924_ _3927_ _3922_ _3923_ vssd1 vssd1 vccd1 vccd1 _3928_ sky130_fd_sc_hd__a32o_1
X_8378_ net171 _3359_ vssd1 vssd1 vccd1 vccd1 _3859_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7329_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.remainingDelayTicks\[19\]
+ _2996_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7205__A _2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9568__496 vssd1 vssd1 vccd1 vccd1 net496 _9568__496/LO sky130_fd_sc_hd__conb_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5959__A0 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8036__A team_08_WB.instance_to_wrap.allocation.game.controller.v\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8373__A1 team_08_WB.instance_to_wrap.allocation.game.controller.v\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7884__B1 _3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4739__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7769__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8061__B1 _0654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5414__A2 _1215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4961_ net138 _0913_ _0912_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_35_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4892_ _0806_ _0843_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__xnor2_1
X_6700_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[7\]
+ _2563_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2566_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_35_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7680_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[4\]
+ _3260_ vssd1 vssd1 vccd1 vccd1 _3270_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6631_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[25\] _2519_
+ net255 vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5717__A3 _0930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9350_ clknet_leaf_31_wb_clk_i _0298_ net244 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.block_done
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8301_ net196 _3526_ net170 vssd1 vssd1 vccd1 vccd1 _3794_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6562_ _2471_ _2474_ _2475_ _2476_ vssd1 vssd1 vccd1 vccd1 _2477_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_15_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5513_ _0856_ _1459_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__xnor2_1
X_9281_ clknet_leaf_5_wb_clk_i _0124_ net203 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6493_ _0513_ net156 vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__and2b_2
XFILLER_0_15_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5444_ _0884_ _1396_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_30_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8232_ _2993_ _3734_ net122 vssd1 vssd1 vccd1 vccd1 _3735_ sky130_fd_sc_hd__a21o_1
X_8163_ net178 _3672_ vssd1 vssd1 vccd1 vccd1 _3683_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5375_ _1309_ _1326_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7114_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[7\]
+ _2844_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__a21oi_1
Xfanout104 _3272_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8094_ net288 _0642_ vssd1 vssd1 vccd1 vccd1 _3623_ sky130_fd_sc_hd__nand2_1
Xfanout137 _2418_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_4
Xfanout115 _0236_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_2
Xfanout126 net127 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_4
Xfanout148 _0777_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
Xfanout159 net160 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_7045_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[0\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.idx\[1\] vssd1
+ vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8996_ clknet_leaf_3_wb_clk_i _0160_ net204 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9483__358 vssd1 vssd1 vccd1 vccd1 _9483__358/HI net358 sky130_fd_sc_hd__conb_1
XFILLER_0_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7947_ net330 _3466_ vssd1 vssd1 vccd1 vccd1 _3487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7878_ _3433_ _3434_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[13\]
+ net166 vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8355__A1 _2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9617_ net264 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5486__Y _1439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6829_ net275 _2651_ _2652_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_46_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6366__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4831__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9524__399 vssd1 vssd1 vccd1 vccd1 _9524__399/HI net399 sky130_fd_sc_hd__conb_1
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9548_ net416 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_45_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6118__B1 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9479_ net354 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XANTENNA__5943__A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7866__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold180 team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[4\] vssd1 vssd1
+ vccd1 vccd1 net689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9067__SET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8830__A2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8594__A1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8346__A1 _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5160_ _1093_ _1110_ _1112_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_20_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5091_ _0757_ _0785_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_3_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4916__B _0861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8850_ _3871_ _3888_ _3895_ _4309_ vssd1 vssd1 vccd1 vccd1 _4328_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5993_ _1942_ _1944_ _1945_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__nand3_1
X_7801_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[5\] team_08_WB.instance_to_wrap.allocation.game.controller.state\[0\]
+ net294 vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__mux2_1
X_8781_ _3871_ _4258_ _4256_ _3933_ vssd1 vssd1 vccd1 vccd1 _4259_ sky130_fd_sc_hd__o211a_1
XANTENNA__6596__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4944_ _0841_ _0894_ _0895_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7732_ net151 _3321_ vssd1 vssd1 vccd1 vccd1 _3322_ sky130_fd_sc_hd__nand2_1
XANTENNA__8404__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8337__A1 _0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4875_ _0820_ _0827_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9402_ clknet_leaf_30_wb_clk_i _0349_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7663_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[5\]
+ net106 vssd1 vssd1 vccd1 vccd1 _3253_ sky130_fd_sc_hd__nand2_1
XANTENNA__8888__A2 _3895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6614_ _2509_ _2510_ vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[18\]
+ sky130_fd_sc_hd__nor2_1
X_7594_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[14\]
+ net184 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[13\]
+ net176 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[15\]
+ vssd1 vssd1 vccd1 vccd1 _3184_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_41_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6545_ net671 _2461_ _2429_ vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__o21ai_1
X_9333_ clknet_leaf_53_wb_clk_i _0016_ net201 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9264_ clknet_leaf_10_wb_clk_i _0086_ net226 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst0.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6476_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.state\[2\]
+ _0635_ _2261_ net574 _0429_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__a32o_1
XANTENNA__7312__A2 _2974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8215_ _3021_ _3031_ _3723_ _3002_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__a22o_1
X_5427_ _1378_ _1379_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__nor2_2
X_9195_ clknet_leaf_11_wb_clk_i _0029_ net228 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst0.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5358_ _1309_ _1310_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__nand2_1
X_8146_ net666 net243 _3668_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__o21a_1
XANTENNA__8273__B1 _3511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8077_ _3606_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\] vssd1
+ vssd1 vccd1 vccd1 _3607_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5289_ _1179_ _1181_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__xor2_1
X_7028_ net3 _2776_ vssd1 vssd1 vccd1 vccd1 _2777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold177_A team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9565__433 vssd1 vssd1 vccd1 vccd1 _9565__433/HI net433 sky130_fd_sc_hd__conb_1
XANTENNA__5003__A _0943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8979_ net311 vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9572__437 vssd1 vssd1 vccd1 vccd1 _9572__437/HI net437 sky130_fd_sc_hd__conb_1
XFILLER_0_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8984__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7067__A1 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8803__A2 _3888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6009__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8567__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8567__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5848__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_85_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8319__B2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7790__A2 _2325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4660_ _0616_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_44_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6330_ net325 _2275_ _2281_ net322 _2277_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_12_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4591_ _0554_ _0555_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6261_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[9\]
+ _2213_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6192_ _2140_ _2142_ _1394_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__a21o_1
X_5212_ _1095_ _1109_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__nor2_1
X_8000_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[4\]
+ net239 _3514_ _3537_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5143_ _0820_ _0826_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__and2_1
XANTENNA__7058__B2 _2805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4927__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _0979_ _0984_ _1026_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__a21oi_1
X_9549__417 vssd1 vssd1 vccd1 vccd1 _9549__417/HI net417 sky130_fd_sc_hd__conb_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6281__A2 _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8902_ _2285_ net125 _3627_ net134 vssd1 vssd1 vccd1 vccd1 _4379_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8833_ _4278_ _4307_ _4310_ _4284_ vssd1 vssd1 vccd1 vccd1 _4311_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9241__RESET_B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5976_ _1890_ _1892_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8134__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8764_ net319 _4232_ vssd1 vssd1 vccd1 vccd1 _4242_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4927_ _0818_ _0878_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7715_ _3261_ net107 vssd1 vssd1 vccd1 vccd1 _3305_ sky130_fd_sc_hd__and2b_2
X_8695_ _4001_ _4155_ _4173_ _4036_ vssd1 vssd1 vccd1 vccd1 _4174_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4595__A2 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4858_ _0573_ _0602_ _0781_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__and3_2
XFILLER_0_35_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7646_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[7\]
+ net110 vssd1 vssd1 vccd1 vccd1 _3236_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9595__459 vssd1 vssd1 vccd1 vccd1 _9595__459/HI net459 sky130_fd_sc_hd__conb_1
XFILLER_0_63_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7692__B net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6741__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4789_ _0736_ _0737_ _0634_ net182 vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__a211oi_4
X_7577_ net694 _2610_ _3015_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__mux2_1
X_9316_ clknet_leaf_3_wb_clk_i _0287_ net202 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.bcd_ones\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_91_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6528_ net616 _2449_ _2429_ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__o21ai_1
X_9247_ clknet_leaf_15_wb_clk_i _0098_ net215 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_6459_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[4\]
+ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.clock_div.counter\[3\]
+ _2400_ vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9178_ clknet_leaf_10_wb_clk_i _0041_ net227 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactus1size.clock_div_inst1.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8003__A_N net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8129_ net162 _0697_ _3630_ team_08_WB.instance_to_wrap.allocation.game.controller.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 _3655_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_89_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4837__A _0602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8309__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7213__A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9489__364 vssd1 vssd1 vccd1 vccd1 _9489__364/HI net364 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_67_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5668__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8979__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8721__A1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4747__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6799__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6681__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5830_ _1778_ _1780_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5761_ _0936_ _1663_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4712_ team_08_WB.instance_to_wrap.allocation.game.cactusMove.x_dist\[2\] _0647_
+ _0664_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__a21oi_1
X_7500_ net304 net308 _3041_ _3048_ vssd1 vssd1 vccd1 vccd1 _3138_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8480_ _3302_ _3959_ _3359_ net171 vssd1 vssd1 vccd1 vccd1 _3960_ sky130_fd_sc_hd__o211a_1
X_5692_ _0746_ _0765_ _1644_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7431_ net305 _3073_ vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4643_ _0574_ _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7362_ team_08_WB.instance_to_wrap.allocation.game.cactusDist.clock_div_inst1.clk1
+ _2666_ _3015_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__mux2_1
X_4574_ team_08_WB.instance_to_wrap.allocation.game.cactus1size.state\[0\] _0538_
+ _0542_ net290 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[6\]
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_97_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7293_ _2968_ vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__inv_2
X_6313_ team_08_WB.instance_to_wrap.allocation.game.cactusHeight2\[2\] _2264_ vssd1
+ vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__or2_2
XANTENNA__7017__B team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9101_ clknet_leaf_52_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.cactusMove.n_count\[31\]
+ net207 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8476__B1 _3279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6244_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.counter\[18\]
+ _2196_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9032_ clknet_leaf_51_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoDelay\[14\]
+ net209 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoDelay\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_6175_ _1785_ _1786_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout297_A team_08_WB.instance_to_wrap.allocation.game.controller.state\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5126_ _0818_ _1071_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__xnor2_1
X_5057_ _0824_ _0835_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__xor2_4
XANTENNA__4804__A3 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout252_X net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8816_ net331 net189 vssd1 vssd1 vccd1 vccd1 _4294_ sky130_fd_sc_hd__nand2b_1
X_5959_ net168 _1911_ _0747_ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_62_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8747_ _4197_ _4198_ _4224_ vssd1 vssd1 vccd1 vccd1 _4225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5935__B _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8678_ net125 _3622_ _4156_ net133 vssd1 vssd1 vccd1 vccd1 _4157_ sky130_fd_sc_hd__a22oi_1
XANTENNA__8703__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8703__B2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5517__A1 _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6714__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7629_ team_08_WB.instance_to_wrap.allocation.game.lcdOutput.framebufferIndex\[9\]
+ _3203_ net124 _3202_ vssd1 vssd1 vccd1 vccd1 _3219_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8467__B1 _3916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4838__Y _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold40 team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[23\]
+ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4854__X _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold51 _3163_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 team_08_WB.instance_to_wrap.allocation.game.cactusMove.count\[7\] vssd1 vssd1
+ vccd1 vccd1 net571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[13\] vssd1 vssd1
+ vccd1 vccd1 net582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.spi.tft_sdi vssd1
+ vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5398__A _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_45_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__8942__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8942__B2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6006__B _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7817__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8221__B team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5861__A _0919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6484__A2 team_08_WB.instance_to_wrap.allocation.game.dinoJump.dinoMovement
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7980_ _0500_ _3516_ vssd1 vssd1 vccd1 vccd1 _3518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6931_ _2400_ net157 _2718_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6862_ net273 _2673_ _2674_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__nor3_1
XFILLER_0_53_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7300__B net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9581_ net445 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
X_5813_ _1763_ _1764_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5747__A1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8933__A1 _0405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8601_ _4002_ _4054_ vssd1 vssd1 vccd1 vccd1 _4080_ sky130_fd_sc_hd__or2_1
X_6793_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[10\]
+ _2625_ team_08_WB.instance_to_wrap.allocation.game.cactus2size.clock_div_inst1.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8532_ _4009_ _4010_ vssd1 vssd1 vccd1 vccd1 _4011_ sky130_fd_sc_hd__nor2_1
X_5744_ _0773_ _0905_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5675_ _1599_ _1627_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8463_ _3302_ _3895_ _3881_ net133 vssd1 vssd1 vccd1 vccd1 _3944_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4626_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[3\]
+ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_end\[3\] vssd1
+ vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__and2b_1
XANTENNA__7028__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout212_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7414_ net302 net301 vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__nor2_2
X_8394_ net105 _3352_ net97 vssd1 vssd1 vccd1 vccd1 _3875_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7345_ _2999_ _3007_ net122 vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9016__Q team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4557_ team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[1\] team_08_WB.instance_to_wrap.allocation.game.dinoJump.count\[0\]
+ _0525_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__nor3_1
XFILLER_0_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7276_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[16\]
+ _2954_ team_08_WB.instance_to_wrap.allocation.game.controller.init_module.delay_counter\[17\]
+ vssd1 vssd1 vccd1 vccd1 _2957_ sky130_fd_sc_hd__a21o_1
X_4488_ team_08_WB.instance_to_wrap.allocation.game.scoreCounter.bcd_tens\[0\] vssd1
+ vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6227_ _2149_ _2179_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__nor2_1
X_9015_ clknet_leaf_7_wb_clk_i team_08_WB.instance_to_wrap.allocation.game.dinoJump.next_dinoY\[5\]
+ net211 vssd1 vssd1 vccd1 vccd1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_6158_ _2102_ _2110_ _2095_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__a21o_1
X_5109_ _0861_ _1003_ _1006_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_51_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7698__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6089_ _2006_ _2008_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_51_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4961__A2 _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4849__X _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_75_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_101_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6662__D _2536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6304__X _2257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5460_ _1217_ _1412_ _1411_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _1340_ _1342_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7130_ _2853_ _2860_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__or2_1
X_7061_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.x_start\[1\]
+ _2799_ _2800_ team_08_WB.instance_to_wrap.allocation.game.controller.drawBlock.y_start\[1\]
+ _2807_ vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__a221o_1
XANTENNA__8851__B1 team_08_WB.instance_to_wrap.allocation.game.collision.dinoY\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
Xfanout308 team_08_WB.instance_to_wrap.allocation.game.lcdOutput.tft.initSeqCounter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_2
X_6012_ _1962_ _1963_ _1961_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__a21bo_1
.ends

